/***********************************





************************************/


module plic(
input [7:0]addr,
input wr_n,
input oe,
input [31:0]dat_i,
output[31:0]dat_o,
output ext_int_o
);



endmodule