// Verilog netlist created by TD v4.5.12562
// Wed Apr  8 15:22:26 2020

`timescale 1ns / 1ps
module prv464_top  // ../../RTL/CPU/prv464_top.v(15)
  (
  cacheability_block,
  clk,
  hrdata,
  hready,
  hreset_n,
  hresp,
  m_ext_int,
  m_soft_int,
  m_time_int,
  mtime,
  rst,
  s_ext_int,
  haddr,
  hburst,
  hmastlock,
  hprot,
  hsize,
  htrans,
  hwdata,
  hwrite
  );

  input [31:0] cacheability_block;  // ../../RTL/CPU/prv464_top.v(17)
  input clk;  // ../../RTL/CPU/prv464_top.v(19)
  input [63:0] hrdata;  // ../../RTL/CPU/prv464_top.v(34)
  input hready;  // ../../RTL/CPU/prv464_top.v(31)
  input hreset_n;  // ../../RTL/CPU/prv464_top.v(33)
  input hresp;  // ../../RTL/CPU/prv464_top.v(32)
  input m_ext_int;  // ../../RTL/CPU/prv464_top.v(39)
  input m_soft_int;  // ../../RTL/CPU/prv464_top.v(38)
  input m_time_int;  // ../../RTL/CPU/prv464_top.v(37)
  input [63:0] mtime;  // ../../RTL/CPU/prv464_top.v(42)
  input rst;  // ../../RTL/CPU/prv464_top.v(20)
  input s_ext_int;  // ../../RTL/CPU/prv464_top.v(40)
  output [63:0] haddr;  // ../../RTL/CPU/prv464_top.v(22)
  output [2:0] hburst;  // ../../RTL/CPU/prv464_top.v(25)
  output hmastlock;  // ../../RTL/CPU/prv464_top.v(28)
  output [3:0] hprot;  // ../../RTL/CPU/prv464_top.v(26)
  output [2:0] hsize;  // ../../RTL/CPU/prv464_top.v(24)
  output [1:0] htrans;  // ../../RTL/CPU/prv464_top.v(27)
  output [63:0] hwdata;  // ../../RTL/CPU/prv464_top.v(29)
  output hwrite;  // ../../RTL/CPU/prv464_top.v(23)

  wire [63:0] addr_ex;  // ../../RTL/CPU/prv464_top.v(74)
  wire [63:0] addr_if;  // ../../RTL/CPU/prv464_top.v(65)
  wire [63:0] as1;  // ../../RTL/CPU/prv464_top.v(155)
  wire [63:0] as2;  // ../../RTL/CPU/prv464_top.v(156)
  wire [8:0] \biu/bus_unit/addr_counter ;  // ../../RTL/CPU/BIU/bus_unit.v(117)
  wire [8:0] \biu/bus_unit/last_addr ;  // ../../RTL/CPU/BIU/bus_unit.v(118)
  wire [1:0] \biu/bus_unit/mmu/i ;  // ../../RTL/CPU/BIU/mmu.v(94)
  wire [2:0] \biu/bus_unit/mmu/n39 ;
  wire [3:0] \biu/bus_unit/mmu/n40 ;
  wire [3:0] \biu/bus_unit/mmu/statu ;  // ../../RTL/CPU/BIU/mmu.v(95)
  wire [63:0] \biu/bus_unit/mmu_hwdata ;  // ../../RTL/CPU/BIU/bus_unit.v(106)
  wire [4:0] \biu/bus_unit/n26 ;
  wire [8:0] \biu/bus_unit/n39 ;
  wire [60:0] \biu/bus_unit/n49 ;
  wire [4:0] \biu/bus_unit/statu ;  // ../../RTL/CPU/BIU/bus_unit.v(115)
  wire [7:0] \biu/cache_ctrl_logic/ex_bsel ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(167)
  wire [127:0] \biu/cache_ctrl_logic/l1d_pa ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(143)
  wire [63:0] \biu/cache_ctrl_logic/l1d_pte ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(147)
  wire [63:0] \biu/cache_ctrl_logic/l1d_va ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(142)
  wire [127:0] \biu/cache_ctrl_logic/l1i_pa ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(141)
  wire [63:0] \biu/cache_ctrl_logic/l1i_pte ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(146)
  wire [63:0] \biu/cache_ctrl_logic/l1i_va ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(140)
  wire [4:0] \biu/cache_ctrl_logic/n100 ;
  wire [4:0] \biu/cache_ctrl_logic/n128 ;
  wire [7:0] \biu/cache_ctrl_logic/n182 ;
  wire [6:0] \biu/cache_ctrl_logic/n185 ;
  wire [6:0] \biu/cache_ctrl_logic/n189 ;
  wire [63:0] \biu/cache_ctrl_logic/n207 ;
  wire [63:0] \biu/cache_ctrl_logic/n209 ;
  wire [63:0] \biu/cache_ctrl_logic/n212 ;
  wire [4:0] \biu/cache_ctrl_logic/n83 ;
  wire [11:0] \biu/cache_ctrl_logic/off ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(165)
  wire [127:0] \biu/cache_ctrl_logic/pa_temp ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(136)
  wire [63:0] \biu/cache_ctrl_logic/pte_temp ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(145)
  wire [4:0] \biu/cache_ctrl_logic/statu ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(133)
  wire [1:0] \biu/ex_data_sel ;  // ../../RTL/CPU/BIU/biu.v(81)
  wire [8:0] \biu/l1d_addr ;  // ../../RTL/CPU/BIU/biu.v(96)
  wire [63:0] \biu/l1d_out ;  // ../../RTL/CPU/BIU/biu.v(92)
  wire [8:0] \biu/l1i_addr ;  // ../../RTL/CPU/BIU/biu.v(95)
  wire [63:0] \biu/l1i_in ;  // ../../RTL/CPU/BIU/biu.v(91)
  wire [63:0] \biu/maddress ;  // ../../RTL/CPU/BIU/biu.v(119)
  wire [127:0] \biu/paddress ;  // ../../RTL/CPU/BIU/biu.v(120)
  wire [31:0] cacheability_block_pad;  // ../../RTL/CPU/prv464_top.v(17)
  wire [63:0] csr_data;  // ../../RTL/CPU/prv464_top.v(54)
  wire [11:0] csr_index;  // ../../RTL/CPU/prv464_top.v(180)
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c0_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c0_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c10_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c10_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c11_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c11_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c12_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c12_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c13_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c13_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c14_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c14_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c15_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c15_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c1_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c1_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c2_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c2_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c3_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c3_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c4_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c4_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c5_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c5_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c6_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c6_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c7_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c7_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c8_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c8_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c9_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r0_c9_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c0_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c0_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c10_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c10_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c11_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c11_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c12_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c12_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c13_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c13_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c14_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c14_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c15_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c15_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c1_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c1_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c2_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c2_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c3_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c3_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c4_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c4_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c5_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c5_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c6_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c6_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c7_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c7_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c8_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c8_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c9_di ;
  wire [3:0] \cu_ru/al_ram_gpr_al_u0_r1_c9_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c0_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c0_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c10_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c10_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c11_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c11_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c12_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c12_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c13_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c13_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c14_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c14_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c15_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c15_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c1_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c1_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c2_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c2_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c3_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c3_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c4_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c4_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c5_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c5_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c6_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c6_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c7_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c7_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c8_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c8_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c9_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r0_c9_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c0_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c0_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c10_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c10_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c11_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c11_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c12_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c12_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c13_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c13_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c14_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c14_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c15_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c15_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c1_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c1_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c2_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c2_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c3_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c3_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c4_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c4_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c5_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c5_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c6_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c6_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c7_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c7_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c8_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c8_waddr ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c9_di ;
  wire [3:0] \cu_ru/al_ram_gpr_r1_c9_waddr ;
  wire [63:0] \cu_ru/m_cycle_event/n2 ;
  wire [63:0] \cu_ru/m_cycle_event/n4 ;
  wire [61:0] \cu_ru/m_s_epc/n0 ;
  wire [63:0] \cu_ru/m_s_epc/n2 ;
  wire [1:0] \cu_ru/m_s_status/n5 ;
  wire [63:0] \cu_ru/m_s_tval/n3 ;
  wire [63:0] \cu_ru/m_sie ;  // ../../RTL/CPU/CU&RU/cu_ru.v(157)
  wire [63:0] \cu_ru/m_sip ;  // ../../RTL/CPU/CU&RU/cu_ru.v(158)
  wire [63:0] \cu_ru/mcause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(161)
  wire [63:0] \cu_ru/mcycle ;  // ../../RTL/CPU/CU&RU/cu_ru.v(170)
  wire [63:0] \cu_ru/medeleg ;  // ../../RTL/CPU/CU&RU/cu_ru.v(156)
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n98 ;
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n99 ;
  wire [63:0] \cu_ru/mepc ;  // ../../RTL/CPU/CU&RU/cu_ru.v(163)
  wire [63:0] \cu_ru/mideleg ;  // ../../RTL/CPU/CU&RU/cu_ru.v(155)
  wire [63:0] \cu_ru/minstret ;  // ../../RTL/CPU/CU&RU/cu_ru.v(171)
  wire [63:0] \cu_ru/mscratch ;  // ../../RTL/CPU/CU&RU/cu_ru.v(172)
  wire [63:0] \cu_ru/mstatus ;  // ../../RTL/CPU/CU&RU/cu_ru.v(153)
  wire [63:0] \cu_ru/mtval ;  // ../../RTL/CPU/CU&RU/cu_ru.v(165)
  wire [63:0] \cu_ru/mtvec ;  // ../../RTL/CPU/CU&RU/cu_ru.v(167)
  wire [61:0] \cu_ru/n43 ;
  wire [4:0] \cu_ru/n46 ;
  wire [4:0] \cu_ru/n49 ;
  wire [4:0] \cu_ru/n52 ;
  wire [63:0] \cu_ru/n64 ;
  wire [63:0] \cu_ru/n82 ;
  wire [63:0] \cu_ru/n84 ;
  wire [63:0] \cu_ru/n90 ;
  wire [63:0] \cu_ru/scause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(162)
  wire [63:0] \cu_ru/sepc ;  // ../../RTL/CPU/CU&RU/cu_ru.v(164)
  wire [63:0] \cu_ru/sscratch ;  // ../../RTL/CPU/CU&RU/cu_ru.v(173)
  wire [63:0] \cu_ru/stval ;  // ../../RTL/CPU/CU&RU/cu_ru.v(166)
  wire [63:0] \cu_ru/stvec ;  // ../../RTL/CPU/CU&RU/cu_ru.v(168)
  wire [63:0] \cu_ru/trap_cause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(131)
  wire [63:0] \cu_ru/tvec ;  // ../../RTL/CPU/CU&RU/cu_ru.v(133)
  wire [63:0] data_csr;  // ../../RTL/CPU/prv464_top.v(182)
  wire [63:0] data_rd;  // ../../RTL/CPU/prv464_top.v(183)
  wire [63:0] ds1;  // ../../RTL/CPU/prv464_top.v(153)
  wire [63:0] ds2;  // ../../RTL/CPU/prv464_top.v(154)
  wire [11:0] ex_csr_index;  // ../../RTL/CPU/prv464_top.v(147)
  wire [63:0] ex_exc_code;  // ../../RTL/CPU/prv464_top.v(99)
  wire [63:0] ex_ins_pc;  // ../../RTL/CPU/prv464_top.v(100)
  wire [4:0] ex_rd_index;  // ../../RTL/CPU/prv464_top.v(150)
  wire [3:0] ex_size;  // ../../RTL/CPU/prv464_top.v(133)
  wire [63:0] \exu/alu_au/add_64 ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(55)
  wire [63:0] \exu/alu_au/alu_and ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(58)
  wire [63:0] \exu/alu_au/n17 ;
  wire [63:0] \exu/alu_au/n31 ;
  wire [63:0] \exu/alu_au/n33 ;
  wire [63:0] \exu/alu_au/n35 ;
  wire [63:0] \exu/alu_au/n37 ;
  wire [63:0] \exu/alu_au/n39 ;
  wire [63:0] \exu/alu_au/n47 ;
  wire [63:0] \exu/alu_au/n53 ;
  wire [63:0] \exu/alu_au/n55 ;
  wire [63:0] \exu/alu_au/sub_64 ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(56)
  wire [63:0] \exu/alu_data_mem_csr ;  // ../../RTL/CPU/EX/exu.v(193)
  wire [63:0] \exu/lsu/n1 ;
  wire [63:0] \exu/lsu/n22 ;
  wire [47:0] \exu/lsu/n25 ;
  wire [63:0] \exu/lsu/n4 ;
  wire [63:0] \exu/lsu/n52 ;
  wire [63:0] \exu/lsu/n59 ;
  wire [3:0] \exu/main_state ;  // ../../RTL/CPU/EX/exu.v(184)
  wire [7:0] \exu/n50 ;
  wire [31:0] \exu/n54 ;
  wire [63:0] \exu/n57 ;
  wire [7:0] \exu/shift_count ;  // ../../RTL/CPU/EX/exu.v(185)
  wire [63:0] haddr_pad;  // ../../RTL/CPU/prv464_top.v(22)
  wire [2:0] hburst_pad;  // ../../RTL/CPU/prv464_top.v(25)
  wire [3:0] hprot_pad;  // ../../RTL/CPU/prv464_top.v(26)
  wire [63:0] hrdata_pad;  // ../../RTL/CPU/prv464_top.v(34)
  wire [2:0] hsize_pad;  // ../../RTL/CPU/prv464_top.v(24)
  wire [1:0] htrans_pad;  // ../../RTL/CPU/prv464_top.v(27)
  wire [63:0] hwdata_pad;  // ../../RTL/CPU/prv464_top.v(29)
  wire [31:0] id_ins;  // ../../RTL/CPU/prv464_top.v(90)
  wire [63:0] id_ins_pc;  // ../../RTL/CPU/prv464_top.v(91)
  wire [4:0] id_rs1_index;  // ../../RTL/CPU/prv464_top.v(57)
  wire [4:0] id_rs2_index;  // ../../RTL/CPU/prv464_top.v(59)
  wire [7:0] \ins_dec/op_count_decode ;  // ../../RTL/CPU/ID/ins_dec.v(239)
  wire [31:0] \ins_fetch/ins_hold ;  // ../../RTL/CPU/IF/ins_fetch.v(55)
  wire [31:0] \ins_fetch/ins_shift ;  // ../../RTL/CPU/IF/ins_fetch.v(59)
  wire [61:0] \ins_fetch/n1 ;
  wire [63:0] ins_read;  // ../../RTL/CPU/prv464_top.v(67)
  wire [63:0] mtime_pad;  // ../../RTL/CPU/prv464_top.v(42)
  wire [63:0] new_pc;  // ../../RTL/CPU/prv464_top.v(184)
  wire [7:0] op_count;  // ../../RTL/CPU/prv464_top.v(157)
  wire [3:0] priv;  // ../../RTL/CPU/prv464_top.v(47)
  wire [63:0] rs1_data;  // ../../RTL/CPU/prv464_top.v(56)
  wire [63:0] satp;  // ../../RTL/CPU/prv464_top.v(46)
  wire [63:0] uncache_data;  // ../../RTL/CPU/prv464_top.v(77)
  wire [63:0] wb_exc_code;  // ../../RTL/CPU/prv464_top.v(185)
  wire [63:0] wb_ins_pc;  // ../../RTL/CPU/prv464_top.v(186)
  wire [4:0] wb_rd_index;  // ../../RTL/CPU/prv464_top.v(181)
  wire _al_n0_en;
  wire _al_u2659_o;
  wire _al_u2660_o;
  wire _al_u2662_o;
  wire _al_u2663_o;
  wire _al_u2667_o;
  wire _al_u2668_o;
  wire _al_u2670_o;
  wire _al_u2671_o;
  wire _al_u2674_o;
  wire _al_u2675_o;
  wire _al_u2677_o;
  wire _al_u2678_o;
  wire _al_u2680_o;
  wire _al_u2681_o;
  wire _al_u2683_o;
  wire _al_u2684_o;
  wire _al_u2691_o;
  wire _al_u2695_o;
  wire _al_u2697_o;
  wire _al_u2698_o;
  wire _al_u2703_o;
  wire _al_u2704_o;
  wire _al_u2705_o;
  wire _al_u2706_o;
  wire _al_u2707_o;
  wire _al_u2833_o;
  wire _al_u2835_o;
  wire _al_u2837_o;
  wire _al_u2838_o;
  wire _al_u2841_o;
  wire _al_u2842_o;
  wire _al_u2844_o;
  wire _al_u2845_o;
  wire _al_u2847_o;
  wire _al_u2848_o;
  wire _al_u2850_o;
  wire _al_u2852_o;
  wire _al_u2855_o;
  wire _al_u2856_o;
  wire _al_u2858_o;
  wire _al_u2860_o;
  wire _al_u2862_o;
  wire _al_u2864_o;
  wire _al_u2866_o;
  wire _al_u2868_o;
  wire _al_u2870_o;
  wire _al_u2873_o;
  wire _al_u2874_o;
  wire _al_u2885_o;
  wire _al_u2886_o;
  wire _al_u2889_o;
  wire _al_u2890_o;
  wire _al_u2891_o;
  wire _al_u2893_o;
  wire _al_u2895_o;
  wire _al_u2897_o;
  wire _al_u2899_o;
  wire _al_u2901_o;
  wire _al_u2903_o;
  wire _al_u2905_o;
  wire _al_u2907_o;
  wire _al_u2909_o;
  wire _al_u2910_o;
  wire _al_u2914_o;
  wire _al_u2915_o;
  wire _al_u2929_o;
  wire _al_u2930_o;
  wire _al_u2931_o;
  wire _al_u2932_o;
  wire _al_u2933_o;
  wire _al_u2934_o;
  wire _al_u2935_o;
  wire _al_u2936_o;
  wire _al_u2937_o;
  wire _al_u2938_o;
  wire _al_u2939_o;
  wire _al_u2940_o;
  wire _al_u2941_o;
  wire _al_u2942_o;
  wire _al_u2943_o;
  wire _al_u2944_o;
  wire _al_u2946_o;
  wire _al_u2948_o;
  wire _al_u2952_o;
  wire _al_u2954_o;
  wire _al_u2955_o;
  wire _al_u2956_o;
  wire _al_u2957_o;
  wire _al_u2958_o;
  wire _al_u2963_o;
  wire _al_u2964_o;
  wire _al_u2966_o;
  wire _al_u2974_o;
  wire _al_u2975_o;
  wire _al_u3033_o;
  wire _al_u3034_o;
  wire _al_u3043_o;
  wire _al_u3044_o;
  wire _al_u3046_o;
  wire _al_u3047_o;
  wire _al_u3049_o;
  wire _al_u3050_o;
  wire _al_u3052_o;
  wire _al_u3053_o;
  wire _al_u3055_o;
  wire _al_u3056_o;
  wire _al_u3058_o;
  wire _al_u3059_o;
  wire _al_u3061_o;
  wire _al_u3062_o;
  wire _al_u3064_o;
  wire _al_u3065_o;
  wire _al_u3067_o;
  wire _al_u3068_o;
  wire _al_u3070_o;
  wire _al_u3071_o;
  wire _al_u3073_o;
  wire _al_u3074_o;
  wire _al_u3076_o;
  wire _al_u3077_o;
  wire _al_u3079_o;
  wire _al_u3080_o;
  wire _al_u3082_o;
  wire _al_u3083_o;
  wire _al_u3085_o;
  wire _al_u3086_o;
  wire _al_u3088_o;
  wire _al_u3089_o;
  wire _al_u3091_o;
  wire _al_u3092_o;
  wire _al_u3094_o;
  wire _al_u3095_o;
  wire _al_u3097_o;
  wire _al_u3098_o;
  wire _al_u3100_o;
  wire _al_u3101_o;
  wire _al_u3103_o;
  wire _al_u3104_o;
  wire _al_u3106_o;
  wire _al_u3107_o;
  wire _al_u3109_o;
  wire _al_u3110_o;
  wire _al_u3112_o;
  wire _al_u3113_o;
  wire _al_u3115_o;
  wire _al_u3116_o;
  wire _al_u3118_o;
  wire _al_u3119_o;
  wire _al_u3121_o;
  wire _al_u3122_o;
  wire _al_u3124_o;
  wire _al_u3125_o;
  wire _al_u3127_o;
  wire _al_u3128_o;
  wire _al_u3130_o;
  wire _al_u3131_o;
  wire _al_u3133_o;
  wire _al_u3134_o;
  wire _al_u3136_o;
  wire _al_u3137_o;
  wire _al_u3139_o;
  wire _al_u3140_o;
  wire _al_u3142_o;
  wire _al_u3143_o;
  wire _al_u3145_o;
  wire _al_u3146_o;
  wire _al_u3148_o;
  wire _al_u3149_o;
  wire _al_u3152_o;
  wire _al_u3153_o;
  wire _al_u3155_o;
  wire _al_u3156_o;
  wire _al_u3158_o;
  wire _al_u3159_o;
  wire _al_u3161_o;
  wire _al_u3162_o;
  wire _al_u3164_o;
  wire _al_u3165_o;
  wire _al_u3167_o;
  wire _al_u3168_o;
  wire _al_u3170_o;
  wire _al_u3171_o;
  wire _al_u3173_o;
  wire _al_u3174_o;
  wire _al_u3179_o;
  wire _al_u3181_o;
  wire _al_u3183_o;
  wire _al_u3184_o;
  wire _al_u3185_o;
  wire _al_u3186_o;
  wire _al_u3187_o;
  wire _al_u3189_o;
  wire _al_u3190_o;
  wire _al_u3191_o;
  wire _al_u3194_o;
  wire _al_u3195_o;
  wire _al_u3197_o;
  wire _al_u3198_o;
  wire _al_u3200_o;
  wire _al_u3201_o;
  wire _al_u3204_o;
  wire _al_u3206_o;
  wire _al_u3209_o;
  wire _al_u3212_o;
  wire _al_u3213_o;
  wire _al_u3214_o;
  wire _al_u3216_o;
  wire _al_u3217_o;
  wire _al_u3222_o;
  wire _al_u3224_o;
  wire _al_u3237_o;
  wire _al_u3238_o;
  wire _al_u3240_o;
  wire _al_u3242_o;
  wire _al_u3244_o;
  wire _al_u3245_o;
  wire _al_u3248_o;
  wire _al_u3250_o;
  wire _al_u3252_o;
  wire _al_u3253_o;
  wire _al_u3254_o;
  wire _al_u3256_o;
  wire _al_u3258_o;
  wire _al_u3260_o;
  wire _al_u3262_o;
  wire _al_u3264_o;
  wire _al_u3266_o;
  wire _al_u3268_o;
  wire _al_u3270_o;
  wire _al_u3272_o;
  wire _al_u3274_o;
  wire _al_u3276_o;
  wire _al_u3278_o;
  wire _al_u3280_o;
  wire _al_u3282_o;
  wire _al_u3284_o;
  wire _al_u3286_o;
  wire _al_u3288_o;
  wire _al_u3290_o;
  wire _al_u3292_o;
  wire _al_u3294_o;
  wire _al_u3296_o;
  wire _al_u3298_o;
  wire _al_u3300_o;
  wire _al_u3302_o;
  wire _al_u3304_o;
  wire _al_u3306_o;
  wire _al_u3308_o;
  wire _al_u3310_o;
  wire _al_u3312_o;
  wire _al_u3314_o;
  wire _al_u3316_o;
  wire _al_u3318_o;
  wire _al_u3320_o;
  wire _al_u3322_o;
  wire _al_u3324_o;
  wire _al_u3326_o;
  wire _al_u3328_o;
  wire _al_u3330_o;
  wire _al_u3332_o;
  wire _al_u3334_o;
  wire _al_u3336_o;
  wire _al_u3338_o;
  wire _al_u3340_o;
  wire _al_u3342_o;
  wire _al_u3344_o;
  wire _al_u3346_o;
  wire _al_u3348_o;
  wire _al_u3350_o;
  wire _al_u3352_o;
  wire _al_u3354_o;
  wire _al_u3356_o;
  wire _al_u3358_o;
  wire _al_u3360_o;
  wire _al_u3362_o;
  wire _al_u3364_o;
  wire _al_u3366_o;
  wire _al_u3368_o;
  wire _al_u3370_o;
  wire _al_u3372_o;
  wire _al_u3374_o;
  wire _al_u3376_o;
  wire _al_u3378_o;
  wire _al_u3380_o;
  wire _al_u3382_o;
  wire _al_u3384_o;
  wire _al_u3387_o;
  wire _al_u3388_o;
  wire _al_u3391_o;
  wire _al_u3392_o;
  wire _al_u3393_o;
  wire _al_u3394_o;
  wire _al_u3395_o;
  wire _al_u3397_o;
  wire _al_u3399_o;
  wire _al_u3400_o;
  wire _al_u3403_o;
  wire _al_u3404_o;
  wire _al_u3407_o;
  wire _al_u3410_o;
  wire _al_u3411_o;
  wire _al_u3415_o;
  wire _al_u3420_o;
  wire _al_u3427_o;
  wire _al_u3430_o;
  wire _al_u3432_o;
  wire _al_u3433_o;
  wire _al_u3434_o;
  wire _al_u3441_o;
  wire _al_u3442_o;
  wire _al_u3443_o;
  wire _al_u3449_o;
  wire _al_u3450_o;
  wire _al_u3451_o;
  wire _al_u3456_o;
  wire _al_u3457_o;
  wire _al_u3459_o;
  wire _al_u3460_o;
  wire _al_u3464_o;
  wire _al_u3465_o;
  wire _al_u3467_o;
  wire _al_u3468_o;
  wire _al_u3472_o;
  wire _al_u3473_o;
  wire _al_u3475_o;
  wire _al_u3476_o;
  wire _al_u3480_o;
  wire _al_u3481_o;
  wire _al_u3483_o;
  wire _al_u3484_o;
  wire _al_u3488_o;
  wire _al_u3489_o;
  wire _al_u3490_o;
  wire _al_u3495_o;
  wire _al_u3496_o;
  wire _al_u3498_o;
  wire _al_u3499_o;
  wire _al_u3503_o;
  wire _al_u3504_o;
  wire _al_u3506_o;
  wire _al_u3507_o;
  wire _al_u3511_o;
  wire _al_u3512_o;
  wire _al_u3514_o;
  wire _al_u3515_o;
  wire _al_u3519_o;
  wire _al_u3520_o;
  wire _al_u3522_o;
  wire _al_u3523_o;
  wire _al_u3527_o;
  wire _al_u3528_o;
  wire _al_u3530_o;
  wire _al_u3531_o;
  wire _al_u3535_o;
  wire _al_u3536_o;
  wire _al_u3538_o;
  wire _al_u3539_o;
  wire _al_u3543_o;
  wire _al_u3544_o;
  wire _al_u3546_o;
  wire _al_u3547_o;
  wire _al_u3551_o;
  wire _al_u3552_o;
  wire _al_u3554_o;
  wire _al_u3555_o;
  wire _al_u3559_o;
  wire _al_u3560_o;
  wire _al_u3562_o;
  wire _al_u3563_o;
  wire _al_u3567_o;
  wire _al_u3568_o;
  wire _al_u3570_o;
  wire _al_u3571_o;
  wire _al_u3575_o;
  wire _al_u3576_o;
  wire _al_u3577_o;
  wire _al_u3582_o;
  wire _al_u3583_o;
  wire _al_u3585_o;
  wire _al_u3586_o;
  wire _al_u3590_o;
  wire _al_u3591_o;
  wire _al_u3593_o;
  wire _al_u3594_o;
  wire _al_u3598_o;
  wire _al_u3599_o;
  wire _al_u3601_o;
  wire _al_u3602_o;
  wire _al_u3606_o;
  wire _al_u3607_o;
  wire _al_u3609_o;
  wire _al_u3610_o;
  wire _al_u3614_o;
  wire _al_u3615_o;
  wire _al_u3617_o;
  wire _al_u3618_o;
  wire _al_u3622_o;
  wire _al_u3623_o;
  wire _al_u3625_o;
  wire _al_u3626_o;
  wire _al_u3630_o;
  wire _al_u3631_o;
  wire _al_u3633_o;
  wire _al_u3634_o;
  wire _al_u3638_o;
  wire _al_u3639_o;
  wire _al_u3641_o;
  wire _al_u3642_o;
  wire _al_u3646_o;
  wire _al_u3647_o;
  wire _al_u3649_o;
  wire _al_u3650_o;
  wire _al_u3654_o;
  wire _al_u3655_o;
  wire _al_u3657_o;
  wire _al_u3658_o;
  wire _al_u3662_o;
  wire _al_u3663_o;
  wire _al_u3664_o;
  wire _al_u3669_o;
  wire _al_u3670_o;
  wire _al_u3672_o;
  wire _al_u3673_o;
  wire _al_u3677_o;
  wire _al_u3678_o;
  wire _al_u3680_o;
  wire _al_u3681_o;
  wire _al_u3685_o;
  wire _al_u3686_o;
  wire _al_u3688_o;
  wire _al_u3689_o;
  wire _al_u3693_o;
  wire _al_u3694_o;
  wire _al_u3696_o;
  wire _al_u3697_o;
  wire _al_u3701_o;
  wire _al_u3702_o;
  wire _al_u3704_o;
  wire _al_u3705_o;
  wire _al_u3709_o;
  wire _al_u3710_o;
  wire _al_u3712_o;
  wire _al_u3713_o;
  wire _al_u3717_o;
  wire _al_u3718_o;
  wire _al_u3720_o;
  wire _al_u3721_o;
  wire _al_u3725_o;
  wire _al_u3726_o;
  wire _al_u3728_o;
  wire _al_u3729_o;
  wire _al_u3733_o;
  wire _al_u3734_o;
  wire _al_u3735_o;
  wire _al_u3740_o;
  wire _al_u3741_o;
  wire _al_u3742_o;
  wire _al_u3747_o;
  wire _al_u3748_o;
  wire _al_u3749_o;
  wire _al_u3754_o;
  wire _al_u3755_o;
  wire _al_u3756_o;
  wire _al_u3761_o;
  wire _al_u3762_o;
  wire _al_u3763_o;
  wire _al_u3768_o;
  wire _al_u3769_o;
  wire _al_u3770_o;
  wire _al_u3775_o;
  wire _al_u3776_o;
  wire _al_u3777_o;
  wire _al_u3782_o;
  wire _al_u3783_o;
  wire _al_u3784_o;
  wire _al_u3789_o;
  wire _al_u3790_o;
  wire _al_u3791_o;
  wire _al_u3796_o;
  wire _al_u3797_o;
  wire _al_u3798_o;
  wire _al_u3803_o;
  wire _al_u3804_o;
  wire _al_u3805_o;
  wire _al_u3810_o;
  wire _al_u3811_o;
  wire _al_u3812_o;
  wire _al_u3817_o;
  wire _al_u3818_o;
  wire _al_u3819_o;
  wire _al_u3824_o;
  wire _al_u3825_o;
  wire _al_u3826_o;
  wire _al_u3831_o;
  wire _al_u3832_o;
  wire _al_u3833_o;
  wire _al_u3838_o;
  wire _al_u3839_o;
  wire _al_u3840_o;
  wire _al_u3845_o;
  wire _al_u3846_o;
  wire _al_u3847_o;
  wire _al_u3852_o;
  wire _al_u3853_o;
  wire _al_u3854_o;
  wire _al_u3859_o;
  wire _al_u3860_o;
  wire _al_u3861_o;
  wire _al_u3866_o;
  wire _al_u3867_o;
  wire _al_u3868_o;
  wire _al_u3874_o;
  wire _al_u3875_o;
  wire _al_u3876_o;
  wire _al_u3882_o;
  wire _al_u3883_o;
  wire _al_u3884_o;
  wire _al_u3890_o;
  wire _al_u3891_o;
  wire _al_u3892_o;
  wire _al_u3898_o;
  wire _al_u3899_o;
  wire _al_u3900_o;
  wire _al_u3906_o;
  wire _al_u3907_o;
  wire _al_u3908_o;
  wire _al_u3913_o;
  wire _al_u3914_o;
  wire _al_u3915_o;
  wire _al_u3919_o;
  wire _al_u3923_o;
  wire _al_u3924_o;
  wire _al_u3925_o;
  wire _al_u3926_o;
  wire _al_u3927_o;
  wire _al_u3928_o;
  wire _al_u3929_o;
  wire _al_u3932_o;
  wire _al_u3938_o;
  wire _al_u3939_o;
  wire _al_u3944_o;
  wire _al_u3945_o;
  wire _al_u3947_o;
  wire _al_u3950_o;
  wire _al_u3955_o;
  wire _al_u3956_o;
  wire _al_u3969_o;
  wire _al_u3972_o;
  wire _al_u4055_o;
  wire _al_u4064_o;
  wire _al_u4066_o;
  wire _al_u4067_o;
  wire _al_u4069_o;
  wire _al_u4071_o;
  wire _al_u4072_o;
  wire _al_u4073_o;
  wire _al_u4075_o;
  wire _al_u4076_o;
  wire _al_u4077_o;
  wire _al_u4079_o;
  wire _al_u4080_o;
  wire _al_u4081_o;
  wire _al_u4083_o;
  wire _al_u4084_o;
  wire _al_u4086_o;
  wire _al_u4092_o;
  wire _al_u4094_o;
  wire _al_u4099_o;
  wire _al_u4100_o;
  wire _al_u4101_o;
  wire _al_u4106_o;
  wire _al_u4107_o;
  wire _al_u4108_o;
  wire _al_u4113_o;
  wire _al_u4117_o;
  wire _al_u4119_o;
  wire _al_u4121_o;
  wire _al_u4122_o;
  wire _al_u4123_o;
  wire _al_u4126_o;
  wire _al_u4127_o;
  wire _al_u4128_o;
  wire _al_u4131_o;
  wire _al_u4132_o;
  wire _al_u4133_o;
  wire _al_u4134_o;
  wire _al_u4135_o;
  wire _al_u4136_o;
  wire _al_u4137_o;
  wire _al_u4138_o;
  wire _al_u4139_o;
  wire _al_u4140_o;
  wire _al_u4141_o;
  wire _al_u4142_o;
  wire _al_u4143_o;
  wire _al_u4161_o;
  wire _al_u4162_o;
  wire _al_u4165_o;
  wire _al_u4166_o;
  wire _al_u4167_o;
  wire _al_u4169_o;
  wire _al_u4170_o;
  wire _al_u4172_o;
  wire _al_u4173_o;
  wire _al_u4175_o;
  wire _al_u4177_o;
  wire _al_u4178_o;
  wire _al_u4180_o;
  wire _al_u4182_o;
  wire _al_u4183_o;
  wire _al_u4185_o;
  wire _al_u4191_o;
  wire _al_u4192_o;
  wire _al_u4193_o;
  wire _al_u4194_o;
  wire _al_u4195_o;
  wire _al_u4197_o;
  wire _al_u4199_o;
  wire _al_u4200_o;
  wire _al_u4201_o;
  wire _al_u4203_o;
  wire _al_u4205_o;
  wire _al_u4207_o;
  wire _al_u4208_o;
  wire _al_u4210_o;
  wire _al_u4211_o;
  wire _al_u4213_o;
  wire _al_u4214_o;
  wire _al_u4216_o;
  wire _al_u4217_o;
  wire _al_u4219_o;
  wire _al_u4220_o;
  wire _al_u4222_o;
  wire _al_u4223_o;
  wire _al_u4225_o;
  wire _al_u4226_o;
  wire _al_u4229_o;
  wire _al_u4230_o;
  wire _al_u4232_o;
  wire _al_u4233_o;
  wire _al_u4234_o;
  wire _al_u4236_o;
  wire _al_u4237_o;
  wire _al_u4238_o;
  wire _al_u4240_o;
  wire _al_u4241_o;
  wire _al_u4242_o;
  wire _al_u4244_o;
  wire _al_u4245_o;
  wire _al_u4246_o;
  wire _al_u4248_o;
  wire _al_u4249_o;
  wire _al_u4250_o;
  wire _al_u4252_o;
  wire _al_u4253_o;
  wire _al_u4254_o;
  wire _al_u4256_o;
  wire _al_u4257_o;
  wire _al_u4258_o;
  wire _al_u4260_o;
  wire _al_u4261_o;
  wire _al_u4262_o;
  wire _al_u4264_o;
  wire _al_u4265_o;
  wire _al_u4266_o;
  wire _al_u4268_o;
  wire _al_u4269_o;
  wire _al_u4270_o;
  wire _al_u4272_o;
  wire _al_u4273_o;
  wire _al_u4274_o;
  wire _al_u4276_o;
  wire _al_u4277_o;
  wire _al_u4278_o;
  wire _al_u4280_o;
  wire _al_u4281_o;
  wire _al_u4282_o;
  wire _al_u4284_o;
  wire _al_u4285_o;
  wire _al_u4286_o;
  wire _al_u4288_o;
  wire _al_u4289_o;
  wire _al_u4290_o;
  wire _al_u4292_o;
  wire _al_u4293_o;
  wire _al_u4294_o;
  wire _al_u4296_o;
  wire _al_u4297_o;
  wire _al_u4298_o;
  wire _al_u4300_o;
  wire _al_u4301_o;
  wire _al_u4302_o;
  wire _al_u4304_o;
  wire _al_u4305_o;
  wire _al_u4306_o;
  wire _al_u4308_o;
  wire _al_u4309_o;
  wire _al_u4310_o;
  wire _al_u4312_o;
  wire _al_u4313_o;
  wire _al_u4314_o;
  wire _al_u4316_o;
  wire _al_u4317_o;
  wire _al_u4318_o;
  wire _al_u4320_o;
  wire _al_u4321_o;
  wire _al_u4322_o;
  wire _al_u4324_o;
  wire _al_u4325_o;
  wire _al_u4326_o;
  wire _al_u4328_o;
  wire _al_u4329_o;
  wire _al_u4330_o;
  wire _al_u4332_o;
  wire _al_u4333_o;
  wire _al_u4334_o;
  wire _al_u4336_o;
  wire _al_u4337_o;
  wire _al_u4338_o;
  wire _al_u4340_o;
  wire _al_u4341_o;
  wire _al_u4342_o;
  wire _al_u4344_o;
  wire _al_u4345_o;
  wire _al_u4346_o;
  wire _al_u4348_o;
  wire _al_u4349_o;
  wire _al_u4350_o;
  wire _al_u4352_o;
  wire _al_u4353_o;
  wire _al_u4354_o;
  wire _al_u4356_o;
  wire _al_u4357_o;
  wire _al_u4358_o;
  wire _al_u4360_o;
  wire _al_u4361_o;
  wire _al_u4362_o;
  wire _al_u4364_o;
  wire _al_u4365_o;
  wire _al_u4366_o;
  wire _al_u4368_o;
  wire _al_u4369_o;
  wire _al_u4370_o;
  wire _al_u4372_o;
  wire _al_u4373_o;
  wire _al_u4374_o;
  wire _al_u4376_o;
  wire _al_u4377_o;
  wire _al_u4378_o;
  wire _al_u4380_o;
  wire _al_u4381_o;
  wire _al_u4382_o;
  wire _al_u4384_o;
  wire _al_u4385_o;
  wire _al_u4386_o;
  wire _al_u4388_o;
  wire _al_u4389_o;
  wire _al_u4390_o;
  wire _al_u4392_o;
  wire _al_u4393_o;
  wire _al_u4394_o;
  wire _al_u4397_o;
  wire _al_u4398_o;
  wire _al_u4399_o;
  wire _al_u4400_o;
  wire _al_u4401_o;
  wire _al_u4402_o;
  wire _al_u4403_o;
  wire _al_u4405_o;
  wire _al_u4406_o;
  wire _al_u4407_o;
  wire _al_u4408_o;
  wire _al_u4409_o;
  wire _al_u4411_o;
  wire _al_u4412_o;
  wire _al_u4413_o;
  wire _al_u4414_o;
  wire _al_u4415_o;
  wire _al_u4417_o;
  wire _al_u4418_o;
  wire _al_u4419_o;
  wire _al_u4420_o;
  wire _al_u4421_o;
  wire _al_u4423_o;
  wire _al_u4424_o;
  wire _al_u4425_o;
  wire _al_u4426_o;
  wire _al_u4427_o;
  wire _al_u4429_o;
  wire _al_u4430_o;
  wire _al_u4431_o;
  wire _al_u4432_o;
  wire _al_u4433_o;
  wire _al_u4435_o;
  wire _al_u4436_o;
  wire _al_u4437_o;
  wire _al_u4438_o;
  wire _al_u4439_o;
  wire _al_u4441_o;
  wire _al_u4442_o;
  wire _al_u4443_o;
  wire _al_u4444_o;
  wire _al_u4445_o;
  wire _al_u4447_o;
  wire _al_u4448_o;
  wire _al_u4449_o;
  wire _al_u4450_o;
  wire _al_u4451_o;
  wire _al_u4453_o;
  wire _al_u4454_o;
  wire _al_u4455_o;
  wire _al_u4456_o;
  wire _al_u4457_o;
  wire _al_u4459_o;
  wire _al_u4460_o;
  wire _al_u4461_o;
  wire _al_u4462_o;
  wire _al_u4463_o;
  wire _al_u4465_o;
  wire _al_u4466_o;
  wire _al_u4467_o;
  wire _al_u4468_o;
  wire _al_u4469_o;
  wire _al_u4471_o;
  wire _al_u4472_o;
  wire _al_u4473_o;
  wire _al_u4474_o;
  wire _al_u4475_o;
  wire _al_u4477_o;
  wire _al_u4478_o;
  wire _al_u4479_o;
  wire _al_u4480_o;
  wire _al_u4481_o;
  wire _al_u4483_o;
  wire _al_u4484_o;
  wire _al_u4485_o;
  wire _al_u4486_o;
  wire _al_u4487_o;
  wire _al_u4489_o;
  wire _al_u4490_o;
  wire _al_u4491_o;
  wire _al_u4492_o;
  wire _al_u4493_o;
  wire _al_u4495_o;
  wire _al_u4496_o;
  wire _al_u4497_o;
  wire _al_u4498_o;
  wire _al_u4499_o;
  wire _al_u4501_o;
  wire _al_u4502_o;
  wire _al_u4503_o;
  wire _al_u4504_o;
  wire _al_u4505_o;
  wire _al_u4507_o;
  wire _al_u4508_o;
  wire _al_u4509_o;
  wire _al_u4510_o;
  wire _al_u4511_o;
  wire _al_u4513_o;
  wire _al_u4514_o;
  wire _al_u4515_o;
  wire _al_u4516_o;
  wire _al_u4517_o;
  wire _al_u4519_o;
  wire _al_u4520_o;
  wire _al_u4521_o;
  wire _al_u4522_o;
  wire _al_u4523_o;
  wire _al_u4525_o;
  wire _al_u4526_o;
  wire _al_u4527_o;
  wire _al_u4528_o;
  wire _al_u4529_o;
  wire _al_u4531_o;
  wire _al_u4532_o;
  wire _al_u4533_o;
  wire _al_u4534_o;
  wire _al_u4535_o;
  wire _al_u4537_o;
  wire _al_u4538_o;
  wire _al_u4539_o;
  wire _al_u4540_o;
  wire _al_u4541_o;
  wire _al_u4543_o;
  wire _al_u4544_o;
  wire _al_u4545_o;
  wire _al_u4546_o;
  wire _al_u4547_o;
  wire _al_u4549_o;
  wire _al_u4550_o;
  wire _al_u4551_o;
  wire _al_u4552_o;
  wire _al_u4553_o;
  wire _al_u4555_o;
  wire _al_u4556_o;
  wire _al_u4557_o;
  wire _al_u4558_o;
  wire _al_u4559_o;
  wire _al_u4561_o;
  wire _al_u4562_o;
  wire _al_u4563_o;
  wire _al_u4564_o;
  wire _al_u4565_o;
  wire _al_u4567_o;
  wire _al_u4568_o;
  wire _al_u4569_o;
  wire _al_u4570_o;
  wire _al_u4571_o;
  wire _al_u4573_o;
  wire _al_u4574_o;
  wire _al_u4575_o;
  wire _al_u4576_o;
  wire _al_u4577_o;
  wire _al_u4579_o;
  wire _al_u4580_o;
  wire _al_u4581_o;
  wire _al_u4582_o;
  wire _al_u4583_o;
  wire _al_u4585_o;
  wire _al_u4586_o;
  wire _al_u4587_o;
  wire _al_u4588_o;
  wire _al_u4589_o;
  wire _al_u4591_o;
  wire _al_u4592_o;
  wire _al_u4593_o;
  wire _al_u4594_o;
  wire _al_u4595_o;
  wire _al_u4597_o;
  wire _al_u4598_o;
  wire _al_u4599_o;
  wire _al_u4600_o;
  wire _al_u4601_o;
  wire _al_u4603_o;
  wire _al_u4604_o;
  wire _al_u4605_o;
  wire _al_u4606_o;
  wire _al_u4607_o;
  wire _al_u4609_o;
  wire _al_u4610_o;
  wire _al_u4611_o;
  wire _al_u4612_o;
  wire _al_u4613_o;
  wire _al_u4615_o;
  wire _al_u4616_o;
  wire _al_u4617_o;
  wire _al_u4618_o;
  wire _al_u4619_o;
  wire _al_u4621_o;
  wire _al_u4622_o;
  wire _al_u4623_o;
  wire _al_u4624_o;
  wire _al_u4625_o;
  wire _al_u4627_o;
  wire _al_u4628_o;
  wire _al_u4629_o;
  wire _al_u4630_o;
  wire _al_u4631_o;
  wire _al_u4633_o;
  wire _al_u4634_o;
  wire _al_u4635_o;
  wire _al_u4636_o;
  wire _al_u4637_o;
  wire _al_u4639_o;
  wire _al_u4640_o;
  wire _al_u4641_o;
  wire _al_u4642_o;
  wire _al_u4643_o;
  wire _al_u4645_o;
  wire _al_u4646_o;
  wire _al_u4647_o;
  wire _al_u4648_o;
  wire _al_u4649_o;
  wire _al_u4651_o;
  wire _al_u4652_o;
  wire _al_u4653_o;
  wire _al_u4654_o;
  wire _al_u4655_o;
  wire _al_u4657_o;
  wire _al_u4658_o;
  wire _al_u4659_o;
  wire _al_u4660_o;
  wire _al_u4661_o;
  wire _al_u4663_o;
  wire _al_u4664_o;
  wire _al_u4665_o;
  wire _al_u4666_o;
  wire _al_u4667_o;
  wire _al_u4669_o;
  wire _al_u4670_o;
  wire _al_u4671_o;
  wire _al_u4672_o;
  wire _al_u4673_o;
  wire _al_u4675_o;
  wire _al_u4676_o;
  wire _al_u4677_o;
  wire _al_u4678_o;
  wire _al_u4679_o;
  wire _al_u4681_o;
  wire _al_u4682_o;
  wire _al_u4683_o;
  wire _al_u4684_o;
  wire _al_u4685_o;
  wire _al_u4687_o;
  wire _al_u4688_o;
  wire _al_u4689_o;
  wire _al_u4690_o;
  wire _al_u4691_o;
  wire _al_u4693_o;
  wire _al_u4694_o;
  wire _al_u4695_o;
  wire _al_u4696_o;
  wire _al_u4697_o;
  wire _al_u4699_o;
  wire _al_u4700_o;
  wire _al_u4701_o;
  wire _al_u4702_o;
  wire _al_u4703_o;
  wire _al_u4705_o;
  wire _al_u4706_o;
  wire _al_u4707_o;
  wire _al_u4708_o;
  wire _al_u4709_o;
  wire _al_u4711_o;
  wire _al_u4712_o;
  wire _al_u4713_o;
  wire _al_u4714_o;
  wire _al_u4715_o;
  wire _al_u4717_o;
  wire _al_u4718_o;
  wire _al_u4719_o;
  wire _al_u4720_o;
  wire _al_u4721_o;
  wire _al_u4723_o;
  wire _al_u4724_o;
  wire _al_u4725_o;
  wire _al_u4726_o;
  wire _al_u4727_o;
  wire _al_u4729_o;
  wire _al_u4730_o;
  wire _al_u4731_o;
  wire _al_u4732_o;
  wire _al_u4733_o;
  wire _al_u4735_o;
  wire _al_u4736_o;
  wire _al_u4737_o;
  wire _al_u4738_o;
  wire _al_u4739_o;
  wire _al_u4741_o;
  wire _al_u4742_o;
  wire _al_u4743_o;
  wire _al_u4744_o;
  wire _al_u4745_o;
  wire _al_u4747_o;
  wire _al_u4748_o;
  wire _al_u4749_o;
  wire _al_u4750_o;
  wire _al_u4751_o;
  wire _al_u4753_o;
  wire _al_u4754_o;
  wire _al_u4755_o;
  wire _al_u4756_o;
  wire _al_u4757_o;
  wire _al_u4759_o;
  wire _al_u4760_o;
  wire _al_u4761_o;
  wire _al_u4762_o;
  wire _al_u4763_o;
  wire _al_u4765_o;
  wire _al_u4766_o;
  wire _al_u4768_o;
  wire _al_u4769_o;
  wire _al_u4770_o;
  wire _al_u4772_o;
  wire _al_u4773_o;
  wire _al_u4774_o;
  wire _al_u4776_o;
  wire _al_u4777_o;
  wire _al_u4778_o;
  wire _al_u4780_o;
  wire _al_u4781_o;
  wire _al_u4782_o;
  wire _al_u4784_o;
  wire _al_u4785_o;
  wire _al_u4786_o;
  wire _al_u4788_o;
  wire _al_u4789_o;
  wire _al_u4790_o;
  wire _al_u4792_o;
  wire _al_u4793_o;
  wire _al_u4794_o;
  wire _al_u4796_o;
  wire _al_u4797_o;
  wire _al_u4798_o;
  wire _al_u4801_o;
  wire _al_u4802_o;
  wire _al_u4804_o;
  wire _al_u4806_o;
  wire _al_u4808_o;
  wire _al_u4809_o;
  wire _al_u4810_o;
  wire _al_u4811_o;
  wire _al_u4812_o;
  wire _al_u4813_o;
  wire _al_u4815_o;
  wire _al_u4816_o;
  wire _al_u4817_o;
  wire _al_u4818_o;
  wire _al_u4819_o;
  wire _al_u4820_o;
  wire _al_u4822_o;
  wire _al_u4823_o;
  wire _al_u4824_o;
  wire _al_u4825_o;
  wire _al_u4826_o;
  wire _al_u4827_o;
  wire _al_u4829_o;
  wire _al_u4830_o;
  wire _al_u4831_o;
  wire _al_u4832_o;
  wire _al_u4833_o;
  wire _al_u4834_o;
  wire _al_u4835_o;
  wire _al_u4837_o;
  wire _al_u4838_o;
  wire _al_u4840_o;
  wire _al_u4841_o;
  wire _al_u4842_o;
  wire _al_u4844_o;
  wire _al_u4845_o;
  wire _al_u4846_o;
  wire _al_u4848_o;
  wire _al_u4849_o;
  wire _al_u4850_o;
  wire _al_u4852_o;
  wire _al_u4853_o;
  wire _al_u4854_o;
  wire _al_u4856_o;
  wire _al_u4857_o;
  wire _al_u4858_o;
  wire _al_u4860_o;
  wire _al_u4861_o;
  wire _al_u4862_o;
  wire _al_u4864_o;
  wire _al_u4865_o;
  wire _al_u4866_o;
  wire _al_u4868_o;
  wire _al_u4869_o;
  wire _al_u4870_o;
  wire _al_u4872_o;
  wire _al_u4875_o;
  wire _al_u5003_o;
  wire _al_u5005_o;
  wire _al_u5007_o;
  wire _al_u5009_o;
  wire _al_u5011_o;
  wire _al_u5013_o;
  wire _al_u5015_o;
  wire _al_u5017_o;
  wire _al_u5019_o;
  wire _al_u5020_o;
  wire _al_u5022_o;
  wire _al_u5023_o;
  wire _al_u5025_o;
  wire _al_u5026_o;
  wire _al_u5028_o;
  wire _al_u5029_o;
  wire _al_u5031_o;
  wire _al_u5032_o;
  wire _al_u5034_o;
  wire _al_u5035_o;
  wire _al_u5037_o;
  wire _al_u5038_o;
  wire _al_u5040_o;
  wire _al_u5041_o;
  wire _al_u5043_o;
  wire _al_u5044_o;
  wire _al_u5046_o;
  wire _al_u5047_o;
  wire _al_u5049_o;
  wire _al_u5050_o;
  wire _al_u5052_o;
  wire _al_u5053_o;
  wire _al_u5055_o;
  wire _al_u5056_o;
  wire _al_u5058_o;
  wire _al_u5059_o;
  wire _al_u5061_o;
  wire _al_u5062_o;
  wire _al_u5064_o;
  wire _al_u5065_o;
  wire _al_u5067_o;
  wire _al_u5068_o;
  wire _al_u5070_o;
  wire _al_u5071_o;
  wire _al_u5073_o;
  wire _al_u5074_o;
  wire _al_u5076_o;
  wire _al_u5077_o;
  wire _al_u5079_o;
  wire _al_u5080_o;
  wire _al_u5082_o;
  wire _al_u5083_o;
  wire _al_u5085_o;
  wire _al_u5086_o;
  wire _al_u5088_o;
  wire _al_u5089_o;
  wire _al_u5091_o;
  wire _al_u5092_o;
  wire _al_u5094_o;
  wire _al_u5095_o;
  wire _al_u5098_o;
  wire _al_u5099_o;
  wire _al_u5100_o;
  wire _al_u5101_o;
  wire _al_u5102_o;
  wire _al_u5104_o;
  wire _al_u5105_o;
  wire _al_u5106_o;
  wire _al_u5107_o;
  wire _al_u5108_o;
  wire _al_u5110_o;
  wire _al_u5111_o;
  wire _al_u5112_o;
  wire _al_u5114_o;
  wire _al_u5115_o;
  wire _al_u5116_o;
  wire _al_u5118_o;
  wire _al_u5119_o;
  wire _al_u5120_o;
  wire _al_u5122_o;
  wire _al_u5123_o;
  wire _al_u5124_o;
  wire _al_u5126_o;
  wire _al_u5127_o;
  wire _al_u5128_o;
  wire _al_u5130_o;
  wire _al_u5131_o;
  wire _al_u5132_o;
  wire _al_u5134_o;
  wire _al_u5135_o;
  wire _al_u5136_o;
  wire _al_u5138_o;
  wire _al_u5139_o;
  wire _al_u5140_o;
  wire _al_u5142_o;
  wire _al_u5143_o;
  wire _al_u5144_o;
  wire _al_u5147_o;
  wire _al_u5149_o;
  wire _al_u5151_o;
  wire _al_u5152_o;
  wire _al_u5154_o;
  wire _al_u5155_o;
  wire _al_u5156_o;
  wire _al_u5157_o;
  wire _al_u5158_o;
  wire _al_u5160_o;
  wire _al_u5161_o;
  wire _al_u5164_o;
  wire _al_u5167_o;
  wire _al_u5170_o;
  wire _al_u5173_o;
  wire _al_u5176_o;
  wire _al_u5179_o;
  wire _al_u5182_o;
  wire _al_u5185_o;
  wire _al_u5188_o;
  wire _al_u5191_o;
  wire _al_u5194_o;
  wire _al_u5197_o;
  wire _al_u5200_o;
  wire _al_u5203_o;
  wire _al_u5206_o;
  wire _al_u5209_o;
  wire _al_u5212_o;
  wire _al_u5215_o;
  wire _al_u5218_o;
  wire _al_u5221_o;
  wire _al_u5224_o;
  wire _al_u5227_o;
  wire _al_u5230_o;
  wire _al_u5233_o;
  wire _al_u5236_o;
  wire _al_u5239_o;
  wire _al_u5242_o;
  wire _al_u5245_o;
  wire _al_u5248_o;
  wire _al_u5251_o;
  wire _al_u5254_o;
  wire _al_u5257_o;
  wire _al_u5260_o;
  wire _al_u5263_o;
  wire _al_u5266_o;
  wire _al_u5269_o;
  wire _al_u5272_o;
  wire _al_u5275_o;
  wire _al_u5278_o;
  wire _al_u5281_o;
  wire _al_u5284_o;
  wire _al_u5287_o;
  wire _al_u5290_o;
  wire _al_u5293_o;
  wire _al_u5296_o;
  wire _al_u5299_o;
  wire _al_u5302_o;
  wire _al_u5305_o;
  wire _al_u5308_o;
  wire _al_u5311_o;
  wire _al_u5314_o;
  wire _al_u5317_o;
  wire _al_u5320_o;
  wire _al_u5323_o;
  wire _al_u5326_o;
  wire _al_u5329_o;
  wire _al_u5332_o;
  wire _al_u5335_o;
  wire _al_u5338_o;
  wire _al_u5341_o;
  wire _al_u5344_o;
  wire _al_u5347_o;
  wire _al_u5350_o;
  wire _al_u5353_o;
  wire _al_u5354_o;
  wire _al_u5357_o;
  wire _al_u5359_o;
  wire _al_u5361_o;
  wire _al_u5363_o;
  wire _al_u5365_o;
  wire _al_u5367_o;
  wire _al_u5369_o;
  wire _al_u5371_o;
  wire _al_u5373_o;
  wire _al_u5375_o;
  wire _al_u5377_o;
  wire _al_u5379_o;
  wire _al_u5381_o;
  wire _al_u5383_o;
  wire _al_u5385_o;
  wire _al_u5387_o;
  wire _al_u5389_o;
  wire _al_u5391_o;
  wire _al_u5393_o;
  wire _al_u5395_o;
  wire _al_u5397_o;
  wire _al_u5399_o;
  wire _al_u5401_o;
  wire _al_u5403_o;
  wire _al_u5405_o;
  wire _al_u5407_o;
  wire _al_u5409_o;
  wire _al_u5411_o;
  wire _al_u5413_o;
  wire _al_u5415_o;
  wire _al_u5417_o;
  wire _al_u5419_o;
  wire _al_u5421_o;
  wire _al_u5423_o;
  wire _al_u5425_o;
  wire _al_u5427_o;
  wire _al_u5429_o;
  wire _al_u5431_o;
  wire _al_u5433_o;
  wire _al_u5435_o;
  wire _al_u5437_o;
  wire _al_u5439_o;
  wire _al_u5441_o;
  wire _al_u5443_o;
  wire _al_u5445_o;
  wire _al_u5447_o;
  wire _al_u5449_o;
  wire _al_u5451_o;
  wire _al_u5453_o;
  wire _al_u5455_o;
  wire _al_u5457_o;
  wire _al_u5459_o;
  wire _al_u5461_o;
  wire _al_u5463_o;
  wire _al_u5465_o;
  wire _al_u5467_o;
  wire _al_u5469_o;
  wire _al_u5471_o;
  wire _al_u5473_o;
  wire _al_u5475_o;
  wire _al_u5477_o;
  wire _al_u5479_o;
  wire _al_u5481_o;
  wire _al_u5483_o;
  wire _al_u5485_o;
  wire _al_u5487_o;
  wire _al_u5489_o;
  wire _al_u5491_o;
  wire _al_u5493_o;
  wire _al_u5495_o;
  wire _al_u5497_o;
  wire _al_u5499_o;
  wire _al_u5501_o;
  wire _al_u5503_o;
  wire _al_u5505_o;
  wire _al_u5507_o;
  wire _al_u5509_o;
  wire _al_u5511_o;
  wire _al_u5513_o;
  wire _al_u5515_o;
  wire _al_u5517_o;
  wire _al_u5519_o;
  wire _al_u5521_o;
  wire _al_u5523_o;
  wire _al_u5525_o;
  wire _al_u5527_o;
  wire _al_u5529_o;
  wire _al_u5531_o;
  wire _al_u5533_o;
  wire _al_u5535_o;
  wire _al_u5537_o;
  wire _al_u5539_o;
  wire _al_u5541_o;
  wire _al_u5543_o;
  wire _al_u5545_o;
  wire _al_u5547_o;
  wire _al_u5549_o;
  wire _al_u5551_o;
  wire _al_u5553_o;
  wire _al_u5555_o;
  wire _al_u5557_o;
  wire _al_u5559_o;
  wire _al_u5561_o;
  wire _al_u5563_o;
  wire _al_u5565_o;
  wire _al_u5567_o;
  wire _al_u5569_o;
  wire _al_u5571_o;
  wire _al_u5573_o;
  wire _al_u5575_o;
  wire _al_u5577_o;
  wire _al_u5579_o;
  wire _al_u5581_o;
  wire _al_u5583_o;
  wire _al_u5585_o;
  wire _al_u5587_o;
  wire _al_u5589_o;
  wire _al_u5591_o;
  wire _al_u5593_o;
  wire _al_u5595_o;
  wire _al_u5597_o;
  wire _al_u5599_o;
  wire _al_u5601_o;
  wire _al_u5604_o;
  wire _al_u5607_o;
  wire _al_u5614_o;
  wire _al_u5662_o;
  wire _al_u5674_o;
  wire _al_u5676_o;
  wire _al_u5677_o;
  wire _al_u5678_o;
  wire _al_u5680_o;
  wire _al_u5681_o;
  wire _al_u5682_o;
  wire _al_u5684_o;
  wire _al_u5685_o;
  wire _al_u5686_o;
  wire _al_u5688_o;
  wire _al_u5689_o;
  wire _al_u5690_o;
  wire _al_u5692_o;
  wire _al_u5693_o;
  wire _al_u5694_o;
  wire _al_u5696_o;
  wire _al_u5697_o;
  wire _al_u5698_o;
  wire _al_u5700_o;
  wire _al_u5701_o;
  wire _al_u5702_o;
  wire _al_u5704_o;
  wire _al_u5705_o;
  wire _al_u5706_o;
  wire _al_u5708_o;
  wire _al_u5709_o;
  wire _al_u5710_o;
  wire _al_u5712_o;
  wire _al_u5713_o;
  wire _al_u5714_o;
  wire _al_u5716_o;
  wire _al_u5717_o;
  wire _al_u5718_o;
  wire _al_u5720_o;
  wire _al_u5721_o;
  wire _al_u5722_o;
  wire _al_u5724_o;
  wire _al_u5725_o;
  wire _al_u5726_o;
  wire _al_u5728_o;
  wire _al_u5729_o;
  wire _al_u5730_o;
  wire _al_u5732_o;
  wire _al_u5733_o;
  wire _al_u5734_o;
  wire _al_u5736_o;
  wire _al_u5737_o;
  wire _al_u5738_o;
  wire _al_u5740_o;
  wire _al_u5741_o;
  wire _al_u5742_o;
  wire _al_u5744_o;
  wire _al_u5745_o;
  wire _al_u5746_o;
  wire _al_u5748_o;
  wire _al_u5749_o;
  wire _al_u5750_o;
  wire _al_u5752_o;
  wire _al_u5753_o;
  wire _al_u5754_o;
  wire _al_u5756_o;
  wire _al_u5757_o;
  wire _al_u5758_o;
  wire _al_u5760_o;
  wire _al_u5761_o;
  wire _al_u5762_o;
  wire _al_u5764_o;
  wire _al_u5765_o;
  wire _al_u5766_o;
  wire _al_u5768_o;
  wire _al_u5769_o;
  wire _al_u5770_o;
  wire _al_u5772_o;
  wire _al_u5773_o;
  wire _al_u5774_o;
  wire _al_u5776_o;
  wire _al_u5777_o;
  wire _al_u5778_o;
  wire _al_u5780_o;
  wire _al_u5781_o;
  wire _al_u5782_o;
  wire _al_u5784_o;
  wire _al_u5785_o;
  wire _al_u5786_o;
  wire _al_u5788_o;
  wire _al_u5789_o;
  wire _al_u5790_o;
  wire _al_u5792_o;
  wire _al_u5793_o;
  wire _al_u5794_o;
  wire _al_u5796_o;
  wire _al_u5797_o;
  wire _al_u5798_o;
  wire _al_u5800_o;
  wire _al_u5801_o;
  wire _al_u5802_o;
  wire _al_u5804_o;
  wire _al_u5805_o;
  wire _al_u5806_o;
  wire _al_u5808_o;
  wire _al_u5809_o;
  wire _al_u5810_o;
  wire _al_u5812_o;
  wire _al_u5813_o;
  wire _al_u5814_o;
  wire _al_u5816_o;
  wire _al_u5817_o;
  wire _al_u5818_o;
  wire _al_u5820_o;
  wire _al_u5821_o;
  wire _al_u5822_o;
  wire _al_u5824_o;
  wire _al_u5825_o;
  wire _al_u5826_o;
  wire _al_u5828_o;
  wire _al_u5829_o;
  wire _al_u5830_o;
  wire _al_u5832_o;
  wire _al_u5833_o;
  wire _al_u5834_o;
  wire _al_u5837_o;
  wire _al_u5839_o;
  wire _al_u5841_o;
  wire _al_u5843_o;
  wire _al_u5845_o;
  wire _al_u5847_o;
  wire _al_u5850_o;
  wire _al_u5851_o;
  wire _al_u5853_o;
  wire _al_u5854_o;
  wire _al_u5856_o;
  wire _al_u5858_o;
  wire _al_u5859_o;
  wire _al_u5860_o;
  wire _al_u5862_o;
  wire _al_u5863_o;
  wire _al_u5865_o;
  wire _al_u5866_o;
  wire _al_u5868_o;
  wire _al_u5869_o;
  wire _al_u5871_o;
  wire _al_u5873_o;
  wire _al_u5874_o;
  wire _al_u5876_o;
  wire _al_u5877_o;
  wire _al_u5879_o;
  wire _al_u5880_o;
  wire _al_u5882_o;
  wire _al_u5883_o;
  wire _al_u5885_o;
  wire _al_u5887_o;
  wire _al_u5888_o;
  wire _al_u5890_o;
  wire _al_u5891_o;
  wire _al_u5893_o;
  wire _al_u5894_o;
  wire _al_u5895_o;
  wire _al_u5896_o;
  wire _al_u5898_o;
  wire _al_u5899_o;
  wire _al_u5900_o;
  wire _al_u5901_o;
  wire _al_u5903_o;
  wire _al_u5904_o;
  wire _al_u5905_o;
  wire _al_u5906_o;
  wire _al_u5908_o;
  wire _al_u5909_o;
  wire _al_u5910_o;
  wire _al_u5911_o;
  wire _al_u5913_o;
  wire _al_u5914_o;
  wire _al_u5915_o;
  wire _al_u5916_o;
  wire _al_u5918_o;
  wire _al_u5919_o;
  wire _al_u5920_o;
  wire _al_u5921_o;
  wire _al_u5923_o;
  wire _al_u5924_o;
  wire _al_u5925_o;
  wire _al_u5926_o;
  wire _al_u5928_o;
  wire _al_u5929_o;
  wire _al_u5930_o;
  wire _al_u5931_o;
  wire _al_u5933_o;
  wire _al_u5934_o;
  wire _al_u5935_o;
  wire _al_u5936_o;
  wire _al_u5938_o;
  wire _al_u5939_o;
  wire _al_u5940_o;
  wire _al_u5941_o;
  wire _al_u5942_o;
  wire _al_u5944_o;
  wire _al_u5945_o;
  wire _al_u5946_o;
  wire _al_u5947_o;
  wire _al_u5948_o;
  wire _al_u5950_o;
  wire _al_u5951_o;
  wire _al_u5952_o;
  wire _al_u5953_o;
  wire _al_u5954_o;
  wire _al_u5956_o;
  wire _al_u5957_o;
  wire _al_u5958_o;
  wire _al_u5959_o;
  wire _al_u5960_o;
  wire _al_u5962_o;
  wire _al_u5963_o;
  wire _al_u5964_o;
  wire _al_u5965_o;
  wire _al_u5966_o;
  wire _al_u5968_o;
  wire _al_u5969_o;
  wire _al_u5970_o;
  wire _al_u5971_o;
  wire _al_u5972_o;
  wire _al_u5974_o;
  wire _al_u5975_o;
  wire _al_u5976_o;
  wire _al_u5977_o;
  wire _al_u5978_o;
  wire _al_u5980_o;
  wire _al_u5981_o;
  wire _al_u5982_o;
  wire _al_u5983_o;
  wire _al_u5984_o;
  wire _al_u5986_o;
  wire _al_u5987_o;
  wire _al_u5988_o;
  wire _al_u5989_o;
  wire _al_u5990_o;
  wire _al_u5992_o;
  wire _al_u6055_o;
  wire _al_u6058_o;
  wire _al_u6059_o;
  wire _al_u6061_o;
  wire _al_u6063_o;
  wire _al_u6064_o;
  wire _al_u6065_o;
  wire _al_u6067_o;
  wire _al_u6068_o;
  wire _al_u6070_o;
  wire _al_u6071_o;
  wire _al_u6073_o;
  wire _al_u6074_o;
  wire _al_u6076_o;
  wire _al_u6077_o;
  wire _al_u6079_o;
  wire _al_u6080_o;
  wire _al_u6082_o;
  wire _al_u6083_o;
  wire _al_u6085_o;
  wire _al_u6086_o;
  wire _al_u6088_o;
  wire _al_u6089_o;
  wire _al_u6091_o;
  wire _al_u6092_o;
  wire _al_u6094_o;
  wire _al_u6095_o;
  wire _al_u6097_o;
  wire _al_u6098_o;
  wire _al_u6100_o;
  wire _al_u6101_o;
  wire _al_u6103_o;
  wire _al_u6104_o;
  wire _al_u6106_o;
  wire _al_u6107_o;
  wire _al_u6109_o;
  wire _al_u6110_o;
  wire _al_u6112_o;
  wire _al_u6113_o;
  wire _al_u6114_o;
  wire _al_u6116_o;
  wire _al_u6117_o;
  wire _al_u6119_o;
  wire _al_u6120_o;
  wire _al_u6122_o;
  wire _al_u6123_o;
  wire _al_u6125_o;
  wire _al_u6126_o;
  wire _al_u6128_o;
  wire _al_u6129_o;
  wire _al_u6131_o;
  wire _al_u6132_o;
  wire _al_u6134_o;
  wire _al_u6135_o;
  wire _al_u6137_o;
  wire _al_u6138_o;
  wire _al_u6140_o;
  wire _al_u6141_o;
  wire _al_u6143_o;
  wire _al_u6144_o;
  wire _al_u6146_o;
  wire _al_u6147_o;
  wire _al_u6149_o;
  wire _al_u6150_o;
  wire _al_u6152_o;
  wire _al_u6153_o;
  wire _al_u6155_o;
  wire _al_u6156_o;
  wire _al_u6158_o;
  wire _al_u6159_o;
  wire _al_u6161_o;
  wire _al_u6162_o;
  wire _al_u6164_o;
  wire _al_u6165_o;
  wire _al_u6167_o;
  wire _al_u6168_o;
  wire _al_u6170_o;
  wire _al_u6171_o;
  wire _al_u6173_o;
  wire _al_u6174_o;
  wire _al_u6176_o;
  wire _al_u6177_o;
  wire _al_u6179_o;
  wire _al_u6180_o;
  wire _al_u6181_o;
  wire _al_u6183_o;
  wire _al_u6184_o;
  wire _al_u6186_o;
  wire _al_u6187_o;
  wire _al_u6189_o;
  wire _al_u6190_o;
  wire _al_u6192_o;
  wire _al_u6193_o;
  wire _al_u6195_o;
  wire _al_u6196_o;
  wire _al_u6198_o;
  wire _al_u6199_o;
  wire _al_u6201_o;
  wire _al_u6202_o;
  wire _al_u6204_o;
  wire _al_u6205_o;
  wire _al_u6207_o;
  wire _al_u6208_o;
  wire _al_u6209_o;
  wire _al_u6211_o;
  wire _al_u6212_o;
  wire _al_u6213_o;
  wire _al_u6215_o;
  wire _al_u6216_o;
  wire _al_u6218_o;
  wire _al_u6219_o;
  wire _al_u6221_o;
  wire _al_u6222_o;
  wire _al_u6224_o;
  wire _al_u6225_o;
  wire _al_u6227_o;
  wire _al_u6228_o;
  wire _al_u6230_o;
  wire _al_u6231_o;
  wire _al_u6233_o;
  wire _al_u6234_o;
  wire _al_u6236_o;
  wire _al_u6237_o;
  wire _al_u6239_o;
  wire _al_u6240_o;
  wire _al_u6243_o;
  wire _al_u6244_o;
  wire _al_u6245_o;
  wire _al_u6246_o;
  wire _al_u6247_o;
  wire _al_u6248_o;
  wire _al_u6249_o;
  wire _al_u6250_o;
  wire _al_u6251_o;
  wire _al_u6254_o;
  wire _al_u6255_o;
  wire _al_u6257_o;
  wire _al_u6258_o;
  wire _al_u6259_o;
  wire _al_u6260_o;
  wire _al_u6261_o;
  wire _al_u6262_o;
  wire _al_u6263_o;
  wire _al_u6264_o;
  wire _al_u6265_o;
  wire _al_u6267_o;
  wire _al_u6268_o;
  wire _al_u6269_o;
  wire _al_u6270_o;
  wire _al_u6271_o;
  wire _al_u6272_o;
  wire _al_u6273_o;
  wire _al_u6274_o;
  wire _al_u6275_o;
  wire _al_u6276_o;
  wire _al_u6277_o;
  wire _al_u6278_o;
  wire _al_u6279_o;
  wire _al_u6280_o;
  wire _al_u6281_o;
  wire _al_u6282_o;
  wire _al_u6283_o;
  wire _al_u6284_o;
  wire _al_u6285_o;
  wire _al_u6286_o;
  wire _al_u6287_o;
  wire _al_u6288_o;
  wire _al_u6289_o;
  wire _al_u6290_o;
  wire _al_u6291_o;
  wire _al_u6292_o;
  wire _al_u6293_o;
  wire _al_u6294_o;
  wire _al_u6295_o;
  wire _al_u6296_o;
  wire _al_u6297_o;
  wire _al_u6298_o;
  wire _al_u6299_o;
  wire _al_u6300_o;
  wire _al_u6301_o;
  wire _al_u6302_o;
  wire _al_u6303_o;
  wire _al_u6304_o;
  wire _al_u6305_o;
  wire _al_u6306_o;
  wire _al_u6307_o;
  wire _al_u6308_o;
  wire _al_u6309_o;
  wire _al_u6311_o;
  wire _al_u6313_o;
  wire _al_u6319_o;
  wire _al_u6320_o;
  wire _al_u6321_o;
  wire _al_u6323_o;
  wire _al_u6326_o;
  wire _al_u6331_o;
  wire _al_u6334_o;
  wire _al_u6336_o;
  wire _al_u6339_o;
  wire _al_u6340_o;
  wire _al_u6341_o;
  wire _al_u6344_o;
  wire _al_u6346_o;
  wire _al_u6348_o;
  wire _al_u6349_o;
  wire _al_u6351_o;
  wire _al_u6352_o;
  wire _al_u6354_o;
  wire _al_u6357_o;
  wire _al_u6359_o;
  wire _al_u6360_o;
  wire _al_u6362_o;
  wire _al_u6363_o;
  wire _al_u6365_o;
  wire _al_u6366_o;
  wire _al_u6367_o;
  wire _al_u6368_o;
  wire _al_u6369_o;
  wire _al_u6370_o;
  wire _al_u6371_o;
  wire _al_u6372_o;
  wire _al_u6373_o;
  wire _al_u6374_o;
  wire _al_u6375_o;
  wire _al_u6376_o;
  wire _al_u6377_o;
  wire _al_u6378_o;
  wire _al_u6379_o;
  wire _al_u6380_o;
  wire _al_u6381_o;
  wire _al_u6382_o;
  wire _al_u6383_o;
  wire _al_u6384_o;
  wire _al_u6385_o;
  wire _al_u6386_o;
  wire _al_u6387_o;
  wire _al_u6388_o;
  wire _al_u6389_o;
  wire _al_u6390_o;
  wire _al_u6391_o;
  wire _al_u6392_o;
  wire _al_u6393_o;
  wire _al_u6394_o;
  wire _al_u6395_o;
  wire _al_u6396_o;
  wire _al_u6397_o;
  wire _al_u6398_o;
  wire _al_u6399_o;
  wire _al_u6400_o;
  wire _al_u6401_o;
  wire _al_u6402_o;
  wire _al_u6403_o;
  wire _al_u6404_o;
  wire _al_u6405_o;
  wire _al_u6406_o;
  wire _al_u6407_o;
  wire _al_u6408_o;
  wire _al_u6409_o;
  wire _al_u6410_o;
  wire _al_u6411_o;
  wire _al_u6412_o;
  wire _al_u6413_o;
  wire _al_u6414_o;
  wire _al_u6415_o;
  wire _al_u6416_o;
  wire _al_u6417_o;
  wire _al_u6418_o;
  wire _al_u6419_o;
  wire _al_u6420_o;
  wire _al_u6423_o;
  wire _al_u6425_o;
  wire _al_u6426_o;
  wire _al_u6436_o;
  wire _al_u6438_o;
  wire _al_u6441_o;
  wire _al_u6443_o;
  wire _al_u6445_o;
  wire _al_u6447_o;
  wire _al_u6449_o;
  wire _al_u6451_o;
  wire _al_u6453_o;
  wire _al_u6455_o;
  wire _al_u6457_o;
  wire _al_u6459_o;
  wire _al_u6461_o;
  wire _al_u6463_o;
  wire _al_u6465_o;
  wire _al_u6467_o;
  wire _al_u6469_o;
  wire _al_u6471_o;
  wire _al_u6473_o;
  wire _al_u6475_o;
  wire _al_u6477_o;
  wire _al_u6479_o;
  wire _al_u6481_o;
  wire _al_u6483_o;
  wire _al_u6485_o;
  wire _al_u6487_o;
  wire _al_u6489_o;
  wire _al_u6491_o;
  wire _al_u6493_o;
  wire _al_u6495_o;
  wire _al_u6497_o;
  wire _al_u6499_o;
  wire _al_u6501_o;
  wire _al_u6503_o;
  wire _al_u6505_o;
  wire _al_u6507_o;
  wire _al_u6509_o;
  wire _al_u6511_o;
  wire _al_u6513_o;
  wire _al_u6515_o;
  wire _al_u6517_o;
  wire _al_u6519_o;
  wire _al_u6521_o;
  wire _al_u6523_o;
  wire _al_u6525_o;
  wire _al_u6527_o;
  wire _al_u6529_o;
  wire _al_u6531_o;
  wire _al_u6533_o;
  wire _al_u6535_o;
  wire _al_u6537_o;
  wire _al_u6539_o;
  wire _al_u6541_o;
  wire _al_u6543_o;
  wire _al_u6545_o;
  wire _al_u6547_o;
  wire _al_u6549_o;
  wire _al_u6551_o;
  wire _al_u6553_o;
  wire _al_u6555_o;
  wire _al_u6557_o;
  wire _al_u6559_o;
  wire _al_u6561_o;
  wire _al_u6563_o;
  wire _al_u6565_o;
  wire _al_u6567_o;
  wire _al_u6570_o;
  wire _al_u6572_o;
  wire _al_u6574_o;
  wire _al_u6576_o;
  wire _al_u6578_o;
  wire _al_u6580_o;
  wire _al_u6582_o;
  wire _al_u6584_o;
  wire _al_u6586_o;
  wire _al_u6588_o;
  wire _al_u6590_o;
  wire _al_u6592_o;
  wire _al_u6594_o;
  wire _al_u6596_o;
  wire _al_u6598_o;
  wire _al_u6600_o;
  wire _al_u6602_o;
  wire _al_u6604_o;
  wire _al_u6606_o;
  wire _al_u6608_o;
  wire _al_u6610_o;
  wire _al_u6612_o;
  wire _al_u6614_o;
  wire _al_u6616_o;
  wire _al_u6618_o;
  wire _al_u6620_o;
  wire _al_u6622_o;
  wire _al_u6624_o;
  wire _al_u6626_o;
  wire _al_u6628_o;
  wire _al_u6630_o;
  wire _al_u6632_o;
  wire _al_u6634_o;
  wire _al_u6636_o;
  wire _al_u6638_o;
  wire _al_u6640_o;
  wire _al_u6642_o;
  wire _al_u6644_o;
  wire _al_u6646_o;
  wire _al_u6648_o;
  wire _al_u6650_o;
  wire _al_u6652_o;
  wire _al_u6654_o;
  wire _al_u6656_o;
  wire _al_u6658_o;
  wire _al_u6660_o;
  wire _al_u6662_o;
  wire _al_u6664_o;
  wire _al_u6666_o;
  wire _al_u6668_o;
  wire _al_u6670_o;
  wire _al_u6672_o;
  wire _al_u6674_o;
  wire _al_u6676_o;
  wire _al_u6678_o;
  wire _al_u6680_o;
  wire _al_u6682_o;
  wire _al_u6684_o;
  wire _al_u6686_o;
  wire _al_u6688_o;
  wire _al_u6690_o;
  wire _al_u6692_o;
  wire _al_u6694_o;
  wire _al_u6696_o;
  wire _al_u6698_o;
  wire _al_u6700_o;
  wire _al_u6702_o;
  wire _al_u6704_o;
  wire _al_u6706_o;
  wire _al_u6708_o;
  wire _al_u6710_o;
  wire _al_u6712_o;
  wire _al_u6714_o;
  wire _al_u6716_o;
  wire _al_u6718_o;
  wire _al_u6720_o;
  wire _al_u6722_o;
  wire _al_u6724_o;
  wire _al_u6725_o;
  wire _al_u6727_o;
  wire _al_u6729_o;
  wire _al_u6731_o;
  wire _al_u6732_o;
  wire _al_u6733_o;
  wire _al_u6734_o;
  wire _al_u6736_o;
  wire _al_u6737_o;
  wire _al_u6738_o;
  wire _al_u6739_o;
  wire _al_u6742_o;
  wire _al_u6743_o;
  wire _al_u6744_o;
  wire _al_u6746_o;
  wire _al_u6747_o;
  wire _al_u6748_o;
  wire _al_u6750_o;
  wire _al_u6751_o;
  wire _al_u6752_o;
  wire _al_u6754_o;
  wire _al_u6755_o;
  wire _al_u6757_o;
  wire _al_u6758_o;
  wire _al_u6760_o;
  wire _al_u6761_o;
  wire _al_u6763_o;
  wire _al_u6764_o;
  wire _al_u6765_o;
  wire _al_u6766_o;
  wire _al_u6768_o;
  wire _al_u6769_o;
  wire _al_u6772_o;
  wire _al_u6775_o;
  wire _al_u6777_o;
  wire _al_u6778_o;
  wire _al_u6780_o;
  wire _al_u6781_o;
  wire _al_u6784_o;
  wire _al_u6785_o;
  wire _al_u6788_o;
  wire _al_u6790_o;
  wire _al_u6791_o;
  wire _al_u6794_o;
  wire _al_u6795_o;
  wire _al_u6796_o;
  wire _al_u6797_o;
  wire _al_u6798_o;
  wire _al_u6799_o;
  wire _al_u6800_o;
  wire _al_u6801_o;
  wire _al_u6803_o;
  wire _al_u6804_o;
  wire _al_u6805_o;
  wire _al_u6806_o;
  wire _al_u6807_o;
  wire _al_u6808_o;
  wire _al_u6809_o;
  wire _al_u6810_o;
  wire _al_u6812_o;
  wire _al_u6813_o;
  wire _al_u6814_o;
  wire _al_u6815_o;
  wire _al_u6816_o;
  wire _al_u6817_o;
  wire _al_u6818_o;
  wire _al_u6819_o;
  wire _al_u6820_o;
  wire _al_u6822_o;
  wire _al_u6823_o;
  wire _al_u6824_o;
  wire _al_u6825_o;
  wire _al_u6826_o;
  wire _al_u6827_o;
  wire _al_u6828_o;
  wire _al_u6829_o;
  wire _al_u6831_o;
  wire _al_u6832_o;
  wire _al_u6833_o;
  wire _al_u6834_o;
  wire _al_u6835_o;
  wire _al_u6836_o;
  wire _al_u6837_o;
  wire _al_u6838_o;
  wire _al_u6839_o;
  wire _al_u6841_o;
  wire _al_u6842_o;
  wire _al_u6843_o;
  wire _al_u6844_o;
  wire _al_u6845_o;
  wire _al_u6846_o;
  wire _al_u6847_o;
  wire _al_u6848_o;
  wire _al_u6850_o;
  wire _al_u6851_o;
  wire _al_u6852_o;
  wire _al_u6853_o;
  wire _al_u6854_o;
  wire _al_u6855_o;
  wire _al_u6856_o;
  wire _al_u6857_o;
  wire _al_u6858_o;
  wire _al_u6860_o;
  wire _al_u6861_o;
  wire _al_u6862_o;
  wire _al_u6863_o;
  wire _al_u6864_o;
  wire _al_u6865_o;
  wire _al_u6866_o;
  wire _al_u6867_o;
  wire _al_u6868_o;
  wire _al_u6870_o;
  wire _al_u6871_o;
  wire _al_u6872_o;
  wire _al_u6873_o;
  wire _al_u6874_o;
  wire _al_u6875_o;
  wire _al_u6876_o;
  wire _al_u6877_o;
  wire _al_u6878_o;
  wire _al_u6880_o;
  wire _al_u6881_o;
  wire _al_u6882_o;
  wire _al_u6883_o;
  wire _al_u6884_o;
  wire _al_u6885_o;
  wire _al_u6886_o;
  wire _al_u6887_o;
  wire _al_u6888_o;
  wire _al_u6890_o;
  wire _al_u6891_o;
  wire _al_u6892_o;
  wire _al_u6893_o;
  wire _al_u6894_o;
  wire _al_u6895_o;
  wire _al_u6896_o;
  wire _al_u6897_o;
  wire _al_u6899_o;
  wire _al_u6900_o;
  wire _al_u6901_o;
  wire _al_u6902_o;
  wire _al_u6903_o;
  wire _al_u6904_o;
  wire _al_u6905_o;
  wire _al_u6906_o;
  wire _al_u6908_o;
  wire _al_u6909_o;
  wire _al_u6910_o;
  wire _al_u6911_o;
  wire _al_u6912_o;
  wire _al_u6913_o;
  wire _al_u6914_o;
  wire _al_u6915_o;
  wire _al_u6917_o;
  wire _al_u6918_o;
  wire _al_u6919_o;
  wire _al_u6920_o;
  wire _al_u6921_o;
  wire _al_u6922_o;
  wire _al_u6923_o;
  wire _al_u6924_o;
  wire _al_u6926_o;
  wire _al_u6927_o;
  wire _al_u6928_o;
  wire _al_u6929_o;
  wire _al_u6930_o;
  wire _al_u6931_o;
  wire _al_u6932_o;
  wire _al_u6933_o;
  wire _al_u6935_o;
  wire _al_u6936_o;
  wire _al_u6938_o;
  wire _al_u6939_o;
  wire _al_u6940_o;
  wire _al_u6942_o;
  wire _al_u6943_o;
  wire _al_u6945_o;
  wire _al_u6947_o;
  wire _al_u6948_o;
  wire _al_u6949_o;
  wire _al_u6950_o;
  wire _al_u6951_o;
  wire _al_u6952_o;
  wire _al_u6953_o;
  wire _al_u6954_o;
  wire _al_u6955_o;
  wire _al_u6957_o;
  wire _al_u6958_o;
  wire _al_u6959_o;
  wire _al_u6960_o;
  wire _al_u6961_o;
  wire _al_u6962_o;
  wire _al_u6963_o;
  wire _al_u6964_o;
  wire _al_u6965_o;
  wire _al_u6967_o;
  wire _al_u6968_o;
  wire _al_u6969_o;
  wire _al_u6970_o;
  wire _al_u6971_o;
  wire _al_u6972_o;
  wire _al_u6973_o;
  wire _al_u6974_o;
  wire _al_u6975_o;
  wire _al_u6977_o;
  wire _al_u6978_o;
  wire _al_u6979_o;
  wire _al_u6980_o;
  wire _al_u6981_o;
  wire _al_u6982_o;
  wire _al_u6983_o;
  wire _al_u6984_o;
  wire _al_u6985_o;
  wire _al_u6987_o;
  wire _al_u6988_o;
  wire _al_u6989_o;
  wire _al_u6990_o;
  wire _al_u6991_o;
  wire _al_u6992_o;
  wire _al_u6993_o;
  wire _al_u6994_o;
  wire _al_u6995_o;
  wire _al_u6997_o;
  wire _al_u6998_o;
  wire _al_u6999_o;
  wire _al_u7000_o;
  wire _al_u7001_o;
  wire _al_u7002_o;
  wire _al_u7003_o;
  wire _al_u7004_o;
  wire _al_u7005_o;
  wire _al_u7006_o;
  wire _al_u7008_o;
  wire _al_u7009_o;
  wire _al_u7010_o;
  wire _al_u7011_o;
  wire _al_u7012_o;
  wire _al_u7013_o;
  wire _al_u7014_o;
  wire _al_u7015_o;
  wire _al_u7016_o;
  wire _al_u7018_o;
  wire _al_u7019_o;
  wire _al_u7020_o;
  wire _al_u7021_o;
  wire _al_u7022_o;
  wire _al_u7023_o;
  wire _al_u7024_o;
  wire _al_u7025_o;
  wire _al_u7026_o;
  wire _al_u7028_o;
  wire _al_u7029_o;
  wire _al_u7030_o;
  wire _al_u7031_o;
  wire _al_u7032_o;
  wire _al_u7033_o;
  wire _al_u7034_o;
  wire _al_u7035_o;
  wire _al_u7036_o;
  wire _al_u7038_o;
  wire _al_u7039_o;
  wire _al_u7040_o;
  wire _al_u7041_o;
  wire _al_u7042_o;
  wire _al_u7043_o;
  wire _al_u7044_o;
  wire _al_u7045_o;
  wire _al_u7046_o;
  wire _al_u7048_o;
  wire _al_u7049_o;
  wire _al_u7050_o;
  wire _al_u7051_o;
  wire _al_u7052_o;
  wire _al_u7053_o;
  wire _al_u7054_o;
  wire _al_u7055_o;
  wire _al_u7056_o;
  wire _al_u7058_o;
  wire _al_u7059_o;
  wire _al_u7060_o;
  wire _al_u7061_o;
  wire _al_u7062_o;
  wire _al_u7063_o;
  wire _al_u7064_o;
  wire _al_u7065_o;
  wire _al_u7066_o;
  wire _al_u7068_o;
  wire _al_u7069_o;
  wire _al_u7070_o;
  wire _al_u7071_o;
  wire _al_u7072_o;
  wire _al_u7073_o;
  wire _al_u7074_o;
  wire _al_u7075_o;
  wire _al_u7076_o;
  wire _al_u7078_o;
  wire _al_u7079_o;
  wire _al_u7080_o;
  wire _al_u7081_o;
  wire _al_u7082_o;
  wire _al_u7083_o;
  wire _al_u7084_o;
  wire _al_u7085_o;
  wire _al_u7086_o;
  wire _al_u7088_o;
  wire _al_u7089_o;
  wire _al_u7090_o;
  wire _al_u7091_o;
  wire _al_u7092_o;
  wire _al_u7093_o;
  wire _al_u7094_o;
  wire _al_u7095_o;
  wire _al_u7096_o;
  wire _al_u7098_o;
  wire _al_u7099_o;
  wire _al_u7100_o;
  wire _al_u7101_o;
  wire _al_u7102_o;
  wire _al_u7103_o;
  wire _al_u7104_o;
  wire _al_u7105_o;
  wire _al_u7106_o;
  wire _al_u7107_o;
  wire _al_u7109_o;
  wire _al_u7110_o;
  wire _al_u7111_o;
  wire _al_u7112_o;
  wire _al_u7113_o;
  wire _al_u7114_o;
  wire _al_u7115_o;
  wire _al_u7116_o;
  wire _al_u7117_o;
  wire _al_u7118_o;
  wire _al_u7120_o;
  wire _al_u7121_o;
  wire _al_u7122_o;
  wire _al_u7123_o;
  wire _al_u7124_o;
  wire _al_u7125_o;
  wire _al_u7126_o;
  wire _al_u7127_o;
  wire _al_u7128_o;
  wire _al_u7129_o;
  wire _al_u7131_o;
  wire _al_u7132_o;
  wire _al_u7133_o;
  wire _al_u7134_o;
  wire _al_u7135_o;
  wire _al_u7136_o;
  wire _al_u7137_o;
  wire _al_u7138_o;
  wire _al_u7139_o;
  wire _al_u7141_o;
  wire _al_u7142_o;
  wire _al_u7145_o;
  wire _al_u7146_o;
  wire _al_u7147_o;
  wire _al_u7149_o;
  wire _al_u7150_o;
  wire _al_u7151_o;
  wire _al_u7152_o;
  wire _al_u7154_o;
  wire _al_u7155_o;
  wire _al_u7156_o;
  wire _al_u7157_o;
  wire _al_u7158_o;
  wire _al_u7159_o;
  wire _al_u7160_o;
  wire _al_u7161_o;
  wire _al_u7162_o;
  wire _al_u7163_o;
  wire _al_u7164_o;
  wire _al_u7165_o;
  wire _al_u7166_o;
  wire _al_u7167_o;
  wire _al_u7168_o;
  wire _al_u7169_o;
  wire _al_u7170_o;
  wire _al_u7171_o;
  wire _al_u7172_o;
  wire _al_u7173_o;
  wire _al_u7174_o;
  wire _al_u7175_o;
  wire _al_u7176_o;
  wire _al_u7177_o;
  wire _al_u7178_o;
  wire _al_u7179_o;
  wire _al_u7180_o;
  wire _al_u7181_o;
  wire _al_u7182_o;
  wire _al_u7183_o;
  wire _al_u7184_o;
  wire _al_u7185_o;
  wire _al_u7186_o;
  wire _al_u7187_o;
  wire _al_u7188_o;
  wire _al_u7190_o;
  wire _al_u7191_o;
  wire _al_u7192_o;
  wire _al_u7193_o;
  wire _al_u7195_o;
  wire _al_u7198_o;
  wire _al_u7199_o;
  wire _al_u7200_o;
  wire _al_u7201_o;
  wire _al_u7202_o;
  wire _al_u7203_o;
  wire _al_u7205_o;
  wire _al_u7206_o;
  wire _al_u7208_o;
  wire _al_u7210_o;
  wire _al_u7211_o;
  wire _al_u7212_o;
  wire _al_u7214_o;
  wire _al_u7215_o;
  wire _al_u7216_o;
  wire _al_u7218_o;
  wire _al_u7219_o;
  wire _al_u7220_o;
  wire _al_u7221_o;
  wire _al_u7222_o;
  wire _al_u7223_o;
  wire _al_u7224_o;
  wire _al_u7226_o;
  wire _al_u7227_o;
  wire _al_u7228_o;
  wire _al_u7229_o;
  wire _al_u7230_o;
  wire _al_u7231_o;
  wire _al_u7232_o;
  wire _al_u7233_o;
  wire _al_u7234_o;
  wire _al_u7235_o;
  wire _al_u7237_o;
  wire _al_u7238_o;
  wire _al_u7239_o;
  wire _al_u7240_o;
  wire _al_u7242_o;
  wire _al_u7243_o;
  wire _al_u7244_o;
  wire _al_u7245_o;
  wire _al_u7246_o;
  wire _al_u7247_o;
  wire _al_u7248_o;
  wire _al_u7249_o;
  wire _al_u7251_o;
  wire _al_u7252_o;
  wire _al_u7253_o;
  wire _al_u7254_o;
  wire _al_u7255_o;
  wire _al_u7256_o;
  wire _al_u7257_o;
  wire _al_u7258_o;
  wire _al_u7259_o;
  wire _al_u7260_o;
  wire _al_u7262_o;
  wire _al_u7263_o;
  wire _al_u7264_o;
  wire _al_u7266_o;
  wire _al_u7267_o;
  wire _al_u7268_o;
  wire _al_u7269_o;
  wire _al_u7270_o;
  wire _al_u7271_o;
  wire _al_u7272_o;
  wire _al_u7274_o;
  wire _al_u7275_o;
  wire _al_u7276_o;
  wire _al_u7277_o;
  wire _al_u7278_o;
  wire _al_u7279_o;
  wire _al_u7280_o;
  wire _al_u7281_o;
  wire _al_u7282_o;
  wire _al_u7283_o;
  wire _al_u7285_o;
  wire _al_u7287_o;
  wire _al_u7288_o;
  wire _al_u7289_o;
  wire _al_u7290_o;
  wire _al_u7291_o;
  wire _al_u7292_o;
  wire _al_u7293_o;
  wire _al_u7294_o;
  wire _al_u7295_o;
  wire _al_u7296_o;
  wire _al_u7330_o;
  wire _al_u7331_o;
  wire _al_u7333_o;
  wire _al_u7335_o;
  wire _al_u7337_o;
  wire _al_u7339_o;
  wire _al_u7340_o;
  wire _al_u7341_o;
  wire _al_u7342_o;
  wire _al_u7343_o;
  wire _al_u7344_o;
  wire _al_u7345_o;
  wire _al_u7346_o;
  wire _al_u7347_o;
  wire _al_u7348_o;
  wire _al_u7349_o;
  wire _al_u7351_o;
  wire _al_u7352_o;
  wire _al_u7353_o;
  wire _al_u7355_o;
  wire _al_u7356_o;
  wire _al_u7358_o;
  wire _al_u7359_o;
  wire _al_u7361_o;
  wire _al_u7362_o;
  wire _al_u7364_o;
  wire _al_u7365_o;
  wire _al_u7367_o;
  wire _al_u7368_o;
  wire _al_u7370_o;
  wire _al_u7371_o;
  wire _al_u7373_o;
  wire _al_u7374_o;
  wire _al_u7376_o;
  wire _al_u7377_o;
  wire _al_u7379_o;
  wire _al_u7380_o;
  wire _al_u7382_o;
  wire _al_u7383_o;
  wire _al_u7385_o;
  wire _al_u7386_o;
  wire _al_u7388_o;
  wire _al_u7389_o;
  wire _al_u7391_o;
  wire _al_u7392_o;
  wire _al_u7394_o;
  wire _al_u7395_o;
  wire _al_u7397_o;
  wire _al_u7398_o;
  wire _al_u7401_o;
  wire _al_u7402_o;
  wire _al_u7403_o;
  wire _al_u7404_o;
  wire _al_u7405_o;
  wire _al_u7406_o;
  wire _al_u7407_o;
  wire _al_u7408_o;
  wire _al_u7409_o;
  wire _al_u7410_o;
  wire _al_u7411_o;
  wire _al_u7413_o;
  wire _al_u7414_o;
  wire _al_u7415_o;
  wire _al_u7416_o;
  wire _al_u7417_o;
  wire _al_u7418_o;
  wire _al_u7419_o;
  wire _al_u7420_o;
  wire _al_u7421_o;
  wire _al_u7422_o;
  wire _al_u7424_o;
  wire _al_u7425_o;
  wire _al_u7426_o;
  wire _al_u7427_o;
  wire _al_u7428_o;
  wire _al_u7429_o;
  wire _al_u7430_o;
  wire _al_u7431_o;
  wire _al_u7432_o;
  wire _al_u7433_o;
  wire _al_u7434_o;
  wire _al_u7436_o;
  wire _al_u7437_o;
  wire _al_u7438_o;
  wire _al_u7439_o;
  wire _al_u7440_o;
  wire _al_u7441_o;
  wire _al_u7442_o;
  wire _al_u7443_o;
  wire _al_u7444_o;
  wire _al_u7445_o;
  wire _al_u7447_o;
  wire _al_u7448_o;
  wire _al_u7449_o;
  wire _al_u7450_o;
  wire _al_u7451_o;
  wire _al_u7452_o;
  wire _al_u7453_o;
  wire _al_u7454_o;
  wire _al_u7455_o;
  wire _al_u7456_o;
  wire _al_u7457_o;
  wire _al_u7459_o;
  wire _al_u7460_o;
  wire _al_u7461_o;
  wire _al_u7462_o;
  wire _al_u7463_o;
  wire _al_u7464_o;
  wire _al_u7465_o;
  wire _al_u7466_o;
  wire _al_u7467_o;
  wire _al_u7468_o;
  wire _al_u7470_o;
  wire _al_u7471_o;
  wire _al_u7472_o;
  wire _al_u7473_o;
  wire _al_u7474_o;
  wire _al_u7475_o;
  wire _al_u7476_o;
  wire _al_u7477_o;
  wire _al_u7478_o;
  wire _al_u7480_o;
  wire _al_u7481_o;
  wire _al_u7482_o;
  wire _al_u7483_o;
  wire _al_u7485_o;
  wire _al_u7486_o;
  wire _al_u7487_o;
  wire _al_u7488_o;
  wire _al_u7489_o;
  wire _al_u7491_o;
  wire _al_u7492_o;
  wire _al_u7493_o;
  wire _al_u7494_o;
  wire _al_u7495_o;
  wire _al_u7497_o;
  wire _al_u7498_o;
  wire _al_u7499_o;
  wire _al_u7500_o;
  wire _al_u7501_o;
  wire _al_u7502_o;
  wire _al_u7503_o;
  wire _al_u7504_o;
  wire _al_u7505_o;
  wire _al_u7506_o;
  wire _al_u7507_o;
  wire _al_u7508_o;
  wire _al_u7510_o;
  wire _al_u7511_o;
  wire _al_u7512_o;
  wire _al_u7514_o;
  wire _al_u7515_o;
  wire _al_u7516_o;
  wire _al_u7518_o;
  wire _al_u7519_o;
  wire _al_u7520_o;
  wire _al_u7522_o;
  wire _al_u7523_o;
  wire _al_u7524_o;
  wire _al_u7526_o;
  wire _al_u7527_o;
  wire _al_u7528_o;
  wire _al_u7530_o;
  wire _al_u7531_o;
  wire _al_u7533_o;
  wire _al_u7534_o;
  wire _al_u7535_o;
  wire _al_u7537_o;
  wire _al_u7538_o;
  wire _al_u7539_o;
  wire _al_u7541_o;
  wire _al_u7542_o;
  wire _al_u7543_o;
  wire _al_u7544_o;
  wire _al_u7545_o;
  wire _al_u7546_o;
  wire _al_u7547_o;
  wire _al_u7548_o;
  wire _al_u7549_o;
  wire _al_u7550_o;
  wire _al_u7551_o;
  wire _al_u7553_o;
  wire _al_u7554_o;
  wire _al_u7555_o;
  wire _al_u7557_o;
  wire _al_u7558_o;
  wire _al_u7559_o;
  wire _al_u7561_o;
  wire _al_u7562_o;
  wire _al_u7563_o;
  wire _al_u7565_o;
  wire _al_u7566_o;
  wire _al_u7567_o;
  wire _al_u7569_o;
  wire _al_u7570_o;
  wire _al_u7571_o;
  wire _al_u7573_o;
  wire _al_u7574_o;
  wire _al_u7575_o;
  wire _al_u7576_o;
  wire _al_u7577_o;
  wire _al_u7578_o;
  wire _al_u7579_o;
  wire _al_u7580_o;
  wire _al_u7581_o;
  wire _al_u7582_o;
  wire _al_u7583_o;
  wire _al_u7585_o;
  wire _al_u7586_o;
  wire _al_u7588_o;
  wire _al_u7589_o;
  wire _al_u7591_o;
  wire _al_u7592_o;
  wire _al_u7594_o;
  wire _al_u7595_o;
  wire _al_u7597_o;
  wire _al_u7598_o;
  wire _al_u7600_o;
  wire _al_u7601_o;
  wire _al_u7602_o;
  wire _al_u7603_o;
  wire _al_u7604_o;
  wire _al_u7605_o;
  wire _al_u7606_o;
  wire _al_u7607_o;
  wire _al_u7608_o;
  wire _al_u7609_o;
  wire _al_u7610_o;
  wire _al_u7612_o;
  wire _al_u7613_o;
  wire _al_u7614_o;
  wire _al_u7615_o;
  wire _al_u7616_o;
  wire _al_u7617_o;
  wire _al_u7618_o;
  wire _al_u7619_o;
  wire _al_u7620_o;
  wire _al_u7621_o;
  wire _al_u7622_o;
  wire _al_u7624_o;
  wire _al_u7625_o;
  wire _al_u7626_o;
  wire _al_u7627_o;
  wire _al_u7628_o;
  wire _al_u7629_o;
  wire _al_u7630_o;
  wire _al_u7631_o;
  wire _al_u7632_o;
  wire _al_u7633_o;
  wire _al_u7634_o;
  wire _al_u7635_o;
  wire _al_u7637_o;
  wire _al_u7638_o;
  wire _al_u7639_o;
  wire _al_u7640_o;
  wire _al_u7641_o;
  wire _al_u7642_o;
  wire _al_u7643_o;
  wire _al_u7644_o;
  wire _al_u7645_o;
  wire _al_u7646_o;
  wire _al_u7647_o;
  wire _al_u7649_o;
  wire _al_u7650_o;
  wire _al_u7652_o;
  wire _al_u7653_o;
  wire _al_u7654_o;
  wire _al_u7655_o;
  wire _al_u7656_o;
  wire _al_u7657_o;
  wire _al_u7658_o;
  wire _al_u7659_o;
  wire _al_u7660_o;
  wire _al_u7661_o;
  wire _al_u7662_o;
  wire _al_u7663_o;
  wire _al_u7665_o;
  wire _al_u7666_o;
  wire _al_u7667_o;
  wire _al_u7668_o;
  wire _al_u7669_o;
  wire _al_u7670_o;
  wire _al_u7671_o;
  wire _al_u7672_o;
  wire _al_u7673_o;
  wire _al_u7674_o;
  wire _al_u7675_o;
  wire _al_u7676_o;
  wire _al_u7678_o;
  wire _al_u7679_o;
  wire _al_u7681_o;
  wire _al_u7682_o;
  wire _al_u7683_o;
  wire _al_u7685_o;
  wire _al_u7686_o;
  wire _al_u7688_o;
  wire _al_u7689_o;
  wire _al_u7691_o;
  wire _al_u7692_o;
  wire _al_u7693_o;
  wire _al_u7694_o;
  wire _al_u7695_o;
  wire _al_u7696_o;
  wire _al_u7697_o;
  wire _al_u7698_o;
  wire _al_u7699_o;
  wire _al_u7700_o;
  wire _al_u7701_o;
  wire _al_u7702_o;
  wire _al_u7704_o;
  wire _al_u7705_o;
  wire _al_u7707_o;
  wire _al_u7708_o;
  wire _al_u7710_o;
  wire _al_u7712_o;
  wire _al_u7713_o;
  wire _al_u7715_o;
  wire _al_u7716_o;
  wire _al_u7717_o;
  wire _al_u7718_o;
  wire _al_u7719_o;
  wire _al_u7720_o;
  wire _al_u7721_o;
  wire _al_u7722_o;
  wire _al_u7723_o;
  wire _al_u7724_o;
  wire _al_u7725_o;
  wire _al_u7726_o;
  wire _al_u7728_o;
  wire _al_u7729_o;
  wire _al_u7730_o;
  wire _al_u7731_o;
  wire _al_u7733_o;
  wire _al_u7734_o;
  wire _al_u7800_o;
  wire _al_u7801_o;
  wire _al_u7803_o;
  wire _al_u7804_o;
  wire _al_u7805_o;
  wire _al_u7806_o;
  wire _al_u7807_o;
  wire _al_u7808_o;
  wire _al_u7809_o;
  wire _al_u7810_o;
  wire _al_u7811_o;
  wire _al_u7812_o;
  wire _al_u7814_o;
  wire _al_u7816_o;
  wire _al_u7817_o;
  wire _al_u7819_o;
  wire _al_u7820_o;
  wire _al_u7822_o;
  wire _al_u7823_o;
  wire _al_u7825_o;
  wire _al_u7826_o;
  wire _al_u7828_o;
  wire _al_u7829_o;
  wire _al_u7831_o;
  wire _al_u7832_o;
  wire _al_u7834_o;
  wire _al_u7836_o;
  wire _al_u7838_o;
  wire _al_u7840_o;
  wire _al_u7842_o;
  wire _al_u7843_o;
  wire _al_u7845_o;
  wire _al_u7846_o;
  wire _al_u7848_o;
  wire _al_u7849_o;
  wire _al_u7851_o;
  wire _al_u7852_o;
  wire _al_u7854_o;
  wire _al_u7855_o;
  wire _al_u7857_o;
  wire _al_u7858_o;
  wire _al_u7859_o;
  wire _al_u7860_o;
  wire _al_u7861_o;
  wire _al_u7862_o;
  wire _al_u7863_o;
  wire _al_u7864_o;
  wire _al_u7865_o;
  wire _al_u7866_o;
  wire _al_u7867_o;
  wire _al_u7868_o;
  wire _al_u7869_o;
  wire _al_u7871_o;
  wire _al_u7873_o;
  wire _al_u7874_o;
  wire _al_u7875_o;
  wire _al_u7876_o;
  wire _al_u7877_o;
  wire _al_u7878_o;
  wire _al_u7879_o;
  wire _al_u7880_o;
  wire _al_u7881_o;
  wire _al_u7882_o;
  wire _al_u7883_o;
  wire _al_u7884_o;
  wire _al_u7885_o;
  wire _al_u7887_o;
  wire _al_u7889_o;
  wire _al_u7891_o;
  wire _al_u7893_o;
  wire _al_u7895_o;
  wire _al_u7897_o;
  wire _al_u7898_o;
  wire _al_u7899_o;
  wire _al_u7900_o;
  wire _al_u7901_o;
  wire _al_u7902_o;
  wire _al_u7905_o;
  wire _al_u7906_o;
  wire _al_u7907_o;
  wire _al_u7908_o;
  wire _al_u7909_o;
  wire _al_u7910_o;
  wire _al_u7911_o;
  wire _al_u7912_o;
  wire _al_u7913_o;
  wire _al_u7915_o;
  wire _al_u7916_o;
  wire _al_u7918_o;
  wire _al_u7919_o;
  wire _al_u7920_o;
  wire _al_u7921_o;
  wire _al_u7922_o;
  wire _al_u7923_o;
  wire _al_u7924_o;
  wire _al_u7925_o;
  wire _al_u7926_o;
  wire _al_u7927_o;
  wire _al_u7928_o;
  wire _al_u7930_o;
  wire _al_u7932_o;
  wire _al_u7933_o;
  wire _al_u7934_o;
  wire _al_u7935_o;
  wire _al_u7936_o;
  wire _al_u7937_o;
  wire _al_u7938_o;
  wire _al_u7939_o;
  wire _al_u7940_o;
  wire _al_u7941_o;
  wire _al_u7942_o;
  wire _al_u7943_o;
  wire _al_u7944_o;
  wire _al_u7945_o;
  wire _al_u7946_o;
  wire _al_u7947_o;
  wire _al_u7948_o;
  wire _al_u7949_o;
  wire _al_u7951_o;
  wire _al_u7953_o;
  wire _al_u7954_o;
  wire _al_u7955_o;
  wire _al_u7956_o;
  wire _al_u7957_o;
  wire _al_u7958_o;
  wire _al_u7959_o;
  wire _al_u7960_o;
  wire _al_u7961_o;
  wire _al_u7963_o;
  wire _al_u7965_o;
  wire _al_u7967_o;
  wire _al_u7968_o;
  wire _al_u7969_o;
  wire _al_u7970_o;
  wire _al_u7971_o;
  wire _al_u7973_o;
  wire _al_u7974_o;
  wire _al_u7975_o;
  wire _al_u7976_o;
  wire _al_u7977_o;
  wire _al_u7978_o;
  wire _al_u7979_o;
  wire _al_u7980_o;
  wire _al_u7981_o;
  wire _al_u7982_o;
  wire _al_u7985_o;
  wire _al_u7986_o;
  wire _al_u7987_o;
  wire _al_u7988_o;
  wire _al_u7990_o;
  wire _al_u7991_o;
  wire _al_u7993_o;
  wire _al_u7994_o;
  wire _al_u7995_o;
  wire _al_u7997_o;
  wire _al_u8000_o;
  wire _al_u8001_o;
  wire _al_u8002_o;
  wire _al_u8005_o;
  wire _al_u8007_o;
  wire _al_u8009_o;
  wire _al_u8011_o;
  wire _al_u8012_o;
  wire _al_u8013_o;
  wire _al_u8014_o;
  wire _al_u8016_o;
  wire _al_u8018_o;
  wire _al_u8019_o;
  wire _al_u8020_o;
  wire _al_u8022_o;
  wire _al_u8025_o;
  wire _al_u8027_o;
  wire _al_u8028_o;
  wire _al_u8029_o;
  wire _al_u8030_o;
  wire _al_u8031_o;
  wire _al_u8032_o;
  wire _al_u8034_o;
  wire _al_u8036_o;
  wire _al_u8037_o;
  wire _al_u8038_o;
  wire _al_u8040_o;
  wire _al_u8041_o;
  wire _al_u8042_o;
  wire _al_u8043_o;
  wire _al_u8045_o;
  wire _al_u8046_o;
  wire _al_u8047_o;
  wire _al_u8048_o;
  wire _al_u8050_o;
  wire _al_u8052_o;
  wire _al_u8053_o;
  wire _al_u8054_o;
  wire _al_u8056_o;
  wire _al_u8057_o;
  wire _al_u8058_o;
  wire _al_u8059_o;
  wire _al_u8061_o;
  wire _al_u8062_o;
  wire _al_u8063_o;
  wire _al_u8064_o;
  wire _al_u8066_o;
  wire _al_u8068_o;
  wire _al_u8069_o;
  wire _al_u8070_o;
  wire _al_u8072_o;
  wire _al_u8074_o;
  wire _al_u8075_o;
  wire _al_u8077_o;
  wire _al_u8078_o;
  wire _al_u8079_o;
  wire _al_u8080_o;
  wire _al_u8082_o;
  wire _al_u8084_o;
  wire _al_u8085_o;
  wire _al_u8086_o;
  wire _al_u8088_o;
  wire _al_u8090_o;
  wire _al_u8091_o;
  wire _al_u8093_o;
  wire _al_u8094_o;
  wire _al_u8095_o;
  wire _al_u8096_o;
  wire _al_u8098_o;
  wire _al_u8100_o;
  wire _al_u8101_o;
  wire _al_u8102_o;
  wire _al_u8104_o;
  wire _al_u8106_o;
  wire _al_u8107_o;
  wire _al_u8109_o;
  wire _al_u8110_o;
  wire _al_u8111_o;
  wire _al_u8112_o;
  wire _al_u8114_o;
  wire _al_u8116_o;
  wire _al_u8117_o;
  wire _al_u8118_o;
  wire _al_u8120_o;
  wire _al_u8122_o;
  wire _al_u8123_o;
  wire _al_u8125_o;
  wire _al_u8126_o;
  wire _al_u8127_o;
  wire _al_u8128_o;
  wire _al_u8129_o;
  wire _al_u8130_o;
  wire _al_u8131_o;
  wire _al_u8132_o;
  wire _al_u8133_o;
  wire _al_u8134_o;
  wire _al_u8136_o;
  wire _al_u8137_o;
  wire _al_u8138_o;
  wire _al_u8140_o;
  wire _al_u8142_o;
  wire _al_u8143_o;
  wire _al_u8145_o;
  wire _al_u8146_o;
  wire _al_u8147_o;
  wire _al_u8148_o;
  wire _al_u8149_o;
  wire _al_u8150_o;
  wire _al_u8151_o;
  wire _al_u8153_o;
  wire _al_u8154_o;
  wire _al_u8155_o;
  wire _al_u8157_o;
  wire _al_u8159_o;
  wire _al_u8160_o;
  wire _al_u8162_o;
  wire _al_u8163_o;
  wire _al_u8164_o;
  wire _al_u8165_o;
  wire _al_u8166_o;
  wire _al_u8167_o;
  wire _al_u8168_o;
  wire _al_u8169_o;
  wire _al_u8171_o;
  wire _al_u8172_o;
  wire _al_u8173_o;
  wire _al_u8175_o;
  wire _al_u8177_o;
  wire _al_u8178_o;
  wire _al_u8180_o;
  wire _al_u8181_o;
  wire _al_u8182_o;
  wire _al_u8183_o;
  wire _al_u8184_o;
  wire _al_u8185_o;
  wire _al_u8186_o;
  wire _al_u8188_o;
  wire _al_u8189_o;
  wire _al_u8190_o;
  wire _al_u8192_o;
  wire _al_u8194_o;
  wire _al_u8195_o;
  wire _al_u8197_o;
  wire _al_u8198_o;
  wire _al_u8199_o;
  wire _al_u8200_o;
  wire _al_u8201_o;
  wire _al_u8202_o;
  wire _al_u8203_o;
  wire _al_u8205_o;
  wire _al_u8206_o;
  wire _al_u8207_o;
  wire _al_u8209_o;
  wire _al_u8211_o;
  wire _al_u8212_o;
  wire _al_u8214_o;
  wire _al_u8215_o;
  wire _al_u8216_o;
  wire _al_u8217_o;
  wire _al_u8218_o;
  wire _al_u8219_o;
  wire _al_u8220_o;
  wire _al_u8222_o;
  wire _al_u8223_o;
  wire _al_u8224_o;
  wire _al_u8226_o;
  wire _al_u8228_o;
  wire _al_u8229_o;
  wire _al_u8231_o;
  wire _al_u8232_o;
  wire _al_u8233_o;
  wire _al_u8234_o;
  wire _al_u8235_o;
  wire _al_u8236_o;
  wire _al_u8237_o;
  wire _al_u8239_o;
  wire _al_u8240_o;
  wire _al_u8241_o;
  wire _al_u8243_o;
  wire _al_u8245_o;
  wire _al_u8246_o;
  wire _al_u8248_o;
  wire _al_u8249_o;
  wire _al_u8250_o;
  wire _al_u8251_o;
  wire _al_u8252_o;
  wire _al_u8253_o;
  wire _al_u8254_o;
  wire _al_u8256_o;
  wire _al_u8257_o;
  wire _al_u8258_o;
  wire _al_u8260_o;
  wire _al_u8262_o;
  wire _al_u8263_o;
  wire _al_u8265_o;
  wire _al_u8266_o;
  wire _al_u8267_o;
  wire _al_u8268_o;
  wire _al_u8269_o;
  wire _al_u8270_o;
  wire _al_u8271_o;
  wire _al_u8272_o;
  wire _al_u8274_o;
  wire _al_u8276_o;
  wire _al_u8277_o;
  wire _al_u8278_o;
  wire _al_u8280_o;
  wire _al_u8282_o;
  wire _al_u8283_o;
  wire _al_u8285_o;
  wire _al_u8286_o;
  wire _al_u8287_o;
  wire _al_u8288_o;
  wire _al_u8289_o;
  wire _al_u8290_o;
  wire _al_u8291_o;
  wire _al_u8293_o;
  wire _al_u8295_o;
  wire _al_u8296_o;
  wire _al_u8297_o;
  wire _al_u8299_o;
  wire _al_u8301_o;
  wire _al_u8302_o;
  wire _al_u8304_o;
  wire _al_u8305_o;
  wire _al_u8306_o;
  wire _al_u8307_o;
  wire _al_u8308_o;
  wire _al_u8309_o;
  wire _al_u8310_o;
  wire _al_u8311_o;
  wire _al_u8313_o;
  wire _al_u8315_o;
  wire _al_u8316_o;
  wire _al_u8317_o;
  wire _al_u8319_o;
  wire _al_u8321_o;
  wire _al_u8322_o;
  wire _al_u8324_o;
  wire _al_u8325_o;
  wire _al_u8326_o;
  wire _al_u8327_o;
  wire _al_u8328_o;
  wire _al_u8329_o;
  wire _al_u8330_o;
  wire _al_u8331_o;
  wire _al_u8333_o;
  wire _al_u8335_o;
  wire _al_u8336_o;
  wire _al_u8337_o;
  wire _al_u8339_o;
  wire _al_u8341_o;
  wire _al_u8342_o;
  wire _al_u8344_o;
  wire _al_u8345_o;
  wire _al_u8346_o;
  wire _al_u8347_o;
  wire _al_u8348_o;
  wire _al_u8349_o;
  wire _al_u8350_o;
  wire _al_u8352_o;
  wire _al_u8354_o;
  wire _al_u8355_o;
  wire _al_u8356_o;
  wire _al_u8358_o;
  wire _al_u8360_o;
  wire _al_u8361_o;
  wire _al_u8363_o;
  wire _al_u8364_o;
  wire _al_u8365_o;
  wire _al_u8366_o;
  wire _al_u8367_o;
  wire _al_u8368_o;
  wire _al_u8369_o;
  wire _al_u8371_o;
  wire _al_u8373_o;
  wire _al_u8374_o;
  wire _al_u8375_o;
  wire _al_u8377_o;
  wire _al_u8379_o;
  wire _al_u8380_o;
  wire _al_u8382_o;
  wire _al_u8383_o;
  wire _al_u8384_o;
  wire _al_u8385_o;
  wire _al_u8386_o;
  wire _al_u8387_o;
  wire _al_u8388_o;
  wire _al_u8390_o;
  wire _al_u8391_o;
  wire _al_u8392_o;
  wire _al_u8393_o;
  wire _al_u8395_o;
  wire _al_u8396_o;
  wire _al_u8397_o;
  wire _al_u8399_o;
  wire _al_u8401_o;
  wire _al_u8402_o;
  wire _al_u8403_o;
  wire _al_u8404_o;
  wire _al_u8405_o;
  wire _al_u8406_o;
  wire _al_u8407_o;
  wire _al_u8409_o;
  wire _al_u8410_o;
  wire _al_u8411_o;
  wire _al_u8412_o;
  wire _al_u8414_o;
  wire _al_u8415_o;
  wire _al_u8416_o;
  wire _al_u8418_o;
  wire _al_u8420_o;
  wire _al_u8421_o;
  wire _al_u8422_o;
  wire _al_u8423_o;
  wire _al_u8424_o;
  wire _al_u8425_o;
  wire _al_u8426_o;
  wire _al_u8427_o;
  wire _al_u8428_o;
  wire _al_u8429_o;
  wire _al_u8430_o;
  wire _al_u8431_o;
  wire _al_u8432_o;
  wire _al_u8433_o;
  wire _al_u8434_o;
  wire _al_u8436_o;
  wire _al_u8437_o;
  wire _al_u8438_o;
  wire _al_u8440_o;
  wire _al_u8442_o;
  wire _al_u8443_o;
  wire _al_u8444_o;
  wire _al_u8445_o;
  wire _al_u8446_o;
  wire _al_u8447_o;
  wire _al_u8448_o;
  wire _al_u8449_o;
  wire _al_u8450_o;
  wire _al_u8451_o;
  wire _al_u8452_o;
  wire _al_u8454_o;
  wire _al_u8455_o;
  wire _al_u8456_o;
  wire _al_u8458_o;
  wire _al_u8459_o;
  wire _al_u8460_o;
  wire _al_u8461_o;
  wire _al_u8463_o;
  wire _al_u8464_o;
  wire _al_u8465_o;
  wire _al_u8466_o;
  wire _al_u8467_o;
  wire _al_u8468_o;
  wire _al_u8469_o;
  wire _al_u8470_o;
  wire _al_u8471_o;
  wire _al_u8472_o;
  wire _al_u8473_o;
  wire _al_u8474_o;
  wire _al_u8476_o;
  wire _al_u8477_o;
  wire _al_u8478_o;
  wire _al_u8480_o;
  wire _al_u8481_o;
  wire _al_u8482_o;
  wire _al_u8483_o;
  wire _al_u8485_o;
  wire _al_u8486_o;
  wire _al_u8487_o;
  wire _al_u8488_o;
  wire _al_u8489_o;
  wire _al_u8490_o;
  wire _al_u8491_o;
  wire _al_u8492_o;
  wire _al_u8493_o;
  wire _al_u8494_o;
  wire _al_u8495_o;
  wire _al_u8496_o;
  wire _al_u8497_o;
  wire _al_u8499_o;
  wire _al_u8500_o;
  wire _al_u8501_o;
  wire _al_u8503_o;
  wire _al_u8505_o;
  wire _al_u8506_o;
  wire _al_u8508_o;
  wire _al_u8509_o;
  wire _al_u8510_o;
  wire _al_u8511_o;
  wire _al_u8512_o;
  wire _al_u8513_o;
  wire _al_u8514_o;
  wire _al_u8515_o;
  wire _al_u8516_o;
  wire _al_u8517_o;
  wire _al_u8518_o;
  wire _al_u8519_o;
  wire _al_u8520_o;
  wire _al_u8521_o;
  wire _al_u8523_o;
  wire _al_u8524_o;
  wire _al_u8525_o;
  wire _al_u8527_o;
  wire _al_u8529_o;
  wire _al_u8530_o;
  wire _al_u8531_o;
  wire _al_u8532_o;
  wire _al_u8533_o;
  wire _al_u8534_o;
  wire _al_u8535_o;
  wire _al_u8536_o;
  wire _al_u8537_o;
  wire _al_u8538_o;
  wire _al_u8539_o;
  wire _al_u8540_o;
  wire _al_u8541_o;
  wire _al_u8542_o;
  wire _al_u8544_o;
  wire _al_u8545_o;
  wire _al_u8546_o;
  wire _al_u8548_o;
  wire _al_u8550_o;
  wire _al_u8551_o;
  wire _al_u8552_o;
  wire _al_u8553_o;
  wire _al_u8554_o;
  wire _al_u8555_o;
  wire _al_u8556_o;
  wire _al_u8557_o;
  wire _al_u8558_o;
  wire _al_u8559_o;
  wire _al_u8561_o;
  wire _al_u8562_o;
  wire _al_u8563_o;
  wire _al_u8565_o;
  wire _al_u8567_o;
  wire _al_u8568_o;
  wire _al_u8570_o;
  wire _al_u8571_o;
  wire _al_u8572_o;
  wire _al_u8573_o;
  wire _al_u8574_o;
  wire _al_u8575_o;
  wire _al_u8576_o;
  wire _al_u8577_o;
  wire _al_u8578_o;
  wire _al_u8579_o;
  wire _al_u8581_o;
  wire _al_u8582_o;
  wire _al_u8583_o;
  wire _al_u8585_o;
  wire _al_u8587_o;
  wire _al_u8588_o;
  wire _al_u8590_o;
  wire _al_u8591_o;
  wire _al_u8592_o;
  wire _al_u8593_o;
  wire _al_u8594_o;
  wire _al_u8595_o;
  wire _al_u8596_o;
  wire _al_u8597_o;
  wire _al_u8598_o;
  wire _al_u8600_o;
  wire _al_u8601_o;
  wire _al_u8602_o;
  wire _al_u8603_o;
  wire _al_u8605_o;
  wire _al_u8606_o;
  wire _al_u8607_o;
  wire _al_u8608_o;
  wire _al_u8609_o;
  wire _al_u8610_o;
  wire _al_u8611_o;
  wire _al_u8612_o;
  wire _al_u8613_o;
  wire _al_u8614_o;
  wire _al_u8615_o;
  wire _al_u8616_o;
  wire _al_u8617_o;
  wire _al_u8618_o;
  wire _al_u8620_o;
  wire _al_u8622_o;
  wire _al_u8624_o;
  wire _al_u8625_o;
  wire _al_u8626_o;
  wire _al_u8627_o;
  wire _al_u8628_o;
  wire _al_u8629_o;
  wire _al_u8630_o;
  wire _al_u8631_o;
  wire _al_u8632_o;
  wire _al_u8633_o;
  wire _al_u8634_o;
  wire _al_u8635_o;
  wire _al_u8636_o;
  wire _al_u8637_o;
  wire _al_u8638_o;
  wire _al_u8640_o;
  wire _al_u8642_o;
  wire _al_u8644_o;
  wire _al_u8645_o;
  wire _al_u8646_o;
  wire _al_u8647_o;
  wire _al_u8648_o;
  wire _al_u8649_o;
  wire _al_u8650_o;
  wire _al_u8651_o;
  wire _al_u8652_o;
  wire _al_u8653_o;
  wire _al_u8654_o;
  wire _al_u8655_o;
  wire _al_u8656_o;
  wire _al_u8657_o;
  wire _al_u8658_o;
  wire _al_u8660_o;
  wire _al_u8662_o;
  wire _al_u8664_o;
  wire _al_u8665_o;
  wire _al_u8666_o;
  wire _al_u8667_o;
  wire _al_u8668_o;
  wire _al_u8669_o;
  wire _al_u8670_o;
  wire _al_u8671_o;
  wire _al_u8672_o;
  wire _al_u8673_o;
  wire _al_u8674_o;
  wire _al_u8675_o;
  wire _al_u8676_o;
  wire _al_u8677_o;
  wire _al_u8679_o;
  wire _al_u8681_o;
  wire _al_u8683_o;
  wire _al_u8684_o;
  wire _al_u8685_o;
  wire _al_u8686_o;
  wire _al_u8687_o;
  wire _al_u8688_o;
  wire _al_u8689_o;
  wire _al_u8690_o;
  wire _al_u8691_o;
  wire _al_u8692_o;
  wire _al_u8693_o;
  wire _al_u8694_o;
  wire _al_u8695_o;
  wire _al_u8696_o;
  wire _al_u8698_o;
  wire _al_u8700_o;
  wire _al_u8702_o;
  wire _al_u8703_o;
  wire _al_u8704_o;
  wire _al_u8705_o;
  wire _al_u8706_o;
  wire _al_u8707_o;
  wire _al_u8708_o;
  wire _al_u8709_o;
  wire _al_u8710_o;
  wire _al_u8711_o;
  wire _al_u8712_o;
  wire _al_u8713_o;
  wire _al_u8714_o;
  wire _al_u8716_o;
  wire _al_u8718_o;
  wire _al_u8720_o;
  wire _al_u8721_o;
  wire _al_u8722_o;
  wire _al_u8723_o;
  wire _al_u8724_o;
  wire _al_u8725_o;
  wire _al_u8726_o;
  wire _al_u8727_o;
  wire _al_u8728_o;
  wire _al_u8729_o;
  wire _al_u8730_o;
  wire _al_u8731_o;
  wire _al_u8732_o;
  wire _al_u8734_o;
  wire _al_u8736_o;
  wire _al_u8738_o;
  wire _al_u8739_o;
  wire _al_u8740_o;
  wire _al_u8741_o;
  wire _al_u8742_o;
  wire _al_u8743_o;
  wire _al_u8744_o;
  wire _al_u8745_o;
  wire _al_u8746_o;
  wire _al_u8747_o;
  wire _al_u8748_o;
  wire _al_u8749_o;
  wire _al_u8750_o;
  wire _al_u8751_o;
  wire _al_u8752_o;
  wire _al_u8753_o;
  wire _al_u8755_o;
  wire _al_u8757_o;
  wire _al_u8759_o;
  wire _al_u8760_o;
  wire _al_u8761_o;
  wire _al_u8762_o;
  wire _al_u8763_o;
  wire _al_u8764_o;
  wire _al_u8765_o;
  wire _al_u8766_o;
  wire _al_u8767_o;
  wire _al_u8768_o;
  wire _al_u8769_o;
  wire _al_u8770_o;
  wire _al_u8771_o;
  wire _al_u8772_o;
  wire _al_u8774_o;
  wire _al_u8776_o;
  wire _al_u8778_o;
  wire _al_u8779_o;
  wire _al_u8780_o;
  wire _al_u8781_o;
  wire _al_u8782_o;
  wire _al_u8783_o;
  wire _al_u8784_o;
  wire _al_u8785_o;
  wire _al_u8786_o;
  wire _al_u8787_o;
  wire _al_u8788_o;
  wire _al_u8789_o;
  wire _al_u8790_o;
  wire _al_u8791_o;
  wire _al_u8793_o;
  wire _al_u8795_o;
  wire _al_u8797_o;
  wire _al_u8798_o;
  wire _al_u8799_o;
  wire _al_u8800_o;
  wire _al_u8801_o;
  wire _al_u8802_o;
  wire _al_u8803_o;
  wire _al_u8804_o;
  wire _al_u8805_o;
  wire _al_u8806_o;
  wire _al_u8807_o;
  wire _al_u8808_o;
  wire _al_u8809_o;
  wire _al_u8810_o;
  wire _al_u8812_o;
  wire _al_u8814_o;
  wire _al_u8816_o;
  wire _al_u8817_o;
  wire _al_u8818_o;
  wire _al_u8819_o;
  wire _al_u8820_o;
  wire _al_u8821_o;
  wire _al_u8822_o;
  wire _al_u8823_o;
  wire _al_u8824_o;
  wire _al_u8825_o;
  wire _al_u8826_o;
  wire _al_u8827_o;
  wire _al_u8828_o;
  wire _al_u8829_o;
  wire _al_u8831_o;
  wire _al_u8833_o;
  wire _al_u8835_o;
  wire _al_u8836_o;
  wire _al_u8837_o;
  wire _al_u8838_o;
  wire _al_u8839_o;
  wire _al_u8840_o;
  wire _al_u8841_o;
  wire _al_u8842_o;
  wire _al_u8843_o;
  wire _al_u8844_o;
  wire _al_u8845_o;
  wire _al_u8846_o;
  wire _al_u8847_o;
  wire _al_u8848_o;
  wire _al_u8850_o;
  wire _al_u8852_o;
  wire _al_u8854_o;
  wire _al_u8855_o;
  wire _al_u8856_o;
  wire _al_u8857_o;
  wire _al_u8858_o;
  wire _al_u8859_o;
  wire _al_u8860_o;
  wire _al_u8861_o;
  wire _al_u8862_o;
  wire _al_u8863_o;
  wire _al_u8864_o;
  wire _al_u8865_o;
  wire _al_u8866_o;
  wire _al_u8868_o;
  wire _al_u8870_o;
  wire _al_u8872_o;
  wire _al_u8873_o;
  wire _al_u8874_o;
  wire _al_u8875_o;
  wire _al_u8876_o;
  wire _al_u8877_o;
  wire _al_u8878_o;
  wire _al_u8879_o;
  wire _al_u8880_o;
  wire _al_u8881_o;
  wire _al_u8882_o;
  wire _al_u8883_o;
  wire _al_u8884_o;
  wire _al_u8886_o;
  wire _al_u8888_o;
  wire _al_u8890_o;
  wire _al_u8891_o;
  wire _al_u8892_o;
  wire _al_u8893_o;
  wire _al_u8894_o;
  wire _al_u8895_o;
  wire _al_u8896_o;
  wire _al_u8897_o;
  wire _al_u8898_o;
  wire _al_u8900_o;
  wire _al_u8902_o;
  wire _al_u8904_o;
  wire _al_u8905_o;
  wire _al_u8906_o;
  wire _al_u8907_o;
  wire _al_u8908_o;
  wire _al_u8909_o;
  wire _al_u8910_o;
  wire _al_u8911_o;
  wire _al_u8912_o;
  wire _al_u8913_o;
  wire _al_u8914_o;
  wire _al_u8915_o;
  wire _al_u8916_o;
  wire _al_u8918_o;
  wire _al_u8920_o;
  wire _al_u8922_o;
  wire _al_u8923_o;
  wire _al_u8924_o;
  wire _al_u8925_o;
  wire _al_u8926_o;
  wire _al_u8927_o;
  wire _al_u8928_o;
  wire _al_u8929_o;
  wire _al_u8930_o;
  wire _al_u8931_o;
  wire _al_u8932_o;
  wire _al_u8933_o;
  wire _al_u8934_o;
  wire _al_u8935_o;
  wire _al_u8937_o;
  wire _al_u8939_o;
  wire _al_u8940_o;
  wire _al_u8941_o;
  wire _al_u8942_o;
  wire _al_u8943_o;
  wire _al_u8944_o;
  wire _al_u8945_o;
  wire _al_u8946_o;
  wire _al_u8947_o;
  wire _al_u8948_o;
  wire _al_u8949_o;
  wire _al_u8950_o;
  wire _al_u8951_o;
  wire _al_u8952_o;
  wire _al_u8953_o;
  wire _al_u8955_o;
  wire _al_u8957_o;
  wire _al_u8959_o;
  wire _al_u8960_o;
  wire _al_u8961_o;
  wire _al_u8962_o;
  wire _al_u8963_o;
  wire _al_u8964_o;
  wire _al_u8965_o;
  wire _al_u8966_o;
  wire _al_u8967_o;
  wire _al_u8968_o;
  wire _al_u8969_o;
  wire _al_u8970_o;
  wire _al_u8971_o;
  wire _al_u8972_o;
  wire _al_u8974_o;
  wire _al_u8976_o;
  wire _al_u8977_o;
  wire _al_u8978_o;
  wire _al_u8979_o;
  wire _al_u8980_o;
  wire _al_u8981_o;
  wire _al_u8982_o;
  wire _al_u8983_o;
  wire _al_u8984_o;
  wire _al_u8985_o;
  wire _al_u8986_o;
  wire _al_u8987_o;
  wire _al_u8988_o;
  wire _al_u8990_o;
  wire _al_u8992_o;
  wire _al_u8994_o;
  wire _al_u8995_o;
  wire _al_u8996_o;
  wire _al_u8997_o;
  wire _al_u8998_o;
  wire _al_u8999_o;
  wire _al_u9000_o;
  wire _al_u9001_o;
  wire _al_u9002_o;
  wire _al_u9003_o;
  wire _al_u9004_o;
  wire _al_u9005_o;
  wire _al_u9006_o;
  wire _al_u9007_o;
  wire _al_u9009_o;
  wire _al_u9011_o;
  wire _al_u9012_o;
  wire _al_u9013_o;
  wire _al_u9014_o;
  wire _al_u9015_o;
  wire _al_u9016_o;
  wire _al_u9017_o;
  wire _al_u9018_o;
  wire _al_u9019_o;
  wire _al_u9020_o;
  wire _al_u9021_o;
  wire _al_u9022_o;
  wire _al_u9023_o;
  wire _al_u9025_o;
  wire _al_u9027_o;
  wire _al_u9029_o;
  wire _al_u9030_o;
  wire _al_u9031_o;
  wire _al_u9032_o;
  wire _al_u9033_o;
  wire _al_u9034_o;
  wire _al_u9035_o;
  wire _al_u9036_o;
  wire _al_u9037_o;
  wire _al_u9038_o;
  wire _al_u9039_o;
  wire _al_u9040_o;
  wire _al_u9041_o;
  wire _al_u9042_o;
  wire _al_u9044_o;
  wire _al_u9046_o;
  wire _al_u9047_o;
  wire _al_u9048_o;
  wire _al_u9049_o;
  wire _al_u9050_o;
  wire _al_u9051_o;
  wire _al_u9052_o;
  wire _al_u9053_o;
  wire _al_u9054_o;
  wire _al_u9055_o;
  wire _al_u9056_o;
  wire _al_u9057_o;
  wire _al_u9058_o;
  wire _al_u9059_o;
  wire _al_u9060_o;
  wire _al_u9062_o;
  wire _al_u9064_o;
  wire _al_u9066_o;
  wire _al_u9067_o;
  wire _al_u9068_o;
  wire _al_u9069_o;
  wire _al_u9070_o;
  wire _al_u9071_o;
  wire _al_u9072_o;
  wire _al_u9073_o;
  wire _al_u9074_o;
  wire _al_u9075_o;
  wire _al_u9076_o;
  wire _al_u9077_o;
  wire _al_u9078_o;
  wire _al_u9079_o;
  wire _al_u9081_o;
  wire _al_u9083_o;
  wire _al_u9084_o;
  wire _al_u9085_o;
  wire _al_u9086_o;
  wire _al_u9087_o;
  wire _al_u9088_o;
  wire _al_u9089_o;
  wire _al_u9090_o;
  wire _al_u9091_o;
  wire _al_u9092_o;
  wire _al_u9093_o;
  wire _al_u9094_o;
  wire _al_u9095_o;
  wire _al_u9096_o;
  wire _al_u9098_o;
  wire _al_u9100_o;
  wire _al_u9102_o;
  wire _al_u9103_o;
  wire _al_u9104_o;
  wire _al_u9105_o;
  wire _al_u9106_o;
  wire _al_u9107_o;
  wire _al_u9108_o;
  wire _al_u9110_o;
  wire _al_u9111_o;
  wire _al_u9112_o;
  wire _al_u9113_o;
  wire _al_u9114_o;
  wire _al_u9117_o;
  wire _al_u9118_o;
  wire _al_u9119_o;
  wire _al_u9121_o;
  wire _al_u9122_o;
  wire _al_u9125_o;
  wire _al_u9126_o;
  wire _al_u9127_o;
  wire _al_u9128_o;
  wire _al_u9129_o;
  wire _al_u9130_o;
  wire _al_u9131_o;
  wire _al_u9133_o;
  wire _al_u9134_o;
  wire _al_u9135_o;
  wire _al_u9137_o;
  wire _al_u9139_o;
  wire _al_u9141_o;
  wire _al_u9142_o;
  wire _al_u9144_o;
  wire _al_u9146_o;
  wire _al_u9147_o;
  wire _al_u9148_o;
  wire _al_u9149_o;
  wire _al_u9151_o;
  wire _al_u9152_o;
  wire _al_u9153_o;
  wire _al_u9154_o;
  wire _al_u9155_o;
  wire _al_u9156_o;
  wire _al_u9158_o;
  wire _al_u9159_o;
  wire _al_u9160_o;
  wire _al_u9161_o;
  wire _al_u9162_o;
  wire _al_u9164_o;
  wire _al_u9165_o;
  wire _al_u9166_o;
  wire _al_u9167_o;
  wire _al_u9168_o;
  wire _al_u9170_o;
  wire _al_u9171_o;
  wire _al_u9173_o;
  wire _al_u9174_o;
  wire _al_u9175_o;
  wire _al_u9176_o;
  wire _al_u9177_o;
  wire _al_u9178_o;
  wire _al_u9179_o;
  wire _al_u9180_o;
  wire _al_u9181_o;
  wire _al_u9182_o;
  wire _al_u9183_o;
  wire _al_u9184_o;
  wire _al_u9186_o;
  wire _al_u9188_o;
  wire _al_u9189_o;
  wire _al_u9190_o;
  wire _al_u9192_o;
  wire _al_u9193_o;
  wire _al_u9195_o;
  wire _al_u9197_o;
  wire _al_u9204_o;
  wire _al_u9205_o;
  wire _al_u9206_o;
  wire _al_u9207_o;
  wire _al_u9208_o;
  wire _al_u9209_o;
  wire _al_u9210_o;
  wire _al_u9211_o;
  wire _al_u9212_o;
  wire _al_u9213_o;
  wire _al_u9214_o;
  wire _al_u9215_o;
  wire _al_u9216_o;
  wire _al_u9217_o;
  wire _al_u9218_o;
  wire _al_u9219_o;
  wire _al_u9220_o;
  wire _al_u9221_o;
  wire _al_u9222_o;
  wire _al_u9223_o;
  wire _al_u9224_o;
  wire _al_u9225_o;
  wire _al_u9226_o;
  wire _al_u9227_o;
  wire _al_u9228_o;
  wire _al_u9229_o;
  wire _al_u9230_o;
  wire _al_u9231_o;
  wire _al_u9232_o;
  wire _al_u9233_o;
  wire _al_u9234_o;
  wire _al_u9235_o;
  wire _al_u9236_o;
  wire _al_u9237_o;
  wire _al_u9238_o;
  wire _al_u9239_o;
  wire _al_u9240_o;
  wire _al_u9241_o;
  wire _al_u9242_o;
  wire _al_u9243_o;
  wire _al_u9244_o;
  wire _al_u9245_o;
  wire _al_u9246_o;
  wire _al_u9247_o;
  wire _al_u9248_o;
  wire _al_u9249_o;
  wire _al_u9250_o;
  wire _al_u9251_o;
  wire _al_u9252_o;
  wire _al_u9253_o;
  wire _al_u9254_o;
  wire _al_u9255_o;
  wire _al_u9256_o;
  wire _al_u9257_o;
  wire _al_u9258_o;
  wire _al_u9259_o;
  wire _al_u9260_o;
  wire _al_u9261_o;
  wire _al_u9262_o;
  wire _al_u9263_o;
  wire _al_u9264_o;
  wire _al_u9265_o;
  wire _al_u9266_o;
  wire _al_u9268_o;
  wire _al_u9270_o;
  wire _al_u9271_o;
  wire _al_u9272_o;
  wire _al_u9273_o;
  wire _al_u9274_o;
  wire _al_u9275_o;
  wire _al_u9276_o;
  wire _al_u9277_o;
  wire _al_u9278_o;
  wire _al_u9279_o;
  wire _al_u9280_o;
  wire _al_u9281_o;
  wire _al_u9283_o;
  wire _al_u9284_o;
  wire _al_u9285_o;
  wire _al_u9286_o;
  wire _al_u9287_o;
  wire _al_u9289_o;
  wire _al_u9290_o;
  wire _al_u9292_o;
  wire _al_u9293_o;
  wire _al_u9294_o;
  wire _al_u9296_o;
  wire _al_u9297_o;
  wire _al_u9298_o;
  wire _al_u9299_o;
  wire _al_u9301_o;
  wire _al_u9302_o;
  wire _al_u9303_o;
  wire _al_u9304_o;
  wire _al_u9306_o;
  wire _al_u9307_o;
  wire _al_u9308_o;
  wire _al_u9309_o;
  wire _al_u9311_o;
  wire _al_u9312_o;
  wire _al_u9313_o;
  wire _al_u9315_o;
  wire _al_u9316_o;
  wire _al_u9317_o;
  wire _al_u9318_o;
  wire _al_u9320_o;
  wire _al_u9321_o;
  wire _al_u9322_o;
  wire _al_u9323_o;
  wire _al_u9325_o;
  wire _al_u9326_o;
  wire _al_u9327_o;
  wire _al_u9328_o;
  wire _al_u9330_o;
  wire _al_u9331_o;
  wire _al_u9332_o;
  wire _al_u9333_o;
  wire _al_u9335_o;
  wire _al_u9336_o;
  wire _al_u9337_o;
  wire _al_u9338_o;
  wire _al_u9340_o;
  wire _al_u9341_o;
  wire _al_u9342_o;
  wire _al_u9343_o;
  wire _al_u9345_o;
  wire _al_u9346_o;
  wire _al_u9347_o;
  wire _al_u9348_o;
  wire _al_u9349_o;
  wire _al_u9350_o;
  wire _al_u9352_o;
  wire _al_u9353_o;
  wire _al_u9354_o;
  wire _al_u9355_o;
  wire _al_u9356_o;
  wire _al_u9357_o;
  wire _al_u9359_o;
  wire _al_u9360_o;
  wire _al_u9361_o;
  wire _al_u9362_o;
  wire _al_u9363_o;
  wire _al_u9364_o;
  wire _al_u9366_o;
  wire _al_u9367_o;
  wire _al_u9368_o;
  wire _al_u9369_o;
  wire _al_u9371_o;
  wire _al_u9372_o;
  wire _al_u9373_o;
  wire _al_u9374_o;
  wire _al_u9375_o;
  wire _al_u9376_o;
  wire _al_u9378_o;
  wire _al_u9379_o;
  wire _al_u9380_o;
  wire _al_u9381_o;
  wire _al_u9382_o;
  wire _al_u9383_o;
  wire _al_u9385_o;
  wire _al_u9386_o;
  wire _al_u9387_o;
  wire _al_u9388_o;
  wire _al_u9389_o;
  wire _al_u9390_o;
  wire _al_u9392_o;
  wire _al_u9393_o;
  wire _al_u9394_o;
  wire _al_u9395_o;
  wire _al_u9396_o;
  wire _al_u9397_o;
  wire _al_u9399_o;
  wire _al_u9400_o;
  wire _al_u9401_o;
  wire _al_u9402_o;
  wire _al_u9404_o;
  wire _al_u9405_o;
  wire _al_u9406_o;
  wire _al_u9407_o;
  wire _al_u9408_o;
  wire _al_u9409_o;
  wire _al_u9411_o;
  wire _al_u9412_o;
  wire _al_u9413_o;
  wire _al_u9414_o;
  wire _al_u9415_o;
  wire _al_u9416_o;
  wire _al_u9418_o;
  wire _al_u9419_o;
  wire _al_u9420_o;
  wire _al_u9421_o;
  wire _al_u9422_o;
  wire _al_u9423_o;
  wire _al_u9425_o;
  wire _al_u9426_o;
  wire _al_u9427_o;
  wire _al_u9428_o;
  wire _al_u9430_o;
  wire _al_u9431_o;
  wire _al_u9432_o;
  wire _al_u9433_o;
  wire _al_u9434_o;
  wire _al_u9435_o;
  wire _al_u9437_o;
  wire _al_u9438_o;
  wire _al_u9439_o;
  wire _al_u9440_o;
  wire _al_u9441_o;
  wire _al_u9442_o;
  wire _al_u9444_o;
  wire _al_u9445_o;
  wire _al_u9446_o;
  wire _al_u9447_o;
  wire _al_u9449_o;
  wire _al_u9450_o;
  wire _al_u9451_o;
  wire _al_u9452_o;
  wire _al_u9453_o;
  wire _al_u9454_o;
  wire _al_u9456_o;
  wire _al_u9457_o;
  wire _al_u9458_o;
  wire _al_u9459_o;
  wire _al_u9461_o;
  wire _al_u9462_o;
  wire _al_u9463_o;
  wire _al_u9464_o;
  wire _al_u9465_o;
  wire _al_u9466_o;
  wire _al_u9468_o;
  wire _al_u9469_o;
  wire _al_u9470_o;
  wire _al_u9471_o;
  wire _al_u9473_o;
  wire _al_u9474_o;
  wire _al_u9475_o;
  wire _al_u9476_o;
  wire _al_u9477_o;
  wire _al_u9478_o;
  wire _al_u9480_o;
  wire _al_u9481_o;
  wire _al_u9482_o;
  wire _al_u9483_o;
  wire _al_u9484_o;
  wire _al_u9485_o;
  wire _al_u9487_o;
  wire _al_u9488_o;
  wire _al_u9489_o;
  wire _al_u9490_o;
  wire _al_u9491_o;
  wire _al_u9492_o;
  wire _al_u9494_o;
  wire _al_u9495_o;
  wire _al_u9496_o;
  wire _al_u9497_o;
  wire _al_u9499_o;
  wire _al_u9500_o;
  wire _al_u9501_o;
  wire _al_u9502_o;
  wire _al_u9503_o;
  wire _al_u9504_o;
  wire _al_u9506_o;
  wire _al_u9507_o;
  wire _al_u9508_o;
  wire _al_u9509_o;
  wire _al_u9510_o;
  wire _al_u9511_o;
  wire _al_u9513_o;
  wire _al_u9514_o;
  wire _al_u9515_o;
  wire _al_u9516_o;
  wire _al_u9518_o;
  wire _al_u9519_o;
  wire _al_u9520_o;
  wire _al_u9521_o;
  wire _al_u9522_o;
  wire _al_u9523_o;
  wire _al_u9525_o;
  wire _al_u9526_o;
  wire _al_u9527_o;
  wire _al_u9528_o;
  wire _al_u9530_o;
  wire _al_u9531_o;
  wire _al_u9532_o;
  wire _al_u9533_o;
  wire _al_u9534_o;
  wire _al_u9535_o;
  wire _al_u9537_o;
  wire _al_u9538_o;
  wire _al_u9539_o;
  wire _al_u9540_o;
  wire _al_u9541_o;
  wire _al_u9542_o;
  wire _al_u9544_o;
  wire _al_u9545_o;
  wire _al_u9546_o;
  wire _al_u9547_o;
  wire _al_u9548_o;
  wire _al_u9549_o;
  wire _al_u9551_o;
  wire _al_u9552_o;
  wire _al_u9553_o;
  wire _al_u9554_o;
  wire _al_u9555_o;
  wire _al_u9556_o;
  wire _al_u9558_o;
  wire _al_u9559_o;
  wire _al_u9560_o;
  wire _al_u9561_o;
  wire _al_u9562_o;
  wire _al_u9563_o;
  wire _al_u9565_o;
  wire _al_u9566_o;
  wire _al_u9567_o;
  wire _al_u9568_o;
  wire _al_u9569_o;
  wire _al_u9570_o;
  wire _al_u9572_o;
  wire _al_u9573_o;
  wire _al_u9574_o;
  wire _al_u9575_o;
  wire _al_u9576_o;
  wire _al_u9577_o;
  wire _al_u9579_o;
  wire _al_u9580_o;
  wire _al_u9581_o;
  wire _al_u9582_o;
  wire _al_u9583_o;
  wire _al_u9584_o;
  wire _al_u9586_o;
  wire _al_u9587_o;
  wire _al_u9588_o;
  wire _al_u9589_o;
  wire _al_u9591_o;
  wire _al_u9592_o;
  wire _al_u9593_o;
  wire _al_u9594_o;
  wire _al_u9595_o;
  wire _al_u9596_o;
  wire _al_u9598_o;
  wire _al_u9599_o;
  wire _al_u9600_o;
  wire _al_u9601_o;
  wire _al_u9602_o;
  wire _al_u9603_o;
  wire _al_u9605_o;
  wire _al_u9606_o;
  wire _al_u9607_o;
  wire _al_u9608_o;
  wire _al_u9609_o;
  wire _al_u9610_o;
  wire _al_u9612_o;
  wire _al_u9613_o;
  wire _al_u9614_o;
  wire _al_u9615_o;
  wire _al_u9616_o;
  wire _al_u9617_o;
  wire _al_u9619_o;
  wire _al_u9620_o;
  wire _al_u9621_o;
  wire _al_u9622_o;
  wire _al_u9624_o;
  wire _al_u9625_o;
  wire _al_u9626_o;
  wire _al_u9627_o;
  wire _al_u9628_o;
  wire _al_u9629_o;
  wire _al_u9631_o;
  wire _al_u9632_o;
  wire _al_u9633_o;
  wire _al_u9634_o;
  wire _al_u9635_o;
  wire _al_u9636_o;
  wire _al_u9638_o;
  wire _al_u9639_o;
  wire _al_u9640_o;
  wire _al_u9641_o;
  wire _al_u9642_o;
  wire _al_u9643_o;
  wire _al_u9645_o;
  wire _al_u9646_o;
  wire _al_u9647_o;
  wire _al_u9648_o;
  wire _al_u9650_o;
  wire _al_u9651_o;
  wire _al_u9652_o;
  wire _al_u9653_o;
  wire _al_u9654_o;
  wire _al_u9655_o;
  wire _al_u9657_o;
  wire _al_u9658_o;
  wire _al_u9659_o;
  wire _al_u9660_o;
  wire _al_u9661_o;
  wire _al_u9662_o;
  wire _al_u9664_o;
  wire _al_u9665_o;
  wire _al_u9666_o;
  wire _al_u9667_o;
  wire _al_u9669_o;
  wire _al_u9670_o;
  wire _al_u9671_o;
  wire _al_u9672_o;
  wire _al_u9673_o;
  wire _al_u9674_o;
  wire _al_u9676_o;
  wire _al_u9677_o;
  wire _al_u9678_o;
  wire _al_u9679_o;
  wire _al_u9680_o;
  wire _al_u9681_o;
  wire _al_u9682_o;
  wire _al_u9683_o;
  wire _al_u9685_o;
  wire _al_u9686_o;
  wire _al_u9687_o;
  wire _al_u9688_o;
  wire _al_u9689_o;
  wire _al_u9690_o;
  wire _al_u9691_o;
  wire _al_u9692_o;
  wire _al_u9693_o;
  wire _al_u9695_o;
  wire _al_u9696_o;
  wire _al_u9697_o;
  wire _al_u9698_o;
  wire _al_u9699_o;
  wire _al_u9700_o;
  wire _al_u9701_o;
  wire _al_u9702_o;
  wire _al_u9704_o;
  wire _al_u9705_o;
  wire _al_u9706_o;
  wire _al_u9707_o;
  wire _al_u9708_o;
  wire _al_u9709_o;
  wire _al_u9710_o;
  wire _al_u9711_o;
  wire _al_u9712_o;
  wire _al_u9713_o;
  wire amo;  // ../../RTL/CPU/prv464_top.v(138)
  wire and_clr;  // ../../RTL/CPU/prv464_top.v(129)
  wire \biu/bus_unit/add0/c1 ;
  wire \biu/bus_unit/add0/c3 ;
  wire \biu/bus_unit/add0/c5 ;
  wire \biu/bus_unit/add0/c7 ;
  wire \biu/bus_unit/add1/c1 ;
  wire \biu/bus_unit/add1/c11 ;
  wire \biu/bus_unit/add1/c13 ;
  wire \biu/bus_unit/add1/c15 ;
  wire \biu/bus_unit/add1/c17 ;
  wire \biu/bus_unit/add1/c19 ;
  wire \biu/bus_unit/add1/c21 ;
  wire \biu/bus_unit/add1/c23 ;
  wire \biu/bus_unit/add1/c25 ;
  wire \biu/bus_unit/add1/c27 ;
  wire \biu/bus_unit/add1/c29 ;
  wire \biu/bus_unit/add1/c3 ;
  wire \biu/bus_unit/add1/c31 ;
  wire \biu/bus_unit/add1/c33 ;
  wire \biu/bus_unit/add1/c35 ;
  wire \biu/bus_unit/add1/c37 ;
  wire \biu/bus_unit/add1/c39 ;
  wire \biu/bus_unit/add1/c41 ;
  wire \biu/bus_unit/add1/c43 ;
  wire \biu/bus_unit/add1/c45 ;
  wire \biu/bus_unit/add1/c47 ;
  wire \biu/bus_unit/add1/c49 ;
  wire \biu/bus_unit/add1/c5 ;
  wire \biu/bus_unit/add1/c51 ;
  wire \biu/bus_unit/add1/c53 ;
  wire \biu/bus_unit/add1/c55 ;
  wire \biu/bus_unit/add1/c57 ;
  wire \biu/bus_unit/add1/c59 ;
  wire \biu/bus_unit/add1/c7 ;
  wire \biu/bus_unit/add1/c9 ;
  wire \biu/bus_unit/mmu/mux10_b0_sel_is_2_o ;
  wire \biu/bus_unit/mmu/mux18_b3_sel_is_2_o ;
  wire \biu/bus_unit/mmu/mux20_b0_sel_is_3_o ;
  wire \biu/bus_unit/mmu/mux24_b0_sel_is_1_o ;
  wire \biu/bus_unit/mmu/mux34_b0_sel_is_3_o ;
  wire \biu/bus_unit/mmu/n12_lutinv ;
  wire \biu/bus_unit/mmu/n19_lutinv ;
  wire \biu/bus_unit/mmu/n2 ;
  wire \biu/bus_unit/mmu/n31_lutinv ;
  wire \biu/bus_unit/mmu/n37_lutinv ;
  wire \biu/bus_unit/mmu/n45_lutinv ;
  wire \biu/bus_unit/mmu/n58 ;
  wire \biu/bus_unit/mmu/n7_lutinv ;
  wire \biu/bus_unit/mmu/n8_lutinv ;
  wire \biu/bus_unit/mux10_b3_sel_is_0_o ;
  wire \biu/bus_unit/mux11_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux15_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux17_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux1_b1_sel_is_0_o ;
  wire \biu/bus_unit/n15_lutinv ;
  wire \biu/bus_unit/n37 ;
  wire \biu/bus_unit/n39[0]_en ;
  wire \biu/bus_unit/n45_lutinv ;
  wire \biu/bus_unit/sub0/c1 ;
  wire \biu/bus_unit/sub0/c3 ;
  wire \biu/bus_unit/sub0/c5 ;
  wire \biu/bus_unit/sub0/c7 ;
  wire \biu/cache/n1 ;
  wire \biu/cache/n11 ;
  wire \biu/cache/n13 ;
  wire \biu/cache/n15 ;
  wire \biu/cache/n17 ;
  wire \biu/cache/n19 ;
  wire \biu/cache/n21 ;
  wire \biu/cache/n23 ;
  wire \biu/cache/n25 ;
  wire \biu/cache/n27 ;
  wire \biu/cache/n29 ;
  wire \biu/cache/n3 ;
  wire \biu/cache/n31 ;
  wire \biu/cache/n5 ;
  wire \biu/cache/n7 ;
  wire \biu/cache/n9 ;
  wire \biu/cache_ctrl_logic/add0/c11 ;
  wire \biu/cache_ctrl_logic/add0/c15 ;
  wire \biu/cache_ctrl_logic/add0/c19 ;
  wire \biu/cache_ctrl_logic/add0/c23 ;
  wire \biu/cache_ctrl_logic/add0/c27 ;
  wire \biu/cache_ctrl_logic/add0/c3 ;
  wire \biu/cache_ctrl_logic/add0/c31 ;
  wire \biu/cache_ctrl_logic/add0/c35 ;
  wire \biu/cache_ctrl_logic/add0/c39 ;
  wire \biu/cache_ctrl_logic/add0/c43 ;
  wire \biu/cache_ctrl_logic/add0/c47 ;
  wire \biu/cache_ctrl_logic/add0/c51 ;
  wire \biu/cache_ctrl_logic/add0/c55 ;
  wire \biu/cache_ctrl_logic/add0/c59 ;
  wire \biu/cache_ctrl_logic/add0/c63 ;
  wire \biu/cache_ctrl_logic/add0/c7 ;
  wire \biu/cache_ctrl_logic/add1/c11 ;
  wire \biu/cache_ctrl_logic/add1/c15 ;
  wire \biu/cache_ctrl_logic/add1/c19 ;
  wire \biu/cache_ctrl_logic/add1/c23 ;
  wire \biu/cache_ctrl_logic/add1/c27 ;
  wire \biu/cache_ctrl_logic/add1/c3 ;
  wire \biu/cache_ctrl_logic/add1/c31 ;
  wire \biu/cache_ctrl_logic/add1/c35 ;
  wire \biu/cache_ctrl_logic/add1/c39 ;
  wire \biu/cache_ctrl_logic/add1/c43 ;
  wire \biu/cache_ctrl_logic/add1/c47 ;
  wire \biu/cache_ctrl_logic/add1/c51 ;
  wire \biu/cache_ctrl_logic/add1/c55 ;
  wire \biu/cache_ctrl_logic/add1/c59 ;
  wire \biu/cache_ctrl_logic/add1/c63 ;
  wire \biu/cache_ctrl_logic/add1/c7 ;
  wire \biu/cache_ctrl_logic/add2/c11 ;
  wire \biu/cache_ctrl_logic/add2/c15 ;
  wire \biu/cache_ctrl_logic/add2/c19 ;
  wire \biu/cache_ctrl_logic/add2/c23 ;
  wire \biu/cache_ctrl_logic/add2/c27 ;
  wire \biu/cache_ctrl_logic/add2/c3 ;
  wire \biu/cache_ctrl_logic/add2/c31 ;
  wire \biu/cache_ctrl_logic/add2/c35 ;
  wire \biu/cache_ctrl_logic/add2/c39 ;
  wire \biu/cache_ctrl_logic/add2/c43 ;
  wire \biu/cache_ctrl_logic/add2/c47 ;
  wire \biu/cache_ctrl_logic/add2/c51 ;
  wire \biu/cache_ctrl_logic/add2/c55 ;
  wire \biu/cache_ctrl_logic/add2/c59 ;
  wire \biu/cache_ctrl_logic/add2/c63 ;
  wire \biu/cache_ctrl_logic/add2/c7 ;
  wire \biu/cache_ctrl_logic/eq1/xor_i0[4]_i1[4]_o_lutinv ;
  wire \biu/cache_ctrl_logic/ex_l1i_hit ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(155)
  wire \biu/cache_ctrl_logic/l1d_value ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(138)
  wire \biu/cache_ctrl_logic/l1d_wr_sel_lutinv ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(435)
  wire \biu/cache_ctrl_logic/l1i_value ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(137)
  wire \biu/cache_ctrl_logic/mux31_b4_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux44_b4_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/n135 ;
  wire \biu/cache_ctrl_logic/n140 ;
  wire \biu/cache_ctrl_logic/n149 ;
  wire \biu/cache_ctrl_logic/n17 ;
  wire \biu/cache_ctrl_logic/n172_lutinv ;
  wire \biu/cache_ctrl_logic/n173_lutinv ;
  wire \biu/cache_ctrl_logic/n174_lutinv ;
  wire \biu/cache_ctrl_logic/n176_lutinv ;
  wire \biu/cache_ctrl_logic/n204_lutinv ;
  wire \biu/cache_ctrl_logic/n26_lutinv ;
  wire \biu/cache_ctrl_logic/n30 ;
  wire \biu/cache_ctrl_logic/n34 ;
  wire \biu/cache_ctrl_logic/n36 ;
  wire \biu/cache_ctrl_logic/n40 ;
  wire \biu/cache_ctrl_logic/n42 ;
  wire \biu/cache_ctrl_logic/n55_lutinv ;
  wire \biu/cache_ctrl_logic/n75_lutinv ;
  wire \biu/cache_ctrl_logic/n97_lutinv ;
  wire \biu/cache_ctrl_logic/u128_sel_is_0_o ;
  wire \biu/cache_write_lutinv ;  // ../../RTL/CPU/BIU/biu.v(115)
  wire \biu/cacheable ;  // ../../RTL/CPU/BIU/biu.v(113)
  wire \biu/l1i_write_lutinv ;  // ../../RTL/CPU/BIU/biu.v(83)
  wire cache_flush;  // ../../RTL/CPU/prv464_top.v(139)
  wire cache_reset;  // ../../RTL/CPU/prv464_top.v(140)
  wire clk_pad;  // ../../RTL/CPU/prv464_top.v(19)
  wire \cu_ru/add0_2/c1 ;
  wire \cu_ru/add0_2/c11 ;
  wire \cu_ru/add0_2/c13 ;
  wire \cu_ru/add0_2/c15 ;
  wire \cu_ru/add0_2/c17 ;
  wire \cu_ru/add0_2/c19 ;
  wire \cu_ru/add0_2/c21 ;
  wire \cu_ru/add0_2/c23 ;
  wire \cu_ru/add0_2/c25 ;
  wire \cu_ru/add0_2/c27 ;
  wire \cu_ru/add0_2/c29 ;
  wire \cu_ru/add0_2/c3 ;
  wire \cu_ru/add0_2/c31 ;
  wire \cu_ru/add0_2/c33 ;
  wire \cu_ru/add0_2/c35 ;
  wire \cu_ru/add0_2/c37 ;
  wire \cu_ru/add0_2/c39 ;
  wire \cu_ru/add0_2/c41 ;
  wire \cu_ru/add0_2/c43 ;
  wire \cu_ru/add0_2/c45 ;
  wire \cu_ru/add0_2/c47 ;
  wire \cu_ru/add0_2/c49 ;
  wire \cu_ru/add0_2/c5 ;
  wire \cu_ru/add0_2/c51 ;
  wire \cu_ru/add0_2/c53 ;
  wire \cu_ru/add0_2/c55 ;
  wire \cu_ru/add0_2/c57 ;
  wire \cu_ru/add0_2/c59 ;
  wire \cu_ru/add0_2/c7 ;
  wire \cu_ru/add0_2/c9 ;
  wire \cu_ru/add0_2_co ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_000 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_001 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_002 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_003 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_004 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_005 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_006 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_007 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_008 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_009 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_010 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_011 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_012 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_013 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_014 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_015 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_016 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_017 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_018 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_019 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_020 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_021 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_022 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_023 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_024 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_025 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_026 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_027 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_028 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_029 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_030 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_031 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_032 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_033 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_034 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_035 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_036 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_037 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_038 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_039 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_040 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_041 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_042 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_043 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_044 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_045 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_046 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_047 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_048 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_049 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_050 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_051 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_052 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_053 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_054 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_055 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_056 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_057 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_058 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_059 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_060 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_061 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_062 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_063 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_000 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_001 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_002 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_003 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_004 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_005 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_006 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_007 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_008 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_009 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_010 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_011 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_012 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_013 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_014 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_015 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_016 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_017 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_018 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_019 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_020 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_021 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_022 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_023 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_024 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_025 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_026 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_027 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_028 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_029 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_030 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_031 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_032 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_033 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_034 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_035 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_036 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_037 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_038 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_039 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_040 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_041 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_042 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_043 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_044 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_045 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_046 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_047 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_048 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_049 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_050 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_051 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_052 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_053 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_054 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_055 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_056 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_057 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_058 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_059 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_060 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_061 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_062 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_063 ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c0_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c0_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c0_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c10_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c10_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c10_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c11_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c11_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c11_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c12_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c12_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c12_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c13_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c13_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c13_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c14_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c14_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c14_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c15_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c15_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c15_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c1_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c1_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c1_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c2_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c2_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c2_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c3_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c3_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c3_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c4_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c4_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c4_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c5_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c5_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c5_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c6_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c6_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c6_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c7_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c7_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c7_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c8_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c8_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c8_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c9_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c9_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r0_c9_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c0_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c0_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c0_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c10_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c10_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c10_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c11_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c11_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c11_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c12_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c12_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c12_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c13_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c13_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c13_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c14_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c14_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c14_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c15_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c15_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c15_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c1_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c1_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c1_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c2_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c2_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c2_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c3_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c3_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c3_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c4_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c4_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c4_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c5_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c5_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c5_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c6_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c6_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c6_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c7_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c7_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c7_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c8_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c8_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c8_we ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c9_mode ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c9_wclk ;
  wire \cu_ru/al_ram_gpr_al_u0_r1_c9_we ;
  wire \cu_ru/al_ram_gpr_do_i0_000 ;
  wire \cu_ru/al_ram_gpr_do_i0_001 ;
  wire \cu_ru/al_ram_gpr_do_i0_002 ;
  wire \cu_ru/al_ram_gpr_do_i0_003 ;
  wire \cu_ru/al_ram_gpr_do_i0_004 ;
  wire \cu_ru/al_ram_gpr_do_i0_005 ;
  wire \cu_ru/al_ram_gpr_do_i0_006 ;
  wire \cu_ru/al_ram_gpr_do_i0_007 ;
  wire \cu_ru/al_ram_gpr_do_i0_008 ;
  wire \cu_ru/al_ram_gpr_do_i0_009 ;
  wire \cu_ru/al_ram_gpr_do_i0_010 ;
  wire \cu_ru/al_ram_gpr_do_i0_011 ;
  wire \cu_ru/al_ram_gpr_do_i0_012 ;
  wire \cu_ru/al_ram_gpr_do_i0_013 ;
  wire \cu_ru/al_ram_gpr_do_i0_014 ;
  wire \cu_ru/al_ram_gpr_do_i0_015 ;
  wire \cu_ru/al_ram_gpr_do_i0_016 ;
  wire \cu_ru/al_ram_gpr_do_i0_017 ;
  wire \cu_ru/al_ram_gpr_do_i0_018 ;
  wire \cu_ru/al_ram_gpr_do_i0_019 ;
  wire \cu_ru/al_ram_gpr_do_i0_020 ;
  wire \cu_ru/al_ram_gpr_do_i0_021 ;
  wire \cu_ru/al_ram_gpr_do_i0_022 ;
  wire \cu_ru/al_ram_gpr_do_i0_023 ;
  wire \cu_ru/al_ram_gpr_do_i0_024 ;
  wire \cu_ru/al_ram_gpr_do_i0_025 ;
  wire \cu_ru/al_ram_gpr_do_i0_026 ;
  wire \cu_ru/al_ram_gpr_do_i0_027 ;
  wire \cu_ru/al_ram_gpr_do_i0_028 ;
  wire \cu_ru/al_ram_gpr_do_i0_029 ;
  wire \cu_ru/al_ram_gpr_do_i0_030 ;
  wire \cu_ru/al_ram_gpr_do_i0_031 ;
  wire \cu_ru/al_ram_gpr_do_i0_032 ;
  wire \cu_ru/al_ram_gpr_do_i0_033 ;
  wire \cu_ru/al_ram_gpr_do_i0_034 ;
  wire \cu_ru/al_ram_gpr_do_i0_035 ;
  wire \cu_ru/al_ram_gpr_do_i0_036 ;
  wire \cu_ru/al_ram_gpr_do_i0_037 ;
  wire \cu_ru/al_ram_gpr_do_i0_038 ;
  wire \cu_ru/al_ram_gpr_do_i0_039 ;
  wire \cu_ru/al_ram_gpr_do_i0_040 ;
  wire \cu_ru/al_ram_gpr_do_i0_041 ;
  wire \cu_ru/al_ram_gpr_do_i0_042 ;
  wire \cu_ru/al_ram_gpr_do_i0_043 ;
  wire \cu_ru/al_ram_gpr_do_i0_044 ;
  wire \cu_ru/al_ram_gpr_do_i0_045 ;
  wire \cu_ru/al_ram_gpr_do_i0_046 ;
  wire \cu_ru/al_ram_gpr_do_i0_047 ;
  wire \cu_ru/al_ram_gpr_do_i0_048 ;
  wire \cu_ru/al_ram_gpr_do_i0_049 ;
  wire \cu_ru/al_ram_gpr_do_i0_050 ;
  wire \cu_ru/al_ram_gpr_do_i0_051 ;
  wire \cu_ru/al_ram_gpr_do_i0_052 ;
  wire \cu_ru/al_ram_gpr_do_i0_053 ;
  wire \cu_ru/al_ram_gpr_do_i0_054 ;
  wire \cu_ru/al_ram_gpr_do_i0_055 ;
  wire \cu_ru/al_ram_gpr_do_i0_056 ;
  wire \cu_ru/al_ram_gpr_do_i0_057 ;
  wire \cu_ru/al_ram_gpr_do_i0_058 ;
  wire \cu_ru/al_ram_gpr_do_i0_059 ;
  wire \cu_ru/al_ram_gpr_do_i0_060 ;
  wire \cu_ru/al_ram_gpr_do_i0_061 ;
  wire \cu_ru/al_ram_gpr_do_i0_062 ;
  wire \cu_ru/al_ram_gpr_do_i0_063 ;
  wire \cu_ru/al_ram_gpr_do_i1_000 ;
  wire \cu_ru/al_ram_gpr_do_i1_001 ;
  wire \cu_ru/al_ram_gpr_do_i1_002 ;
  wire \cu_ru/al_ram_gpr_do_i1_003 ;
  wire \cu_ru/al_ram_gpr_do_i1_004 ;
  wire \cu_ru/al_ram_gpr_do_i1_005 ;
  wire \cu_ru/al_ram_gpr_do_i1_006 ;
  wire \cu_ru/al_ram_gpr_do_i1_007 ;
  wire \cu_ru/al_ram_gpr_do_i1_008 ;
  wire \cu_ru/al_ram_gpr_do_i1_009 ;
  wire \cu_ru/al_ram_gpr_do_i1_010 ;
  wire \cu_ru/al_ram_gpr_do_i1_011 ;
  wire \cu_ru/al_ram_gpr_do_i1_012 ;
  wire \cu_ru/al_ram_gpr_do_i1_013 ;
  wire \cu_ru/al_ram_gpr_do_i1_014 ;
  wire \cu_ru/al_ram_gpr_do_i1_015 ;
  wire \cu_ru/al_ram_gpr_do_i1_016 ;
  wire \cu_ru/al_ram_gpr_do_i1_017 ;
  wire \cu_ru/al_ram_gpr_do_i1_018 ;
  wire \cu_ru/al_ram_gpr_do_i1_019 ;
  wire \cu_ru/al_ram_gpr_do_i1_020 ;
  wire \cu_ru/al_ram_gpr_do_i1_021 ;
  wire \cu_ru/al_ram_gpr_do_i1_022 ;
  wire \cu_ru/al_ram_gpr_do_i1_023 ;
  wire \cu_ru/al_ram_gpr_do_i1_024 ;
  wire \cu_ru/al_ram_gpr_do_i1_025 ;
  wire \cu_ru/al_ram_gpr_do_i1_026 ;
  wire \cu_ru/al_ram_gpr_do_i1_027 ;
  wire \cu_ru/al_ram_gpr_do_i1_028 ;
  wire \cu_ru/al_ram_gpr_do_i1_029 ;
  wire \cu_ru/al_ram_gpr_do_i1_030 ;
  wire \cu_ru/al_ram_gpr_do_i1_031 ;
  wire \cu_ru/al_ram_gpr_do_i1_032 ;
  wire \cu_ru/al_ram_gpr_do_i1_033 ;
  wire \cu_ru/al_ram_gpr_do_i1_034 ;
  wire \cu_ru/al_ram_gpr_do_i1_035 ;
  wire \cu_ru/al_ram_gpr_do_i1_036 ;
  wire \cu_ru/al_ram_gpr_do_i1_037 ;
  wire \cu_ru/al_ram_gpr_do_i1_038 ;
  wire \cu_ru/al_ram_gpr_do_i1_039 ;
  wire \cu_ru/al_ram_gpr_do_i1_040 ;
  wire \cu_ru/al_ram_gpr_do_i1_041 ;
  wire \cu_ru/al_ram_gpr_do_i1_042 ;
  wire \cu_ru/al_ram_gpr_do_i1_043 ;
  wire \cu_ru/al_ram_gpr_do_i1_044 ;
  wire \cu_ru/al_ram_gpr_do_i1_045 ;
  wire \cu_ru/al_ram_gpr_do_i1_046 ;
  wire \cu_ru/al_ram_gpr_do_i1_047 ;
  wire \cu_ru/al_ram_gpr_do_i1_048 ;
  wire \cu_ru/al_ram_gpr_do_i1_049 ;
  wire \cu_ru/al_ram_gpr_do_i1_050 ;
  wire \cu_ru/al_ram_gpr_do_i1_051 ;
  wire \cu_ru/al_ram_gpr_do_i1_052 ;
  wire \cu_ru/al_ram_gpr_do_i1_053 ;
  wire \cu_ru/al_ram_gpr_do_i1_054 ;
  wire \cu_ru/al_ram_gpr_do_i1_055 ;
  wire \cu_ru/al_ram_gpr_do_i1_056 ;
  wire \cu_ru/al_ram_gpr_do_i1_057 ;
  wire \cu_ru/al_ram_gpr_do_i1_058 ;
  wire \cu_ru/al_ram_gpr_do_i1_059 ;
  wire \cu_ru/al_ram_gpr_do_i1_060 ;
  wire \cu_ru/al_ram_gpr_do_i1_061 ;
  wire \cu_ru/al_ram_gpr_do_i1_062 ;
  wire \cu_ru/al_ram_gpr_do_i1_063 ;
  wire \cu_ru/al_ram_gpr_r0_c0_mode ;
  wire \cu_ru/al_ram_gpr_r0_c0_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c0_we ;
  wire \cu_ru/al_ram_gpr_r0_c10_mode ;
  wire \cu_ru/al_ram_gpr_r0_c10_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c10_we ;
  wire \cu_ru/al_ram_gpr_r0_c11_mode ;
  wire \cu_ru/al_ram_gpr_r0_c11_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c11_we ;
  wire \cu_ru/al_ram_gpr_r0_c12_mode ;
  wire \cu_ru/al_ram_gpr_r0_c12_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c12_we ;
  wire \cu_ru/al_ram_gpr_r0_c13_mode ;
  wire \cu_ru/al_ram_gpr_r0_c13_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c13_we ;
  wire \cu_ru/al_ram_gpr_r0_c14_mode ;
  wire \cu_ru/al_ram_gpr_r0_c14_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c14_we ;
  wire \cu_ru/al_ram_gpr_r0_c15_mode ;
  wire \cu_ru/al_ram_gpr_r0_c15_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c15_we ;
  wire \cu_ru/al_ram_gpr_r0_c1_mode ;
  wire \cu_ru/al_ram_gpr_r0_c1_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c1_we ;
  wire \cu_ru/al_ram_gpr_r0_c2_mode ;
  wire \cu_ru/al_ram_gpr_r0_c2_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c2_we ;
  wire \cu_ru/al_ram_gpr_r0_c3_mode ;
  wire \cu_ru/al_ram_gpr_r0_c3_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c3_we ;
  wire \cu_ru/al_ram_gpr_r0_c4_mode ;
  wire \cu_ru/al_ram_gpr_r0_c4_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c4_we ;
  wire \cu_ru/al_ram_gpr_r0_c5_mode ;
  wire \cu_ru/al_ram_gpr_r0_c5_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c5_we ;
  wire \cu_ru/al_ram_gpr_r0_c6_mode ;
  wire \cu_ru/al_ram_gpr_r0_c6_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c6_we ;
  wire \cu_ru/al_ram_gpr_r0_c7_mode ;
  wire \cu_ru/al_ram_gpr_r0_c7_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c7_we ;
  wire \cu_ru/al_ram_gpr_r0_c8_mode ;
  wire \cu_ru/al_ram_gpr_r0_c8_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c8_we ;
  wire \cu_ru/al_ram_gpr_r0_c9_mode ;
  wire \cu_ru/al_ram_gpr_r0_c9_wclk ;
  wire \cu_ru/al_ram_gpr_r0_c9_we ;
  wire \cu_ru/al_ram_gpr_r1_c0_mode ;
  wire \cu_ru/al_ram_gpr_r1_c0_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c0_we ;
  wire \cu_ru/al_ram_gpr_r1_c10_mode ;
  wire \cu_ru/al_ram_gpr_r1_c10_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c10_we ;
  wire \cu_ru/al_ram_gpr_r1_c11_mode ;
  wire \cu_ru/al_ram_gpr_r1_c11_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c11_we ;
  wire \cu_ru/al_ram_gpr_r1_c12_mode ;
  wire \cu_ru/al_ram_gpr_r1_c12_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c12_we ;
  wire \cu_ru/al_ram_gpr_r1_c13_mode ;
  wire \cu_ru/al_ram_gpr_r1_c13_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c13_we ;
  wire \cu_ru/al_ram_gpr_r1_c14_mode ;
  wire \cu_ru/al_ram_gpr_r1_c14_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c14_we ;
  wire \cu_ru/al_ram_gpr_r1_c15_mode ;
  wire \cu_ru/al_ram_gpr_r1_c15_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c15_we ;
  wire \cu_ru/al_ram_gpr_r1_c1_mode ;
  wire \cu_ru/al_ram_gpr_r1_c1_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c1_we ;
  wire \cu_ru/al_ram_gpr_r1_c2_mode ;
  wire \cu_ru/al_ram_gpr_r1_c2_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c2_we ;
  wire \cu_ru/al_ram_gpr_r1_c3_mode ;
  wire \cu_ru/al_ram_gpr_r1_c3_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c3_we ;
  wire \cu_ru/al_ram_gpr_r1_c4_mode ;
  wire \cu_ru/al_ram_gpr_r1_c4_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c4_we ;
  wire \cu_ru/al_ram_gpr_r1_c5_mode ;
  wire \cu_ru/al_ram_gpr_r1_c5_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c5_we ;
  wire \cu_ru/al_ram_gpr_r1_c6_mode ;
  wire \cu_ru/al_ram_gpr_r1_c6_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c6_we ;
  wire \cu_ru/al_ram_gpr_r1_c7_mode ;
  wire \cu_ru/al_ram_gpr_r1_c7_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c7_we ;
  wire \cu_ru/al_ram_gpr_r1_c8_mode ;
  wire \cu_ru/al_ram_gpr_r1_c8_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c8_we ;
  wire \cu_ru/al_ram_gpr_r1_c9_mode ;
  wire \cu_ru/al_ram_gpr_r1_c9_wclk ;
  wire \cu_ru/al_ram_gpr_r1_c9_we ;
  wire \cu_ru/csr_satp/n0 ;
  wire \cu_ru/m_cycle_event/add0/c11 ;
  wire \cu_ru/m_cycle_event/add0/c15 ;
  wire \cu_ru/m_cycle_event/add0/c19 ;
  wire \cu_ru/m_cycle_event/add0/c23 ;
  wire \cu_ru/m_cycle_event/add0/c27 ;
  wire \cu_ru/m_cycle_event/add0/c3 ;
  wire \cu_ru/m_cycle_event/add0/c31 ;
  wire \cu_ru/m_cycle_event/add0/c35 ;
  wire \cu_ru/m_cycle_event/add0/c39 ;
  wire \cu_ru/m_cycle_event/add0/c43 ;
  wire \cu_ru/m_cycle_event/add0/c47 ;
  wire \cu_ru/m_cycle_event/add0/c51 ;
  wire \cu_ru/m_cycle_event/add0/c55 ;
  wire \cu_ru/m_cycle_event/add0/c59 ;
  wire \cu_ru/m_cycle_event/add0/c63 ;
  wire \cu_ru/m_cycle_event/add0/c7 ;
  wire \cu_ru/m_cycle_event/add1/c11 ;
  wire \cu_ru/m_cycle_event/add1/c15 ;
  wire \cu_ru/m_cycle_event/add1/c19 ;
  wire \cu_ru/m_cycle_event/add1/c23 ;
  wire \cu_ru/m_cycle_event/add1/c27 ;
  wire \cu_ru/m_cycle_event/add1/c3 ;
  wire \cu_ru/m_cycle_event/add1/c31 ;
  wire \cu_ru/m_cycle_event/add1/c35 ;
  wire \cu_ru/m_cycle_event/add1/c39 ;
  wire \cu_ru/m_cycle_event/add1/c43 ;
  wire \cu_ru/m_cycle_event/add1/c47 ;
  wire \cu_ru/m_cycle_event/add1/c51 ;
  wire \cu_ru/m_cycle_event/add1/c55 ;
  wire \cu_ru/m_cycle_event/add1/c59 ;
  wire \cu_ru/m_cycle_event/add1/c63 ;
  wire \cu_ru/m_cycle_event/add1/c7 ;
  wire \cu_ru/m_cycle_event/mcountinhibit[2] ;  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(16)
  wire \cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ;
  wire \cu_ru/m_cycle_event/n13 ;
  wire \cu_ru/m_s_cause/mux2_b0_sel_is_2_o ;
  wire \cu_ru/m_s_cause/mux4_b0_sel_is_2_o ;
  wire \cu_ru/m_s_cause/mux7_b10_sel_is_0_o ;
  wire \cu_ru/m_s_epc/add0/c11 ;
  wire \cu_ru/m_s_epc/add0/c15 ;
  wire \cu_ru/m_s_epc/add0/c19 ;
  wire \cu_ru/m_s_epc/add0/c23 ;
  wire \cu_ru/m_s_epc/add0/c27 ;
  wire \cu_ru/m_s_epc/add0/c3 ;
  wire \cu_ru/m_s_epc/add0/c31 ;
  wire \cu_ru/m_s_epc/add0/c35 ;
  wire \cu_ru/m_s_epc/add0/c39 ;
  wire \cu_ru/m_s_epc/add0/c43 ;
  wire \cu_ru/m_s_epc/add0/c47 ;
  wire \cu_ru/m_s_epc/add0/c51 ;
  wire \cu_ru/m_s_epc/add0/c55 ;
  wire \cu_ru/m_s_epc/add0/c59 ;
  wire \cu_ru/m_s_epc/add0/c7 ;
  wire \cu_ru/m_s_epc/mux4_b0_sel_is_2_o ;
  wire \cu_ru/m_s_epc/mux6_b0_sel_is_2_o ;
  wire \cu_ru/m_s_ie/n0 ;
  wire \cu_ru/m_s_ie/u11_sel_is_0_o ;
  wire \cu_ru/m_s_ip/n0 ;
  wire \cu_ru/m_s_ip/seip ;  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(28)
  wire \cu_ru/m_s_ip/u11_sel_is_0_o ;
  wire \cu_ru/m_s_ip/u12_sel_is_2_o ;
  wire \cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ;
  wire \cu_ru/m_s_scratch/n0 ;
  wire \cu_ru/m_s_status/mux3_b0_sel_is_2_o ;
  wire \cu_ru/m_s_status/n0 ;
  wire \cu_ru/m_s_status/n2 ;
  wire \cu_ru/m_s_status/u14_sel_is_2_o ;
  wire \cu_ru/m_s_status/u34_sel_is_0_o ;
  wire \cu_ru/m_s_tval/mux3_b0_sel_is_2_o ;
  wire \cu_ru/m_s_tval/mux5_b0_sel_is_2_o ;
  wire \cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ;
  wire \cu_ru/m_s_tvec/n0 ;
  wire \cu_ru/mcountinhibit ;  // ../../RTL/CPU/CU&RU/cu_ru.v(639)
  wire \cu_ru/medeleg_exc_ctrl/ecu_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(78)
  wire \cu_ru/medeleg_exc_ctrl/ecu_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(92)
  wire \cu_ru/medeleg_exc_ctrl/iaf_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(71)
  wire \cu_ru/medeleg_exc_ctrl/iam_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(70)
  wire \cu_ru/medeleg_exc_ctrl/iam_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(84)
  wire \cu_ru/medeleg_exc_ctrl/ii_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(86)
  wire \cu_ru/medeleg_exc_ctrl/laf_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(75)
  wire \cu_ru/medeleg_exc_ctrl/laf_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(89)
  wire \cu_ru/medeleg_exc_ctrl/lam_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(74)
  wire \cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/n0 ;
  wire \cu_ru/medeleg_exc_ctrl/n80_neg_lutinv ;
  wire \cu_ru/medeleg_exc_ctrl/n84_neg_lutinv ;
  wire \cu_ru/medeleg_exc_ctrl/n85_neg_lutinv ;
  wire \cu_ru/medeleg_exc_ctrl/n87_neg_lutinv ;
  wire \cu_ru/medeleg_exc_ctrl/saf_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(77)
  wire \cu_ru/medeleg_exc_ctrl/sam_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(90)
  wire \cu_ru/medeleg_exc_ctrl/spf_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(82)
  wire \cu_ru/medeleg_exc_ctrl/spf_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(96)
  wire \cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o ;
  wire \cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ;
  wire \cu_ru/mideleg_int_ctrl/n0 ;
  wire \cu_ru/mideleg_int_ctrl/n28_lutinv ;
  wire \cu_ru/mideleg_int_ctrl/n29_lutinv ;
  wire \cu_ru/mideleg_int_ctrl/n33_neg_lutinv ;
  wire \cu_ru/mideleg_int_ctrl/sei_ack_m ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(61)
  wire \cu_ru/mideleg_int_ctrl/sti_ack_s ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(67)
  wire \cu_ru/mie ;  // ../../RTL/CPU/CU&RU/cu_ru.v(381)
  wire \cu_ru/mux34_b0_sel_is_2_o ;
  wire \cu_ru/n41 ;
  wire \cu_ru/n45_lutinv ;
  wire \cu_ru/n53_0_al_n1985 ;
  wire \cu_ru/n53_1_al_n1986 ;
  wire \cu_ru/n53_lutinv ;
  wire \cu_ru/n66_lutinv ;
  wire \cu_ru/read_cycle_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(220)
  wire \cu_ru/read_instret_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(222)
  wire \cu_ru/read_mcause_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(248)
  wire \cu_ru/read_mcycle_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(254)
  wire \cu_ru/read_medeleg_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(241)
  wire \cu_ru/read_mepc_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(247)
  wire \cu_ru/read_mideleg_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(242)
  wire \cu_ru/read_minstret_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(255)
  wire \cu_ru/read_mip_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(250)
  wire \cu_ru/read_mscratch_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(246)
  wire \cu_ru/read_mtval_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(249)
  wire \cu_ru/read_mtvec_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(244)
  wire \cu_ru/read_satp_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(234)
  wire \cu_ru/read_scause_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(231)
  wire \cu_ru/read_sepc_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(230)
  wire \cu_ru/read_sscratch_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(229)
  wire \cu_ru/read_stval_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(232)
  wire \cu_ru/read_stvec_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(227)
  wire \cu_ru/read_time_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(221)
  wire \cu_ru/sub0/c1 ;
  wire \cu_ru/sub0/c3 ;
  wire \cu_ru/sub1/c1 ;
  wire \cu_ru/sub1/c3 ;
  wire \cu_ru/sub2/c1 ;
  wire \cu_ru/sub2/c3 ;
  wire \cu_ru/trap_target_m ;  // ../../RTL/CPU/CU&RU/cu_ru.v(148)
  wire ex_csr_write;  // ../../RTL/CPU/prv464_top.v(145)
  wire ex_ebreak;  // ../../RTL/CPU/prv464_top.v(171)
  wire ex_ecall;  // ../../RTL/CPU/prv464_top.v(170)
  wire ex_gpr_write;  // ../../RTL/CPU/prv464_top.v(146)
  wire ex_ill_ins;  // ../../RTL/CPU/prv464_top.v(167)
  wire ex_ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(162)
  wire ex_ins_addr_mis;  // ../../RTL/CPU/prv464_top.v(163)
  wire ex_ins_page_fault;  // ../../RTL/CPU/prv464_top.v(164)
  wire ex_int_acc;  // ../../RTL/CPU/prv464_top.v(165)
  wire ex_jmp;  // ../../RTL/CPU/prv464_top.v(161)
  wire ex_more_exception_neg_lutinv;
  wire ex_nop;  // ../../RTL/CPU/prv464_top.v(580)
  wire ex_system;  // ../../RTL/CPU/prv464_top.v(160)
  wire ex_valid;  // ../../RTL/CPU/prv464_top.v(166)
  wire \exu/alu_au/add0/c11 ;
  wire \exu/alu_au/add0/c15 ;
  wire \exu/alu_au/add0/c19 ;
  wire \exu/alu_au/add0/c23 ;
  wire \exu/alu_au/add0/c27 ;
  wire \exu/alu_au/add0/c3 ;
  wire \exu/alu_au/add0/c31 ;
  wire \exu/alu_au/add0/c35 ;
  wire \exu/alu_au/add0/c39 ;
  wire \exu/alu_au/add0/c43 ;
  wire \exu/alu_au/add0/c47 ;
  wire \exu/alu_au/add0/c51 ;
  wire \exu/alu_au/add0/c55 ;
  wire \exu/alu_au/add0/c59 ;
  wire \exu/alu_au/add0/c63 ;
  wire \exu/alu_au/add0/c7 ;
  wire \exu/alu_au/add1/c1 ;
  wire \exu/alu_au/add1/c11 ;
  wire \exu/alu_au/add1/c13 ;
  wire \exu/alu_au/add1/c15 ;
  wire \exu/alu_au/add1/c17 ;
  wire \exu/alu_au/add1/c19 ;
  wire \exu/alu_au/add1/c21 ;
  wire \exu/alu_au/add1/c23 ;
  wire \exu/alu_au/add1/c25 ;
  wire \exu/alu_au/add1/c27 ;
  wire \exu/alu_au/add1/c29 ;
  wire \exu/alu_au/add1/c3 ;
  wire \exu/alu_au/add1/c31 ;
  wire \exu/alu_au/add1/c5 ;
  wire \exu/alu_au/add1/c7 ;
  wire \exu/alu_au/add1/c9 ;
  wire \exu/alu_au/add2/c11 ;
  wire \exu/alu_au/add2/c15 ;
  wire \exu/alu_au/add2/c19 ;
  wire \exu/alu_au/add2/c23 ;
  wire \exu/alu_au/add2/c27 ;
  wire \exu/alu_au/add2/c3 ;
  wire \exu/alu_au/add2/c31 ;
  wire \exu/alu_au/add2/c35 ;
  wire \exu/alu_au/add2/c39 ;
  wire \exu/alu_au/add2/c43 ;
  wire \exu/alu_au/add2/c47 ;
  wire \exu/alu_au/add2/c51 ;
  wire \exu/alu_au/add2/c55 ;
  wire \exu/alu_au/add2/c59 ;
  wire \exu/alu_au/add2/c63 ;
  wire \exu/alu_au/add2/c7 ;
  wire \exu/alu_au/ds1_light_than_ds2_lutinv ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(67)
  wire \exu/alu_au/lt0_c1 ;
  wire \exu/alu_au/lt0_c11 ;
  wire \exu/alu_au/lt0_c13 ;
  wire \exu/alu_au/lt0_c15 ;
  wire \exu/alu_au/lt0_c17 ;
  wire \exu/alu_au/lt0_c19 ;
  wire \exu/alu_au/lt0_c21 ;
  wire \exu/alu_au/lt0_c23 ;
  wire \exu/alu_au/lt0_c25 ;
  wire \exu/alu_au/lt0_c27 ;
  wire \exu/alu_au/lt0_c29 ;
  wire \exu/alu_au/lt0_c3 ;
  wire \exu/alu_au/lt0_c31 ;
  wire \exu/alu_au/lt0_c33 ;
  wire \exu/alu_au/lt0_c35 ;
  wire \exu/alu_au/lt0_c37 ;
  wire \exu/alu_au/lt0_c39 ;
  wire \exu/alu_au/lt0_c41 ;
  wire \exu/alu_au/lt0_c43 ;
  wire \exu/alu_au/lt0_c45 ;
  wire \exu/alu_au/lt0_c47 ;
  wire \exu/alu_au/lt0_c49 ;
  wire \exu/alu_au/lt0_c5 ;
  wire \exu/alu_au/lt0_c51 ;
  wire \exu/alu_au/lt0_c53 ;
  wire \exu/alu_au/lt0_c55 ;
  wire \exu/alu_au/lt0_c57 ;
  wire \exu/alu_au/lt0_c59 ;
  wire \exu/alu_au/lt0_c61 ;
  wire \exu/alu_au/lt0_c63 ;
  wire \exu/alu_au/lt0_c7 ;
  wire \exu/alu_au/lt0_c9 ;
  wire \exu/alu_au/lt1_c1 ;
  wire \exu/alu_au/lt1_c11 ;
  wire \exu/alu_au/lt1_c13 ;
  wire \exu/alu_au/lt1_c15 ;
  wire \exu/alu_au/lt1_c17 ;
  wire \exu/alu_au/lt1_c19 ;
  wire \exu/alu_au/lt1_c21 ;
  wire \exu/alu_au/lt1_c23 ;
  wire \exu/alu_au/lt1_c25 ;
  wire \exu/alu_au/lt1_c27 ;
  wire \exu/alu_au/lt1_c29 ;
  wire \exu/alu_au/lt1_c3 ;
  wire \exu/alu_au/lt1_c31 ;
  wire \exu/alu_au/lt1_c33 ;
  wire \exu/alu_au/lt1_c35 ;
  wire \exu/alu_au/lt1_c37 ;
  wire \exu/alu_au/lt1_c39 ;
  wire \exu/alu_au/lt1_c41 ;
  wire \exu/alu_au/lt1_c43 ;
  wire \exu/alu_au/lt1_c45 ;
  wire \exu/alu_au/lt1_c47 ;
  wire \exu/alu_au/lt1_c49 ;
  wire \exu/alu_au/lt1_c5 ;
  wire \exu/alu_au/lt1_c51 ;
  wire \exu/alu_au/lt1_c53 ;
  wire \exu/alu_au/lt1_c55 ;
  wire \exu/alu_au/lt1_c57 ;
  wire \exu/alu_au/lt1_c59 ;
  wire \exu/alu_au/lt1_c61 ;
  wire \exu/alu_au/lt1_c63 ;
  wire \exu/alu_au/lt1_c7 ;
  wire \exu/alu_au/lt1_c9 ;
  wire \exu/alu_au/n12 ;
  wire \exu/alu_au/n15 ;
  wire \exu/alu_au/n5 ;
  wire \exu/c_fence_lutinv ;  // ../../RTL/CPU/EX/exu.v(182)
  wire \exu/c_load_1_lutinv ;  // ../../RTL/CPU/EX/exu.v(176)
  wire \exu/c_stb_lutinv ;  // ../../RTL/CPU/EX/exu.v(173)
  wire \exu/load_addr_mis ;  // ../../RTL/CPU/EX/exu.v(202)
  wire \exu/lsu/mux27_b56_sel_is_3_o ;
  wire \exu/lsu/n0_lutinv ;
  wire \exu/lsu/n2_lutinv ;
  wire \exu/lsu/n51 ;
  wire \exu/lsu/n53 ;
  wire \exu/lsu/n56 ;
  wire \exu/lsu/n5_lutinv ;
  wire \exu/lsu/n8_lutinv ;
  wire \exu/mux27_b32_sel_is_1_o ;
  wire \exu/n10 ;
  wire \exu/n138_lutinv ;
  wire \exu/n17_lutinv ;
  wire \exu/n19 ;
  wire \exu/n49 ;
  wire \exu/n59_lutinv ;
  wire \exu/n60_lutinv ;
  wire \exu/n86 ;
  wire \exu/shift_multi_ready ;  // ../../RTL/CPU/EX/exu.v(209)
  wire \exu/store_addr_mis ;  // ../../RTL/CPU/EX/exu.v(203)
  wire \exu/sub0/c1 ;
  wire \exu/sub0/c3 ;
  wire \exu/sub0/c5 ;
  wire \exu/sub0/c7 ;
  wire hready_pad;  // ../../RTL/CPU/prv464_top.v(31)
  wire hresp_pad;  // ../../RTL/CPU/prv464_top.v(32)
  wire hwrite_pad;  // ../../RTL/CPU/prv464_top.v(23)
  wire id_hold;  // ../../RTL/CPU/prv464_top.v(177)
  wire id_ill_ins;  // ../../RTL/CPU/prv464_top.v(176)
  wire id_ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(92)
  wire id_ins_addr_mis;  // ../../RTL/CPU/prv464_top.v(93)
  wire id_ins_page_fault;  // ../../RTL/CPU/prv464_top.v(94)
  wire id_int_acc;  // ../../RTL/CPU/prv464_top.v(95)
  wire id_nop_neg_lutinv;
  wire id_system;  // ../../RTL/CPU/prv464_top.v(175)
  wire id_valid;  // ../../RTL/CPU/prv464_top.v(96)
  wire if_hold;  // ../../RTL/CPU/prv464_top.v(263)
  wire \ins_dec/dec_ins_dec_fault_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(336)
  wire \ins_dec/funct3_0_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(172)
  wire \ins_dec/funct5_8_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(189)
  wire \ins_dec/funct6_0_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(214)
  wire \ins_dec/funct7_0_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(220)
  wire \ins_dec/funct7_32_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(217)
  wire \ins_dec/funct7_8_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(219)
  wire \ins_dec/ins_addw ;  // ../../RTL/CPU/ID/ins_dec.v(299)
  wire \ins_dec/ins_fence ;  // ../../RTL/CPU/ID/ins_dec.v(282)
  wire \ins_dec/ins_sfencevma ;  // ../../RTL/CPU/ID/ins_dec.v(331)
  wire \ins_dec/ins_slli ;  // ../../RTL/CPU/ID/ins_dec.v(269)
  wire \ins_dec/ins_srai ;  // ../../RTL/CPU/ID/ins_dec.v(271)
  wire \ins_dec/ins_srli ;  // ../../RTL/CPU/ID/ins_dec.v(270)
  wire \ins_dec/mux13_b0_sel_is_0_o ;
  wire \ins_dec/mux19_b10_sel_is_2_o ;
  wire \ins_dec/mux24_b10_sel_is_0_o ;
  wire \ins_dec/mux27_b12_sel_is_0_o ;
  wire \ins_dec/mux27_b56_sel_is_0_o ;
  wire \ins_dec/n107 ;
  wire \ins_dec/n141_lutinv ;
  wire \ins_dec/n149_lutinv ;
  wire \ins_dec/n198_lutinv ;
  wire \ins_dec/n232 ;
  wire \ins_dec/n235 ;
  wire \ins_dec/n239 ;
  wire \ins_dec/n302 ;
  wire \ins_dec/n35_lutinv ;
  wire \ins_dec/n38 ;
  wire \ins_dec/n48_lutinv ;
  wire \ins_dec/n57_neg_lutinv ;
  wire \ins_dec/n59 ;
  wire \ins_dec/n71 ;
  wire \ins_dec/n80_lutinv ;
  wire \ins_dec/op_32_imm_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(158)
  wire \ins_dec/op_32_reg_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(167)
  wire \ins_dec/op_amo ;  // ../../RTL/CPU/ID/ins_dec.v(168)
  wire \ins_dec/op_load ;  // ../../RTL/CPU/ID/ins_dec.v(165)
  wire \ins_dec/op_lui_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(159)
  wire \ins_dec/op_store ;  // ../../RTL/CPU/ID/ins_dec.v(164)
  wire \ins_dec/qbyte ;  // ../../RTL/CPU/ID/ins_dec.v(236)
  wire \ins_dec/u461_sel_is_0_o ;
  wire \ins_dec/u478_sel_is_0_o ;
  wire \ins_fetch/add0/c1 ;
  wire \ins_fetch/add0/c11 ;
  wire \ins_fetch/add0/c13 ;
  wire \ins_fetch/add0/c15 ;
  wire \ins_fetch/add0/c17 ;
  wire \ins_fetch/add0/c19 ;
  wire \ins_fetch/add0/c21 ;
  wire \ins_fetch/add0/c23 ;
  wire \ins_fetch/add0/c25 ;
  wire \ins_fetch/add0/c27 ;
  wire \ins_fetch/add0/c29 ;
  wire \ins_fetch/add0/c3 ;
  wire \ins_fetch/add0/c31 ;
  wire \ins_fetch/add0/c33 ;
  wire \ins_fetch/add0/c35 ;
  wire \ins_fetch/add0/c37 ;
  wire \ins_fetch/add0/c39 ;
  wire \ins_fetch/add0/c41 ;
  wire \ins_fetch/add0/c43 ;
  wire \ins_fetch/add0/c45 ;
  wire \ins_fetch/add0/c47 ;
  wire \ins_fetch/add0/c49 ;
  wire \ins_fetch/add0/c5 ;
  wire \ins_fetch/add0/c51 ;
  wire \ins_fetch/add0/c53 ;
  wire \ins_fetch/add0/c55 ;
  wire \ins_fetch/add0/c57 ;
  wire \ins_fetch/add0/c59 ;
  wire \ins_fetch/add0/c61 ;
  wire \ins_fetch/add0/c7 ;
  wire \ins_fetch/add0/c9 ;
  wire \ins_fetch/n25 ;
  wire \ins_fetch/n27 ;
  wire \ins_fetch/n9 ;
  wire int_req;  // ../../RTL/CPU/prv464_top.v(259)
  wire jmp;  // ../../RTL/CPU/prv464_top.v(127)
  wire load;  // ../../RTL/CPU/prv464_top.v(136)
  wire load_acc_fault;  // ../../RTL/CPU/prv464_top.v(83)
  wire mem_csr_data_add;  // ../../RTL/CPU/prv464_top.v(116)
  wire mem_csr_data_and;  // ../../RTL/CPU/prv464_top.v(117)
  wire mem_csr_data_ds2;  // ../../RTL/CPU/prv464_top.v(115)
  wire mem_csr_data_max;  // ../../RTL/CPU/prv464_top.v(120)
  wire mem_csr_data_min;  // ../../RTL/CPU/prv464_top.v(121)
  wire mem_csr_data_or;  // ../../RTL/CPU/prv464_top.v(118)
  wire mem_csr_data_xor;  // ../../RTL/CPU/prv464_top.v(119)
  wire mprv;  // ../../RTL/CPU/prv464_top.v(53)
  wire mxr;  // ../../RTL/CPU/prv464_top.v(52)
  wire pc_jmp;  // ../../RTL/CPU/prv464_top.v(522)
  wire \pip_ctrl/eq2/xor_i0[1]_i1[1]_o_lutinv ;
  wire \pip_ctrl/ex_exception ;  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(80)
  wire \pip_ctrl/id_ex_war_lutinv ;  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(83)
  wire \pip_ctrl/id_exception ;  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(79)
  wire \pip_ctrl/n34 ;
  wire \pip_ctrl/n36_lutinv ;
  wire pip_flush;  // ../../RTL/CPU/prv464_top.v(265)
  wire rd_data_add;  // ../../RTL/CPU/prv464_top.v(104)
  wire rd_data_and;  // ../../RTL/CPU/prv464_top.v(106)
  wire rd_data_ds1;  // ../../RTL/CPU/prv464_top.v(103)
  wire rd_data_or;  // ../../RTL/CPU/prv464_top.v(107)
  wire rd_data_slt;  // ../../RTL/CPU/prv464_top.v(109)
  wire rd_data_sub;  // ../../RTL/CPU/prv464_top.v(105)
  wire rd_data_xor;  // ../../RTL/CPU/prv464_top.v(108)
  wire read;  // ../../RTL/CPU/prv464_top.v(81)
  wire rst_pad;  // ../../RTL/CPU/prv464_top.v(20)
  wire s_ext_int_pad;  // ../../RTL/CPU/prv464_top.v(40)
  wire shift_l;  // ../../RTL/CPU/prv464_top.v(142)
  wire shift_r;  // ../../RTL/CPU/prv464_top.v(141)
  wire store;  // ../../RTL/CPU/prv464_top.v(137)
  wire sum;  // ../../RTL/CPU/prv464_top.v(51)
  wire tsr;  // ../../RTL/CPU/prv464_top.v(50)
  wire tvm;  // ../../RTL/CPU/prv464_top.v(49)
  wire tw;  // ../../RTL/CPU/prv464_top.v(309)
  wire unsign;  // ../../RTL/CPU/prv464_top.v(128)
  wire wb_csr_write;  // ../../RTL/CPU/prv464_top.v(520)
  wire wb_ebreak;  // ../../RTL/CPU/prv464_top.v(547)
  wire wb_ecall;  // ../../RTL/CPU/prv464_top.v(546)
  wire wb_gpr_write;  // ../../RTL/CPU/prv464_top.v(521)
  wire wb_ill_ins;  // ../../RTL/CPU/prv464_top.v(543)
  wire wb_ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(532)
  wire wb_ins_addr_mis;  // ../../RTL/CPU/prv464_top.v(533)
  wire wb_ins_page_fault;  // ../../RTL/CPU/prv464_top.v(534)
  wire wb_int_acc;  // ../../RTL/CPU/prv464_top.v(541)
  wire wb_jmp;  // ../../RTL/CPU/prv464_top.v(531)
  wire wb_ld_acc_fault;  // ../../RTL/CPU/prv464_top.v(537)
  wire wb_ld_addr_mis;  // ../../RTL/CPU/prv464_top.v(535)
  wire wb_ld_page_fault;  // ../../RTL/CPU/prv464_top.v(539)
  wire wb_st_acc_fault;  // ../../RTL/CPU/prv464_top.v(538)
  wire wb_st_addr_mis;  // ../../RTL/CPU/prv464_top.v(536)
  wire wb_st_page_fault;  // ../../RTL/CPU/prv464_top.v(540)
  wire wb_system;  // ../../RTL/CPU/prv464_top.v(530)
  wire wb_valid;  // ../../RTL/CPU/prv464_top.v(542)
  wire write;  // ../../RTL/CPU/prv464_top.v(82)

  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1926 (
    .ipad(cacheability_block[31]),
    .di(cacheability_block_pad[31]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1927 (
    .ipad(cacheability_block[30]),
    .di(cacheability_block_pad[30]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1928 (
    .ipad(cacheability_block[29]),
    .di(cacheability_block_pad[29]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1929 (
    .ipad(cacheability_block[28]),
    .di(cacheability_block_pad[28]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1930 (
    .ipad(cacheability_block[27]),
    .di(cacheability_block_pad[27]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1931 (
    .ipad(cacheability_block[26]),
    .di(cacheability_block_pad[26]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1932 (
    .ipad(cacheability_block[25]),
    .di(cacheability_block_pad[25]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1933 (
    .ipad(cacheability_block[24]),
    .di(cacheability_block_pad[24]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1934 (
    .ipad(cacheability_block[23]),
    .di(cacheability_block_pad[23]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1935 (
    .ipad(cacheability_block[22]),
    .di(cacheability_block_pad[22]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1936 (
    .ipad(cacheability_block[21]),
    .di(cacheability_block_pad[21]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1937 (
    .ipad(cacheability_block[20]),
    .di(cacheability_block_pad[20]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1938 (
    .ipad(cacheability_block[19]),
    .di(cacheability_block_pad[19]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1939 (
    .ipad(cacheability_block[18]),
    .di(cacheability_block_pad[18]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1940 (
    .ipad(cacheability_block[17]),
    .di(cacheability_block_pad[17]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1941 (
    .ipad(cacheability_block[16]),
    .di(cacheability_block_pad[16]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1942 (
    .ipad(cacheability_block[15]),
    .di(cacheability_block_pad[15]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1943 (
    .ipad(cacheability_block[14]),
    .di(cacheability_block_pad[14]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1944 (
    .ipad(cacheability_block[13]),
    .di(cacheability_block_pad[13]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1945 (
    .ipad(cacheability_block[12]),
    .di(cacheability_block_pad[12]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1946 (
    .ipad(cacheability_block[11]),
    .di(cacheability_block_pad[11]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1947 (
    .ipad(cacheability_block[10]),
    .di(cacheability_block_pad[10]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1948 (
    .ipad(cacheability_block[9]),
    .di(cacheability_block_pad[9]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1949 (
    .ipad(cacheability_block[8]),
    .di(cacheability_block_pad[8]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1950 (
    .ipad(cacheability_block[7]),
    .di(cacheability_block_pad[7]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1951 (
    .ipad(cacheability_block[6]),
    .di(cacheability_block_pad[6]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1952 (
    .ipad(cacheability_block[5]),
    .di(cacheability_block_pad[5]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1953 (
    .ipad(cacheability_block[4]),
    .di(cacheability_block_pad[4]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1954 (
    .ipad(cacheability_block[3]),
    .di(cacheability_block_pad[3]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1955 (
    .ipad(cacheability_block[2]),
    .di(cacheability_block_pad[2]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1956 (
    .ipad(cacheability_block[1]),
    .di(cacheability_block_pad[1]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1957 (
    .ipad(cacheability_block[0]),
    .di(cacheability_block_pad[0]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1958 (
    .ipad(clk),
    .di(clk_pad));  // ../../RTL/CPU/prv464_top.v(19)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1959 (
    .do({open_n562,open_n563,open_n564,haddr_pad[63]}),
    .opad(haddr[63]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1960 (
    .do({open_n579,open_n580,open_n581,haddr_pad[62]}),
    .opad(haddr[62]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1961 (
    .do({open_n596,open_n597,open_n598,haddr_pad[61]}),
    .opad(haddr[61]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1962 (
    .do({open_n613,open_n614,open_n615,haddr_pad[60]}),
    .opad(haddr[60]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1963 (
    .do({open_n630,open_n631,open_n632,haddr_pad[59]}),
    .opad(haddr[59]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1964 (
    .do({open_n647,open_n648,open_n649,haddr_pad[58]}),
    .opad(haddr[58]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1965 (
    .do({open_n664,open_n665,open_n666,haddr_pad[57]}),
    .opad(haddr[57]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1966 (
    .do({open_n681,open_n682,open_n683,haddr_pad[56]}),
    .opad(haddr[56]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1967 (
    .do({open_n698,open_n699,open_n700,haddr_pad[55]}),
    .opad(haddr[55]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1968 (
    .do({open_n715,open_n716,open_n717,haddr_pad[54]}),
    .opad(haddr[54]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1969 (
    .do({open_n732,open_n733,open_n734,haddr_pad[53]}),
    .opad(haddr[53]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1970 (
    .do({open_n749,open_n750,open_n751,haddr_pad[52]}),
    .opad(haddr[52]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1971 (
    .do({open_n766,open_n767,open_n768,haddr_pad[51]}),
    .opad(haddr[51]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1972 (
    .do({open_n783,open_n784,open_n785,haddr_pad[50]}),
    .opad(haddr[50]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1973 (
    .do({open_n800,open_n801,open_n802,haddr_pad[49]}),
    .opad(haddr[49]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1974 (
    .do({open_n817,open_n818,open_n819,haddr_pad[48]}),
    .opad(haddr[48]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1975 (
    .do({open_n834,open_n835,open_n836,haddr_pad[47]}),
    .opad(haddr[47]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1976 (
    .do({open_n851,open_n852,open_n853,haddr_pad[46]}),
    .opad(haddr[46]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1977 (
    .do({open_n868,open_n869,open_n870,haddr_pad[45]}),
    .opad(haddr[45]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1978 (
    .do({open_n885,open_n886,open_n887,haddr_pad[44]}),
    .opad(haddr[44]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1979 (
    .do({open_n902,open_n903,open_n904,haddr_pad[43]}),
    .opad(haddr[43]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1980 (
    .do({open_n919,open_n920,open_n921,haddr_pad[42]}),
    .opad(haddr[42]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1981 (
    .do({open_n936,open_n937,open_n938,haddr_pad[41]}),
    .opad(haddr[41]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1982 (
    .do({open_n953,open_n954,open_n955,haddr_pad[40]}),
    .opad(haddr[40]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1983 (
    .do({open_n970,open_n971,open_n972,haddr_pad[39]}),
    .opad(haddr[39]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1984 (
    .do({open_n987,open_n988,open_n989,haddr_pad[38]}),
    .opad(haddr[38]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1985 (
    .do({open_n1004,open_n1005,open_n1006,haddr_pad[37]}),
    .opad(haddr[37]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1986 (
    .do({open_n1021,open_n1022,open_n1023,haddr_pad[36]}),
    .opad(haddr[36]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1987 (
    .do({open_n1038,open_n1039,open_n1040,haddr_pad[35]}),
    .opad(haddr[35]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1988 (
    .do({open_n1055,open_n1056,open_n1057,haddr_pad[34]}),
    .opad(haddr[34]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1989 (
    .do({open_n1072,open_n1073,open_n1074,haddr_pad[33]}),
    .opad(haddr[33]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1990 (
    .do({open_n1089,open_n1090,open_n1091,haddr_pad[32]}),
    .opad(haddr[32]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1991 (
    .do({open_n1106,open_n1107,open_n1108,haddr_pad[31]}),
    .opad(haddr[31]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1992 (
    .do({open_n1123,open_n1124,open_n1125,haddr_pad[30]}),
    .opad(haddr[30]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1993 (
    .do({open_n1140,open_n1141,open_n1142,haddr_pad[29]}),
    .opad(haddr[29]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1994 (
    .do({open_n1157,open_n1158,open_n1159,haddr_pad[28]}),
    .opad(haddr[28]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1995 (
    .do({open_n1174,open_n1175,open_n1176,haddr_pad[27]}),
    .opad(haddr[27]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1996 (
    .do({open_n1191,open_n1192,open_n1193,haddr_pad[26]}),
    .opad(haddr[26]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1997 (
    .do({open_n1208,open_n1209,open_n1210,haddr_pad[25]}),
    .opad(haddr[25]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1998 (
    .do({open_n1225,open_n1226,open_n1227,haddr_pad[24]}),
    .opad(haddr[24]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1999 (
    .do({open_n1242,open_n1243,open_n1244,haddr_pad[23]}),
    .opad(haddr[23]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2000 (
    .do({open_n1259,open_n1260,open_n1261,haddr_pad[22]}),
    .opad(haddr[22]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2001 (
    .do({open_n1276,open_n1277,open_n1278,haddr_pad[21]}),
    .opad(haddr[21]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2002 (
    .do({open_n1293,open_n1294,open_n1295,haddr_pad[20]}),
    .opad(haddr[20]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2003 (
    .do({open_n1310,open_n1311,open_n1312,haddr_pad[19]}),
    .opad(haddr[19]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2004 (
    .do({open_n1327,open_n1328,open_n1329,haddr_pad[18]}),
    .opad(haddr[18]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2005 (
    .do({open_n1344,open_n1345,open_n1346,haddr_pad[17]}),
    .opad(haddr[17]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2006 (
    .do({open_n1361,open_n1362,open_n1363,haddr_pad[16]}),
    .opad(haddr[16]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2007 (
    .do({open_n1378,open_n1379,open_n1380,haddr_pad[15]}),
    .opad(haddr[15]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2008 (
    .do({open_n1395,open_n1396,open_n1397,haddr_pad[14]}),
    .opad(haddr[14]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2009 (
    .do({open_n1412,open_n1413,open_n1414,haddr_pad[13]}),
    .opad(haddr[13]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2010 (
    .do({open_n1429,open_n1430,open_n1431,haddr_pad[12]}),
    .opad(haddr[12]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2011 (
    .do({open_n1446,open_n1447,open_n1448,haddr_pad[11]}),
    .opad(haddr[11]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2012 (
    .do({open_n1463,open_n1464,open_n1465,haddr_pad[10]}),
    .opad(haddr[10]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2013 (
    .do({open_n1480,open_n1481,open_n1482,haddr_pad[9]}),
    .opad(haddr[9]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2014 (
    .do({open_n1497,open_n1498,open_n1499,haddr_pad[8]}),
    .opad(haddr[8]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2015 (
    .do({open_n1514,open_n1515,open_n1516,haddr_pad[7]}),
    .opad(haddr[7]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2016 (
    .do({open_n1531,open_n1532,open_n1533,haddr_pad[6]}),
    .opad(haddr[6]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2017 (
    .do({open_n1548,open_n1549,open_n1550,haddr_pad[5]}),
    .opad(haddr[5]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2018 (
    .do({open_n1565,open_n1566,open_n1567,haddr_pad[4]}),
    .opad(haddr[4]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2019 (
    .do({open_n1582,open_n1583,open_n1584,haddr_pad[3]}),
    .opad(haddr[3]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2020 (
    .do({open_n1599,open_n1600,open_n1601,haddr_pad[2]}),
    .opad(haddr[2]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2021 (
    .do({open_n1616,open_n1617,open_n1618,haddr_pad[1]}),
    .opad(haddr[1]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2022 (
    .do({open_n1633,open_n1634,open_n1635,haddr_pad[0]}),
    .opad(haddr[0]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2023 (
    .do({open_n1650,open_n1651,open_n1652,1'b0}),
    .opad(hburst[2]));  // ../../RTL/CPU/prv464_top.v(25)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2024 (
    .do({open_n1667,open_n1668,open_n1669,1'b0}),
    .opad(hburst[1]));  // ../../RTL/CPU/prv464_top.v(25)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2025 (
    .do({open_n1684,open_n1685,open_n1686,hburst_pad[0]}),
    .opad(hburst[0]));  // ../../RTL/CPU/prv464_top.v(25)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2026 (
    .do({open_n1701,open_n1702,open_n1703,1'b0}),
    .opad(hmastlock));  // ../../RTL/CPU/prv464_top.v(28)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2027 (
    .do({open_n1718,open_n1719,open_n1720,1'b0}),
    .opad(hprot[3]));  // ../../RTL/CPU/prv464_top.v(26)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2028 (
    .do({open_n1735,open_n1736,open_n1737,1'b0}),
    .opad(hprot[2]));  // ../../RTL/CPU/prv464_top.v(26)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2029 (
    .do({open_n1752,open_n1753,open_n1754,1'b1}),
    .opad(hprot[1]));  // ../../RTL/CPU/prv464_top.v(26)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2030 (
    .do({open_n1769,open_n1770,open_n1771,1'b1}),
    .opad(hprot[0]));  // ../../RTL/CPU/prv464_top.v(26)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2031 (
    .ipad(hrdata[63]),
    .di(hrdata_pad[63]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2032 (
    .ipad(hrdata[62]),
    .di(hrdata_pad[62]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2033 (
    .ipad(hrdata[61]),
    .di(hrdata_pad[61]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2034 (
    .ipad(hrdata[60]),
    .di(hrdata_pad[60]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2035 (
    .ipad(hrdata[59]),
    .di(hrdata_pad[59]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2036 (
    .ipad(hrdata[58]),
    .di(hrdata_pad[58]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2037 (
    .ipad(hrdata[57]),
    .di(hrdata_pad[57]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2038 (
    .ipad(hrdata[56]),
    .di(hrdata_pad[56]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2039 (
    .ipad(hrdata[55]),
    .di(hrdata_pad[55]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2040 (
    .ipad(hrdata[54]),
    .di(hrdata_pad[54]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2041 (
    .ipad(hrdata[53]),
    .di(hrdata_pad[53]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2042 (
    .ipad(hrdata[52]),
    .di(hrdata_pad[52]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2043 (
    .ipad(hrdata[51]),
    .di(hrdata_pad[51]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2044 (
    .ipad(hrdata[50]),
    .di(hrdata_pad[50]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2045 (
    .ipad(hrdata[49]),
    .di(hrdata_pad[49]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2046 (
    .ipad(hrdata[48]),
    .di(hrdata_pad[48]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2047 (
    .ipad(hrdata[47]),
    .di(hrdata_pad[47]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2048 (
    .ipad(hrdata[46]),
    .di(hrdata_pad[46]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2049 (
    .ipad(hrdata[45]),
    .di(hrdata_pad[45]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2050 (
    .ipad(hrdata[44]),
    .di(hrdata_pad[44]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2051 (
    .ipad(hrdata[43]),
    .di(hrdata_pad[43]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2052 (
    .ipad(hrdata[42]),
    .di(hrdata_pad[42]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2053 (
    .ipad(hrdata[41]),
    .di(hrdata_pad[41]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2054 (
    .ipad(hrdata[40]),
    .di(hrdata_pad[40]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2055 (
    .ipad(hrdata[39]),
    .di(hrdata_pad[39]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2056 (
    .ipad(hrdata[38]),
    .di(hrdata_pad[38]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2057 (
    .ipad(hrdata[37]),
    .di(hrdata_pad[37]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2058 (
    .ipad(hrdata[36]),
    .di(hrdata_pad[36]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2059 (
    .ipad(hrdata[35]),
    .di(hrdata_pad[35]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2060 (
    .ipad(hrdata[34]),
    .di(hrdata_pad[34]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2061 (
    .ipad(hrdata[33]),
    .di(hrdata_pad[33]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2062 (
    .ipad(hrdata[32]),
    .di(hrdata_pad[32]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2063 (
    .ipad(hrdata[31]),
    .di(hrdata_pad[31]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2064 (
    .ipad(hrdata[30]),
    .di(hrdata_pad[30]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2065 (
    .ipad(hrdata[29]),
    .di(hrdata_pad[29]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2066 (
    .ipad(hrdata[28]),
    .di(hrdata_pad[28]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2067 (
    .ipad(hrdata[27]),
    .di(hrdata_pad[27]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2068 (
    .ipad(hrdata[26]),
    .di(hrdata_pad[26]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2069 (
    .ipad(hrdata[25]),
    .di(hrdata_pad[25]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2070 (
    .ipad(hrdata[24]),
    .di(hrdata_pad[24]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2071 (
    .ipad(hrdata[23]),
    .di(hrdata_pad[23]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2072 (
    .ipad(hrdata[22]),
    .di(hrdata_pad[22]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2073 (
    .ipad(hrdata[21]),
    .di(hrdata_pad[21]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2074 (
    .ipad(hrdata[20]),
    .di(hrdata_pad[20]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2075 (
    .ipad(hrdata[19]),
    .di(hrdata_pad[19]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2076 (
    .ipad(hrdata[18]),
    .di(hrdata_pad[18]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2077 (
    .ipad(hrdata[17]),
    .di(hrdata_pad[17]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2078 (
    .ipad(hrdata[16]),
    .di(hrdata_pad[16]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2079 (
    .ipad(hrdata[15]),
    .di(hrdata_pad[15]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2080 (
    .ipad(hrdata[14]),
    .di(hrdata_pad[14]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2081 (
    .ipad(hrdata[13]),
    .di(hrdata_pad[13]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2082 (
    .ipad(hrdata[12]),
    .di(hrdata_pad[12]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2083 (
    .ipad(hrdata[11]),
    .di(hrdata_pad[11]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2084 (
    .ipad(hrdata[10]),
    .di(hrdata_pad[10]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2085 (
    .ipad(hrdata[9]),
    .di(hrdata_pad[9]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2086 (
    .ipad(hrdata[8]),
    .di(hrdata_pad[8]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2087 (
    .ipad(hrdata[7]),
    .di(hrdata_pad[7]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2088 (
    .ipad(hrdata[6]),
    .di(hrdata_pad[6]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2089 (
    .ipad(hrdata[5]),
    .di(hrdata_pad[5]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2090 (
    .ipad(hrdata[4]),
    .di(hrdata_pad[4]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2091 (
    .ipad(hrdata[3]),
    .di(hrdata_pad[3]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2092 (
    .ipad(hrdata[2]),
    .di(hrdata_pad[2]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2093 (
    .ipad(hrdata[1]),
    .di(hrdata_pad[1]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2094 (
    .ipad(hrdata[0]),
    .di(hrdata_pad[0]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2095 (
    .ipad(hready),
    .di(hready_pad));  // ../../RTL/CPU/prv464_top.v(31)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2096 (
    .ipad(hreset_n));  // ../../RTL/CPU/prv464_top.v(33)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2097 (
    .ipad(hresp),
    .di(hresp_pad));  // ../../RTL/CPU/prv464_top.v(32)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2098 (
    .do({open_n2926,open_n2927,open_n2928,1'b0}),
    .opad(hsize[2]));  // ../../RTL/CPU/prv464_top.v(24)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2099 (
    .do({open_n2943,open_n2944,open_n2945,hsize_pad[1]}),
    .opad(hsize[1]));  // ../../RTL/CPU/prv464_top.v(24)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2100 (
    .do({open_n2960,open_n2961,open_n2962,hsize_pad[0]}),
    .opad(hsize[0]));  // ../../RTL/CPU/prv464_top.v(24)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2101 (
    .do({open_n2977,open_n2978,open_n2979,htrans_pad[1]}),
    .opad(htrans[1]));  // ../../RTL/CPU/prv464_top.v(27)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2102 (
    .do({open_n2994,open_n2995,open_n2996,htrans_pad[0]}),
    .opad(htrans[0]));  // ../../RTL/CPU/prv464_top.v(27)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2103 (
    .do({open_n3011,open_n3012,open_n3013,hwdata_pad[63]}),
    .opad(hwdata[63]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2104 (
    .do({open_n3028,open_n3029,open_n3030,hwdata_pad[62]}),
    .opad(hwdata[62]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2105 (
    .do({open_n3045,open_n3046,open_n3047,hwdata_pad[61]}),
    .opad(hwdata[61]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2106 (
    .do({open_n3062,open_n3063,open_n3064,hwdata_pad[60]}),
    .opad(hwdata[60]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2107 (
    .do({open_n3079,open_n3080,open_n3081,hwdata_pad[59]}),
    .opad(hwdata[59]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2108 (
    .do({open_n3096,open_n3097,open_n3098,hwdata_pad[58]}),
    .opad(hwdata[58]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2109 (
    .do({open_n3113,open_n3114,open_n3115,hwdata_pad[57]}),
    .opad(hwdata[57]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2110 (
    .do({open_n3130,open_n3131,open_n3132,hwdata_pad[56]}),
    .opad(hwdata[56]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2111 (
    .do({open_n3147,open_n3148,open_n3149,hwdata_pad[55]}),
    .opad(hwdata[55]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2112 (
    .do({open_n3164,open_n3165,open_n3166,hwdata_pad[54]}),
    .opad(hwdata[54]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2113 (
    .do({open_n3181,open_n3182,open_n3183,hwdata_pad[53]}),
    .opad(hwdata[53]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2114 (
    .do({open_n3198,open_n3199,open_n3200,hwdata_pad[52]}),
    .opad(hwdata[52]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2115 (
    .do({open_n3215,open_n3216,open_n3217,hwdata_pad[51]}),
    .opad(hwdata[51]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2116 (
    .do({open_n3232,open_n3233,open_n3234,hwdata_pad[50]}),
    .opad(hwdata[50]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2117 (
    .do({open_n3249,open_n3250,open_n3251,hwdata_pad[49]}),
    .opad(hwdata[49]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2118 (
    .do({open_n3266,open_n3267,open_n3268,hwdata_pad[48]}),
    .opad(hwdata[48]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2119 (
    .do({open_n3283,open_n3284,open_n3285,hwdata_pad[47]}),
    .opad(hwdata[47]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2120 (
    .do({open_n3300,open_n3301,open_n3302,hwdata_pad[46]}),
    .opad(hwdata[46]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2121 (
    .do({open_n3317,open_n3318,open_n3319,hwdata_pad[45]}),
    .opad(hwdata[45]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2122 (
    .do({open_n3334,open_n3335,open_n3336,hwdata_pad[44]}),
    .opad(hwdata[44]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2123 (
    .do({open_n3351,open_n3352,open_n3353,hwdata_pad[43]}),
    .opad(hwdata[43]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2124 (
    .do({open_n3368,open_n3369,open_n3370,hwdata_pad[42]}),
    .opad(hwdata[42]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2125 (
    .do({open_n3385,open_n3386,open_n3387,hwdata_pad[41]}),
    .opad(hwdata[41]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2126 (
    .do({open_n3402,open_n3403,open_n3404,hwdata_pad[40]}),
    .opad(hwdata[40]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2127 (
    .do({open_n3419,open_n3420,open_n3421,hwdata_pad[39]}),
    .opad(hwdata[39]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2128 (
    .do({open_n3436,open_n3437,open_n3438,hwdata_pad[38]}),
    .opad(hwdata[38]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2129 (
    .do({open_n3453,open_n3454,open_n3455,hwdata_pad[37]}),
    .opad(hwdata[37]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2130 (
    .do({open_n3470,open_n3471,open_n3472,hwdata_pad[36]}),
    .opad(hwdata[36]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2131 (
    .do({open_n3487,open_n3488,open_n3489,hwdata_pad[35]}),
    .opad(hwdata[35]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2132 (
    .do({open_n3504,open_n3505,open_n3506,hwdata_pad[34]}),
    .opad(hwdata[34]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2133 (
    .do({open_n3521,open_n3522,open_n3523,hwdata_pad[33]}),
    .opad(hwdata[33]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2134 (
    .do({open_n3538,open_n3539,open_n3540,hwdata_pad[32]}),
    .opad(hwdata[32]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2135 (
    .do({open_n3555,open_n3556,open_n3557,hwdata_pad[31]}),
    .opad(hwdata[31]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2136 (
    .do({open_n3572,open_n3573,open_n3574,hwdata_pad[30]}),
    .opad(hwdata[30]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2137 (
    .do({open_n3589,open_n3590,open_n3591,hwdata_pad[29]}),
    .opad(hwdata[29]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2138 (
    .do({open_n3606,open_n3607,open_n3608,hwdata_pad[28]}),
    .opad(hwdata[28]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2139 (
    .do({open_n3623,open_n3624,open_n3625,hwdata_pad[27]}),
    .opad(hwdata[27]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2140 (
    .do({open_n3640,open_n3641,open_n3642,hwdata_pad[26]}),
    .opad(hwdata[26]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2141 (
    .do({open_n3657,open_n3658,open_n3659,hwdata_pad[25]}),
    .opad(hwdata[25]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2142 (
    .do({open_n3674,open_n3675,open_n3676,hwdata_pad[24]}),
    .opad(hwdata[24]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2143 (
    .do({open_n3691,open_n3692,open_n3693,hwdata_pad[23]}),
    .opad(hwdata[23]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2144 (
    .do({open_n3708,open_n3709,open_n3710,hwdata_pad[22]}),
    .opad(hwdata[22]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2145 (
    .do({open_n3725,open_n3726,open_n3727,hwdata_pad[21]}),
    .opad(hwdata[21]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2146 (
    .do({open_n3742,open_n3743,open_n3744,hwdata_pad[20]}),
    .opad(hwdata[20]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2147 (
    .do({open_n3759,open_n3760,open_n3761,hwdata_pad[19]}),
    .opad(hwdata[19]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2148 (
    .do({open_n3776,open_n3777,open_n3778,hwdata_pad[18]}),
    .opad(hwdata[18]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2149 (
    .do({open_n3793,open_n3794,open_n3795,hwdata_pad[17]}),
    .opad(hwdata[17]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2150 (
    .do({open_n3810,open_n3811,open_n3812,hwdata_pad[16]}),
    .opad(hwdata[16]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2151 (
    .do({open_n3827,open_n3828,open_n3829,hwdata_pad[15]}),
    .opad(hwdata[15]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2152 (
    .do({open_n3844,open_n3845,open_n3846,hwdata_pad[14]}),
    .opad(hwdata[14]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2153 (
    .do({open_n3861,open_n3862,open_n3863,hwdata_pad[13]}),
    .opad(hwdata[13]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2154 (
    .do({open_n3878,open_n3879,open_n3880,hwdata_pad[12]}),
    .opad(hwdata[12]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2155 (
    .do({open_n3895,open_n3896,open_n3897,hwdata_pad[11]}),
    .opad(hwdata[11]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2156 (
    .do({open_n3912,open_n3913,open_n3914,hwdata_pad[10]}),
    .opad(hwdata[10]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2157 (
    .do({open_n3929,open_n3930,open_n3931,hwdata_pad[9]}),
    .opad(hwdata[9]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2158 (
    .do({open_n3946,open_n3947,open_n3948,hwdata_pad[8]}),
    .opad(hwdata[8]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2159 (
    .do({open_n3963,open_n3964,open_n3965,hwdata_pad[7]}),
    .opad(hwdata[7]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2160 (
    .do({open_n3980,open_n3981,open_n3982,hwdata_pad[6]}),
    .opad(hwdata[6]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2161 (
    .do({open_n3997,open_n3998,open_n3999,hwdata_pad[5]}),
    .opad(hwdata[5]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2162 (
    .do({open_n4014,open_n4015,open_n4016,hwdata_pad[4]}),
    .opad(hwdata[4]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2163 (
    .do({open_n4031,open_n4032,open_n4033,hwdata_pad[3]}),
    .opad(hwdata[3]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2164 (
    .do({open_n4048,open_n4049,open_n4050,hwdata_pad[2]}),
    .opad(hwdata[2]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2165 (
    .do({open_n4065,open_n4066,open_n4067,hwdata_pad[1]}),
    .opad(hwdata[1]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2166 (
    .do({open_n4082,open_n4083,open_n4084,hwdata_pad[0]}),
    .opad(hwdata[0]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2167 (
    .do({open_n4099,open_n4100,open_n4101,hwrite_pad}),
    .opad(hwrite));  // ../../RTL/CPU/prv464_top.v(23)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2168 (
    .ipad(mtime[63]),
    .di(mtime_pad[63]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2169 (
    .ipad(mtime[62]),
    .di(mtime_pad[62]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2170 (
    .ipad(mtime[61]),
    .di(mtime_pad[61]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2171 (
    .ipad(mtime[60]),
    .di(mtime_pad[60]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2172 (
    .ipad(mtime[59]),
    .di(mtime_pad[59]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2173 (
    .ipad(mtime[58]),
    .di(mtime_pad[58]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2174 (
    .ipad(mtime[57]),
    .di(mtime_pad[57]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2175 (
    .ipad(mtime[56]),
    .di(mtime_pad[56]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2176 (
    .ipad(mtime[55]),
    .di(mtime_pad[55]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2177 (
    .ipad(mtime[54]),
    .di(mtime_pad[54]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2178 (
    .ipad(mtime[53]),
    .di(mtime_pad[53]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2179 (
    .ipad(mtime[52]),
    .di(mtime_pad[52]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2180 (
    .ipad(mtime[51]),
    .di(mtime_pad[51]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2181 (
    .ipad(mtime[50]),
    .di(mtime_pad[50]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2182 (
    .ipad(mtime[49]),
    .di(mtime_pad[49]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2183 (
    .ipad(mtime[48]),
    .di(mtime_pad[48]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2184 (
    .ipad(mtime[47]),
    .di(mtime_pad[47]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2185 (
    .ipad(mtime[46]),
    .di(mtime_pad[46]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2186 (
    .ipad(mtime[45]),
    .di(mtime_pad[45]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2187 (
    .ipad(mtime[44]),
    .di(mtime_pad[44]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2188 (
    .ipad(mtime[43]),
    .di(mtime_pad[43]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2189 (
    .ipad(mtime[42]),
    .di(mtime_pad[42]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2190 (
    .ipad(mtime[41]),
    .di(mtime_pad[41]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2191 (
    .ipad(mtime[40]),
    .di(mtime_pad[40]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2192 (
    .ipad(mtime[39]),
    .di(mtime_pad[39]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2193 (
    .ipad(mtime[38]),
    .di(mtime_pad[38]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2194 (
    .ipad(mtime[37]),
    .di(mtime_pad[37]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2195 (
    .ipad(mtime[36]),
    .di(mtime_pad[36]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2196 (
    .ipad(mtime[35]),
    .di(mtime_pad[35]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2197 (
    .ipad(mtime[34]),
    .di(mtime_pad[34]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2198 (
    .ipad(mtime[33]),
    .di(mtime_pad[33]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2199 (
    .ipad(mtime[32]),
    .di(mtime_pad[32]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2200 (
    .ipad(mtime[31]),
    .di(mtime_pad[31]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2201 (
    .ipad(mtime[30]),
    .di(mtime_pad[30]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2202 (
    .ipad(mtime[29]),
    .di(mtime_pad[29]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2203 (
    .ipad(mtime[28]),
    .di(mtime_pad[28]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2204 (
    .ipad(mtime[27]),
    .di(mtime_pad[27]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2205 (
    .ipad(mtime[26]),
    .di(mtime_pad[26]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2206 (
    .ipad(mtime[25]),
    .di(mtime_pad[25]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2207 (
    .ipad(mtime[24]),
    .di(mtime_pad[24]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2208 (
    .ipad(mtime[23]),
    .di(mtime_pad[23]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2209 (
    .ipad(mtime[22]),
    .di(mtime_pad[22]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2210 (
    .ipad(mtime[21]),
    .di(mtime_pad[21]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2211 (
    .ipad(mtime[20]),
    .di(mtime_pad[20]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2212 (
    .ipad(mtime[19]),
    .di(mtime_pad[19]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2213 (
    .ipad(mtime[18]),
    .di(mtime_pad[18]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2214 (
    .ipad(mtime[17]),
    .di(mtime_pad[17]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2215 (
    .ipad(mtime[16]),
    .di(mtime_pad[16]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2216 (
    .ipad(mtime[15]),
    .di(mtime_pad[15]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2217 (
    .ipad(mtime[14]),
    .di(mtime_pad[14]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2218 (
    .ipad(mtime[13]),
    .di(mtime_pad[13]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2219 (
    .ipad(mtime[12]),
    .di(mtime_pad[12]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2220 (
    .ipad(mtime[11]),
    .di(mtime_pad[11]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2221 (
    .ipad(mtime[10]),
    .di(mtime_pad[10]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2222 (
    .ipad(mtime[9]),
    .di(mtime_pad[9]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2223 (
    .ipad(mtime[8]),
    .di(mtime_pad[8]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2224 (
    .ipad(mtime[7]),
    .di(mtime_pad[7]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2225 (
    .ipad(mtime[6]),
    .di(mtime_pad[6]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2226 (
    .ipad(mtime[5]),
    .di(mtime_pad[5]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2227 (
    .ipad(mtime[4]),
    .di(mtime_pad[4]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2228 (
    .ipad(mtime[3]),
    .di(mtime_pad[3]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2229 (
    .ipad(mtime[2]),
    .di(mtime_pad[2]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2230 (
    .ipad(mtime[1]),
    .di(mtime_pad[1]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2231 (
    .ipad(mtime[0]),
    .di(mtime_pad[0]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2232 (
    .ipad(rst),
    .di(rst_pad));  // ../../RTL/CPU/prv464_top.v(20)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2233 (
    .ipad(s_ext_int),
    .di(s_ext_int_pad));  // ../../RTL/CPU/prv464_top.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(C@D)"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(C@D)"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000111111110000),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000111111110000),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2592|_al_u2652  (
    .c({ds2[0],ds2[63]}),
    .d({rd_data_sub,rd_data_sub}),
    .f({\exu/alu_au/n17 [0],\exu/alu_au/n17 [63]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2593|_al_u3906  (
    .a({open_n5265,\exu/alu_au/add_64 [1]}),
    .b({open_n5266,mem_csr_data_add}),
    .c({ds2[1],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[1]}),
    .f({\exu/alu_au/n17 [1],_al_u3906_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2594|_al_u3898  (
    .a({open_n5291,\exu/alu_au/add_64 [10]}),
    .b({open_n5292,mem_csr_data_add}),
    .c({ds2[10],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[10]}),
    .f({\exu/alu_au/n17 [10],_al_u3898_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2595|_al_u3890  (
    .a({open_n5317,\exu/alu_au/add_64 [11]}),
    .b({open_n5318,mem_csr_data_add}),
    .c({ds2[11],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[11]}),
    .f({\exu/alu_au/n17 [11],_al_u3890_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2596|_al_u3882  (
    .a({open_n5343,\exu/alu_au/add_64 [12]}),
    .b({open_n5344,mem_csr_data_add}),
    .c({ds2[12],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[12]}),
    .f({\exu/alu_au/n17 [12],_al_u3882_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2597|_al_u3874  (
    .a({open_n5365,\exu/alu_au/add_64 [13]}),
    .b({open_n5366,mem_csr_data_add}),
    .c({ds2[13],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[13]}),
    .f({\exu/alu_au/n17 [13],_al_u3874_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2598|_al_u3866  (
    .a({open_n5387,\exu/alu_au/add_64 [14]}),
    .b({open_n5388,mem_csr_data_add}),
    .c({ds2[14],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[14]}),
    .f({\exu/alu_au/n17 [14],_al_u3866_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2599|_al_u3859  (
    .a({open_n5413,\exu/alu_au/add_64 [15]}),
    .b({open_n5414,mem_csr_data_add}),
    .c({ds2[15],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[15]}),
    .f({\exu/alu_au/n17 [15],_al_u3859_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2600|_al_u3852  (
    .a({open_n5435,\exu/alu_au/add_64 [16]}),
    .b({open_n5436,mem_csr_data_add}),
    .c({ds2[16],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[16]}),
    .f({\exu/alu_au/n17 [16],_al_u3852_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2601|_al_u3845  (
    .a({open_n5457,\exu/alu_au/add_64 [17]}),
    .b({open_n5458,mem_csr_data_add}),
    .c({ds2[17],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[17]}),
    .f({\exu/alu_au/n17 [17],_al_u3845_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2602|_al_u3838  (
    .a({open_n5483,\exu/alu_au/add_64 [18]}),
    .b({open_n5484,mem_csr_data_add}),
    .c({ds2[18],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[18]}),
    .f({\exu/alu_au/n17 [18],_al_u3838_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2603|_al_u3831  (
    .a({open_n5509,\exu/alu_au/add_64 [19]}),
    .b({open_n5510,mem_csr_data_add}),
    .c({ds2[19],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[19]}),
    .f({\exu/alu_au/n17 [19],_al_u3831_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2604|_al_u3824  (
    .a({open_n5531,\exu/alu_au/add_64 [2]}),
    .b({open_n5532,mem_csr_data_add}),
    .c({ds2[2],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[2]}),
    .f({\exu/alu_au/n17 [2],_al_u3824_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2605|_al_u3817  (
    .a({open_n5553,\exu/alu_au/add_64 [20]}),
    .b({open_n5554,mem_csr_data_add}),
    .c({ds2[20],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[20]}),
    .f({\exu/alu_au/n17 [20],_al_u3817_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2606|_al_u3810  (
    .a({open_n5579,\exu/alu_au/add_64 [21]}),
    .b({open_n5580,mem_csr_data_add}),
    .c({ds2[21],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[21]}),
    .f({\exu/alu_au/n17 [21],_al_u3810_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2607|_al_u3803  (
    .a({open_n5605,\exu/alu_au/add_64 [22]}),
    .b({open_n5606,mem_csr_data_add}),
    .c({ds2[22],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[22]}),
    .f({\exu/alu_au/n17 [22],_al_u3803_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2608|_al_u3796  (
    .a({open_n5627,\exu/alu_au/add_64 [23]}),
    .b({open_n5628,mem_csr_data_add}),
    .c({ds2[23],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[23]}),
    .f({\exu/alu_au/n17 [23],_al_u3796_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2609|_al_u3789  (
    .a({open_n5649,\exu/alu_au/add_64 [24]}),
    .b({open_n5650,mem_csr_data_add}),
    .c({ds2[24],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[24]}),
    .f({\exu/alu_au/n17 [24],_al_u3789_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2610|_al_u3782  (
    .a({open_n5675,\exu/alu_au/add_64 [25]}),
    .b({open_n5676,mem_csr_data_add}),
    .c({ds2[25],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[25]}),
    .f({\exu/alu_au/n17 [25],_al_u3782_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2611|_al_u3775  (
    .a({open_n5701,\exu/alu_au/add_64 [26]}),
    .b({open_n5702,mem_csr_data_add}),
    .c({ds2[26],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[26]}),
    .f({\exu/alu_au/n17 [26],_al_u3775_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2612|_al_u3768  (
    .a({open_n5723,\exu/alu_au/add_64 [27]}),
    .b({open_n5724,mem_csr_data_add}),
    .c({ds2[27],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[27]}),
    .f({\exu/alu_au/n17 [27],_al_u3768_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2613|_al_u3761  (
    .a({open_n5745,\exu/alu_au/add_64 [28]}),
    .b({open_n5746,mem_csr_data_add}),
    .c({ds2[28],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[28]}),
    .f({\exu/alu_au/n17 [28],_al_u3761_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2614|_al_u3754  (
    .a({open_n5771,\exu/alu_au/add_64 [29]}),
    .b({open_n5772,mem_csr_data_add}),
    .c({ds2[29],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[29]}),
    .f({\exu/alu_au/n17 [29],_al_u3754_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2615|_al_u3747  (
    .a({open_n5797,\exu/alu_au/add_64 [3]}),
    .b({open_n5798,mem_csr_data_add}),
    .c({ds2[3],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[3]}),
    .f({\exu/alu_au/n17 [3],_al_u3747_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2616|_al_u3740  (
    .a({open_n5819,\exu/alu_au/add_64 [30]}),
    .b({open_n5820,mem_csr_data_add}),
    .c({ds2[30],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[30]}),
    .f({\exu/alu_au/n17 [30],_al_u3740_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2617|_al_u3733  (
    .a({open_n5841,\exu/alu_au/add_64 [31]}),
    .b({open_n5842,mem_csr_data_add}),
    .c({ds2[31],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[31]}),
    .f({\exu/alu_au/n17 [31],_al_u3733_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2618|_al_u3725  (
    .b({open_n5865,mem_csr_data_or}),
    .c({ds2[32],ds2[32]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [32],_al_u3725_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2619|_al_u3717  (
    .b({open_n5888,mem_csr_data_or}),
    .c({ds2[33],ds2[33]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [33],_al_u3717_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2620|_al_u3709  (
    .b({open_n5915,mem_csr_data_or}),
    .c({ds2[34],ds2[34]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [34],_al_u3709_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2621|_al_u3701  (
    .b({open_n5942,mem_csr_data_or}),
    .c({ds2[35],ds2[35]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [35],_al_u3701_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2622|_al_u3693  (
    .b({open_n5965,mem_csr_data_or}),
    .c({ds2[36],ds2[36]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [36],_al_u3693_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2623|_al_u3685  (
    .b({open_n5988,mem_csr_data_or}),
    .c({ds2[37],ds2[37]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [37],_al_u3685_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2624|_al_u3677  (
    .b({open_n6015,mem_csr_data_or}),
    .c({ds2[38],ds2[38]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [38],_al_u3677_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2625|_al_u3669  (
    .b({open_n6042,mem_csr_data_or}),
    .c({ds2[39],ds2[39]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [39],_al_u3669_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2626|_al_u3662  (
    .a({open_n6063,\exu/alu_au/add_64 [4]}),
    .b({open_n6064,mem_csr_data_add}),
    .c({ds2[4],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[4]}),
    .f({\exu/alu_au/n17 [4],_al_u3662_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2627|_al_u3654  (
    .b({open_n6091,mem_csr_data_or}),
    .c({ds2[40],ds2[40]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [40],_al_u3654_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2628|_al_u3646  (
    .b({open_n6114,mem_csr_data_or}),
    .c({ds2[41],ds2[41]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [41],_al_u3646_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2629|_al_u3638  (
    .b({open_n6141,mem_csr_data_or}),
    .c({ds2[42],ds2[42]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [42],_al_u3638_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2630|_al_u3630  (
    .b({open_n6168,mem_csr_data_or}),
    .c({ds2[43],ds2[43]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [43],_al_u3630_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2631|_al_u3622  (
    .b({open_n6191,mem_csr_data_or}),
    .c({ds2[44],ds2[44]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [44],_al_u3622_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2632|_al_u3614  (
    .b({open_n6214,mem_csr_data_or}),
    .c({ds2[45],ds2[45]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [45],_al_u3614_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2633|_al_u3606  (
    .b({open_n6241,mem_csr_data_or}),
    .c({ds2[46],ds2[46]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [46],_al_u3606_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2634|_al_u3598  (
    .b({open_n6268,mem_csr_data_or}),
    .c({ds2[47],ds2[47]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [47],_al_u3598_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2635|_al_u3590  (
    .b({open_n6291,mem_csr_data_or}),
    .c({ds2[48],ds2[48]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [48],_al_u3590_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2636|_al_u3582  (
    .b({open_n6314,mem_csr_data_or}),
    .c({ds2[49],ds2[49]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [49],_al_u3582_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2637|_al_u3575  (
    .a({open_n6339,\exu/alu_au/add_64 [5]}),
    .b({open_n6340,mem_csr_data_add}),
    .c({ds2[5],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[5]}),
    .f({\exu/alu_au/n17 [5],_al_u3575_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2638|_al_u3567  (
    .b({open_n6367,mem_csr_data_or}),
    .c({ds2[50],ds2[50]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [50],_al_u3567_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2639|_al_u3559  (
    .b({open_n6394,mem_csr_data_or}),
    .c({ds2[51],ds2[51]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [51],_al_u3559_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2640|_al_u3551  (
    .b({open_n6417,mem_csr_data_or}),
    .c({ds2[52],ds2[52]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [52],_al_u3551_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2641|_al_u3543  (
    .b({open_n6440,mem_csr_data_or}),
    .c({ds2[53],ds2[53]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [53],_al_u3543_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2642|_al_u3535  (
    .b({open_n6467,mem_csr_data_or}),
    .c({ds2[54],ds2[54]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [54],_al_u3535_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2643|_al_u3527  (
    .b({open_n6494,mem_csr_data_or}),
    .c({ds2[55],ds2[55]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [55],_al_u3527_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2644|_al_u3519  (
    .b({open_n6517,mem_csr_data_or}),
    .c({ds2[56],ds2[56]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [56],_al_u3519_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2645|_al_u3511  (
    .b({open_n6540,mem_csr_data_or}),
    .c({ds2[57],ds2[57]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [57],_al_u3511_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2646|_al_u3503  (
    .b({open_n6567,mem_csr_data_or}),
    .c({ds2[58],ds2[58]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [58],_al_u3503_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2647|_al_u3495  (
    .b({open_n6594,mem_csr_data_or}),
    .c({ds2[59],ds2[59]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [59],_al_u3495_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2648|_al_u3488  (
    .a({open_n6615,\exu/alu_au/add_64 [6]}),
    .b({open_n6616,mem_csr_data_add}),
    .c({ds2[6],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[6]}),
    .f({\exu/alu_au/n17 [6],_al_u3488_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2649|_al_u3480  (
    .b({open_n6639,mem_csr_data_or}),
    .c({ds2[60],ds2[60]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [60],_al_u3480_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2650|_al_u3472  (
    .b({open_n6662,mem_csr_data_or}),
    .c({ds2[61],ds2[61]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [61],_al_u3472_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2651|_al_u3464  (
    .b({open_n6689,mem_csr_data_or}),
    .c({ds2[62],ds2[62]}),
    .d({rd_data_sub,mem_csr_data_ds2}),
    .f({\exu/alu_au/n17 [62],_al_u3464_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2653|_al_u3449  (
    .a({open_n6714,\exu/alu_au/add_64 [7]}),
    .b({open_n6715,mem_csr_data_add}),
    .c({ds2[7],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[7]}),
    .f({\exu/alu_au/n17 [7],_al_u3449_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*C)*~(B*A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(D*C)*~(B*A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b0000011101110111),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b0000011101110111),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2654|_al_u3441  (
    .a({open_n6736,\exu/alu_au/add_64 [8]}),
    .b({open_n6737,mem_csr_data_add}),
    .c({ds2[8],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[8]}),
    .f({\exu/alu_au/n17 [8],_al_u3441_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(C@D)"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"))
    \_al_u2655|_al_u3432  (
    .a({open_n6762,\exu/alu_au/add_64 [9]}),
    .b({open_n6763,mem_csr_data_add}),
    .c({ds2[9],mem_csr_data_ds2}),
    .d({rd_data_sub,ds2[9]}),
    .f({\exu/alu_au/n17 [9],_al_u3432_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0000001100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2659|ins_fetch/reg1_b31  (
    .a({ins_read[31],open_n6784}),
    .b({ins_read[63],ins_read[63]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[31]}),
    .sr(rst_pad),
    .f({_al_u2659_o,open_n6797}),
    .q({open_n6801,\ins_fetch/ins_hold [31]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2660|ins_dec/reg1_b11  (
    .c({\ins_fetch/ins_hold [31],_al_u2660_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({1'b0,_al_u2659_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u2660_o,id_ins[31]}),
    .q({open_n6821,ex_csr_index[11]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0000001100000101),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0000001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2662|ins_fetch/reg1_b30  (
    .a({ins_read[30],open_n6822}),
    .b({ins_read[62],ins_read[62]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[30]}),
    .sr(rst_pad),
    .f({_al_u2662_o,open_n6839}),
    .q({open_n6843,\ins_fetch/ins_hold [30]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2663|ins_dec/reg1_b10  (
    .c({\ins_fetch/ins_hold [30],_al_u2663_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({1'b0,_al_u2662_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u2663_o,id_ins[30]}),
    .q({open_n6867,ex_csr_index[10]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0000001100000101),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0000001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2667|ins_fetch/reg1_b27  (
    .a({ins_read[27],open_n6868}),
    .b({ins_read[59],ins_read[59]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[27]}),
    .sr(rst_pad),
    .f({_al_u2667_o,open_n6885}),
    .q({open_n6889,\ins_fetch/ins_hold [27]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0000001100000101),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0000001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2670|ins_fetch/reg1_b26  (
    .a({ins_read[26],open_n6890}),
    .b({ins_read[58],ins_read[58]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[26]}),
    .sr(rst_pad),
    .f({_al_u2670_o,open_n6907}),
    .q({open_n6911,\ins_fetch/ins_hold [26]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2671|ins_dec/reg1_b6  (
    .c({\ins_fetch/ins_hold [26],_al_u2671_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({1'b0,_al_u2670_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u2671_o,id_ins[26]}),
    .q({open_n6935,ex_csr_index[6]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0000001100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2674|ins_fetch/reg1_b24  (
    .a({ins_read[24],open_n6936}),
    .b({ins_read[56],ins_read[56]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[24]}),
    .sr(rst_pad),
    .f({_al_u2674_o,open_n6949}),
    .q({open_n6953,\ins_fetch/ins_hold [24]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0000001100000101),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0000001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2677|ins_fetch/reg1_b23  (
    .a({ins_read[23],open_n6954}),
    .b({ins_read[55],ins_read[55]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[23]}),
    .sr(rst_pad),
    .f({_al_u2677_o,open_n6971}),
    .q({open_n6975,\ins_fetch/ins_hold [23]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2678|ins_dec/reg1_b3  (
    .c({\ins_fetch/ins_hold [23],_al_u2678_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({1'b0,_al_u2677_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u2678_o,id_ins[23]}),
    .q({open_n6999,ex_csr_index[3]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0000001100000101),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0000001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2680|ins_fetch/reg1_b22  (
    .a({ins_read[22],open_n7000}),
    .b({ins_read[54],ins_read[54]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[22]}),
    .sr(rst_pad),
    .f({_al_u2680_o,open_n7017}),
    .q({open_n7021,\ins_fetch/ins_hold [22]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0000001100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2683|ins_fetch/reg1_b21  (
    .a({ins_read[21],open_n7022}),
    .b({ins_read[53],ins_read[53]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[21]}),
    .sr(rst_pad),
    .f({_al_u2683_o,open_n7035}),
    .q({open_n7039,\ins_fetch/ins_hold [21]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2684|ins_dec/reg1_b1  (
    .c({\ins_fetch/ins_hold [21],_al_u2684_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({1'b0,_al_u2683_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u2684_o,id_ins[21]}),
    .q({open_n7063,ex_csr_index[1]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(B*~(~D*~C*A))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1100110011000100),
    .MODE("LOGIC"))
    \_al_u2692|_al_u2694  (
    .a({_al_u2691_o,open_n7064}),
    .b({wb_gpr_write,open_n7065}),
    .c({wb_rd_index[0],\cu_ru/n52 [4]}),
    .d({wb_rd_index[1],\cu_ru/n53_lutinv }),
    .f({\cu_ru/n53_lutinv ,\cu_ru/n53_0_al_n1985 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2693|_al_u8586  (
    .b({open_n7088,data_rd[32]}),
    .c({\cu_ru/n52 [4],data_rd[33]}),
    .d({\cu_ru/n53_lutinv ,\exu/mux27_b32_sel_is_1_o }),
    .f({\cu_ru/n53_1_al_n1986 ,\exu/n57 [32]}));
  // ../../RTL/CPU/IF/ins_fetch.v(154)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("~(~C*D)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("~(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1111000011111111),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1111000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2696|ins_fetch/valid_reg  (
    .a({open_n7113,_al_u9189_o}),
    .b({open_n7114,_al_u9195_o}),
    .c({rst_pad,_al_u9268_o}),
    .ce(_al_n0_en),
    .clk(clk_pad),
    .d({_al_u2695_o,_al_u9264_o}),
    .sr(\ins_fetch/n25 ),
    .f({\ins_fetch/n25 ,\ins_fetch/n27 }),
    .q({open_n7134,id_valid}));  // ../../RTL/CPU/IF/ins_fetch.v(154)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*~B*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"))
    \_al_u2697|_al_u2698  (
    .b({\biu/bus_unit/mmu/statu [2],open_n7137}),
    .c({\biu/bus_unit/mmu/statu [3],\biu/bus_unit/mmu/statu [0]}),
    .d({\biu/bus_unit/mmu/statu [1],_al_u2697_o}),
    .f({_al_u2697_o,_al_u2698_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~B*~A)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(~D*C*~B*~A)"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b0000000000010000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000000000010000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2700|_al_u2915  (
    .a({\biu/bus_unit/mmu/statu [0],\biu/bus_unit/mmu/statu [0]}),
    .b({\biu/bus_unit/mmu/statu [1],\biu/bus_unit/mmu/statu [1]}),
    .c({\biu/bus_unit/mmu/statu [2],\biu/bus_unit/mmu/statu [2]}),
    .d({\biu/bus_unit/mmu/statu [3],\biu/bus_unit/mmu/statu [3]}),
    .f({\biu/bus_unit/mmu/n37_lutinv ,_al_u2915_o}));
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2701|biu/bus_unit/mmu/reg3_b3  (
    .a({open_n7182,_al_u2963_o}),
    .b({open_n7183,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [3],\biu/bus_unit/mmu_hwdata [3]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [1],hrdata_pad[3]}),
    .sr(rst_pad),
    .f({\biu/bus_unit/mmu/n39 [0],open_n7201}),
    .q({open_n7205,\biu/bus_unit/mmu_hwdata [3]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2702|biu/bus_unit/mmu/reg3_b2  (
    .a({open_n7206,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/n39 [0],\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [2],\biu/bus_unit/mmu_hwdata [2]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu/n37_lutinv ,hrdata_pad[2]}),
    .sr(rst_pad),
    .f({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,open_n7220}),
    .q({open_n7224,\biu/bus_unit/mmu_hwdata [2]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u2703|_al_u2955  (
    .b({open_n7227,\biu/bus_unit/statu [3]}),
    .c({\biu/bus_unit/statu [4],\biu/bus_unit/statu [4]}),
    .d({\biu/bus_unit/statu [2],\biu/bus_unit/statu [2]}),
    .f({_al_u2703_o,_al_u2955_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(~C*~B*D)"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"))
    \_al_u2704|_al_u3409  (
    .a({open_n7248,_al_u2703_o}),
    .b(\biu/bus_unit/statu [1:0]),
    .c({\biu/bus_unit/statu [3],\biu/bus_unit/statu [1]}),
    .d({_al_u2703_o,\biu/bus_unit/statu [3]}),
    .f({_al_u2704_o,\biu/bus_unit/n45_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*~B*A)"),
    //.LUTF1("(~D*C*~B*A)"),
    //.LUTG0("(D*C*~B*A)"),
    //.LUTG1("(~D*C*~B*A)"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0000000000100000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2706|_al_u2951  (
    .a({_al_u2703_o,_al_u2703_o}),
    .b({\biu/bus_unit/statu [0],\biu/bus_unit/statu [0]}),
    .c({\biu/bus_unit/statu [1],\biu/bus_unit/statu [1]}),
    .d({\biu/bus_unit/statu [3],\biu/bus_unit/statu [3]}),
    .f({_al_u2706_o,htrans_pad[0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*~A)"),
    //.LUT1("(~D*C*~B*A)"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"))
    \_al_u2707|_al_u2964  (
    .a({\biu/bus_unit/mmu/statu [0],\biu/bus_unit/mmu/statu [0]}),
    .b({\biu/bus_unit/mmu/statu [1],\biu/bus_unit/mmu/statu [1]}),
    .c({\biu/bus_unit/mmu/statu [2],\biu/bus_unit/mmu/statu [2]}),
    .d({\biu/bus_unit/mmu/statu [3],\biu/bus_unit/mmu/statu [3]}),
    .f({_al_u2707_o,_al_u2964_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2784|biu/cache_ctrl_logic/reg6_b119  (
    .a({open_n7313,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [52],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [119],\biu/paddress [119]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [53]}),
    .mi({open_n7324,\biu/paddress [119]}),
    .sr(rst_pad),
    .f({haddr_pad[55],_al_u3044_o}),
    .q({open_n7328,\biu/cache_ctrl_logic/pa_temp [119]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2785|biu/cache_ctrl_logic/reg6_b118  (
    .a({open_n7329,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [51],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [118],\biu/paddress [118]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [52]}),
    .mi({open_n7340,\biu/paddress [118]}),
    .sr(rst_pad),
    .f({haddr_pad[54],_al_u3047_o}),
    .q({open_n7344,\biu/cache_ctrl_logic/pa_temp [118]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2786|biu/cache_ctrl_logic/reg6_b117  (
    .a({open_n7345,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [50],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [117],\biu/paddress [117]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [51]}),
    .mi({open_n7349,\biu/paddress [117]}),
    .sr(rst_pad),
    .f({haddr_pad[53],_al_u3050_o}),
    .q({open_n7364,\biu/cache_ctrl_logic/pa_temp [117]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2787|biu/bus_unit/mmu/reg2_b52  (
    .b({\biu/bus_unit/n49 [49],open_n7367}),
    .c({\biu/paddress [116],_al_u3053_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3052_o}),
    .sr(rst_pad),
    .f({haddr_pad[52],open_n7385}),
    .q({open_n7389,\biu/paddress [116]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2788|biu/bus_unit/mmu/reg2_b51  (
    .b({\biu/bus_unit/n49 [48],open_n7392}),
    .c({\biu/paddress [115],_al_u3056_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3055_o}),
    .sr(rst_pad),
    .f({haddr_pad[51],open_n7410}),
    .q({open_n7414,\biu/paddress [115]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2789|biu/bus_unit/mmu/reg2_b50  (
    .b({\biu/bus_unit/n49 [47],open_n7417}),
    .c({\biu/paddress [114],_al_u3059_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3058_o}),
    .sr(rst_pad),
    .f({haddr_pad[50],open_n7431}),
    .q({open_n7435,\biu/paddress [114]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2791|biu/bus_unit/mmu/reg2_b49  (
    .b({\biu/bus_unit/n49 [46],open_n7438}),
    .c({\biu/paddress [113],_al_u3062_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3061_o}),
    .sr(rst_pad),
    .f({haddr_pad[49],open_n7452}),
    .q({open_n7456,\biu/paddress [113]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2792|biu/bus_unit/mmu/reg2_b48  (
    .b({\biu/bus_unit/n49 [45],open_n7459}),
    .c({\biu/paddress [112],_al_u3065_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3064_o}),
    .sr(rst_pad),
    .f({haddr_pad[48],open_n7477}),
    .q({open_n7481,\biu/paddress [112]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2793|biu/bus_unit/mmu/reg2_b47  (
    .b({\biu/bus_unit/n49 [44],open_n7484}),
    .c({\biu/paddress [111],_al_u3068_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3067_o}),
    .sr(rst_pad),
    .f({haddr_pad[47],open_n7502}),
    .q({open_n7506,\biu/paddress [111]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2794|biu/bus_unit/mmu/reg2_b46  (
    .b({\biu/bus_unit/n49 [43],open_n7509}),
    .c({\biu/paddress [110],_al_u3071_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3070_o}),
    .sr(rst_pad),
    .f({haddr_pad[46],open_n7523}),
    .q({open_n7527,\biu/paddress [110]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2795|biu/bus_unit/mmu/reg2_b45  (
    .b({\biu/bus_unit/n49 [42],open_n7530}),
    .c({\biu/paddress [109],_al_u3074_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3073_o}),
    .sr(rst_pad),
    .f({haddr_pad[45],open_n7544}),
    .q({open_n7548,\biu/paddress [109]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2796|biu/bus_unit/mmu/reg2_b44  (
    .b({\biu/bus_unit/n49 [41],open_n7551}),
    .c({\biu/paddress [108],_al_u3077_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3076_o}),
    .sr(rst_pad),
    .f({haddr_pad[44],open_n7569}),
    .q({open_n7573,\biu/paddress [108]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2797|biu/bus_unit/mmu/reg2_b43  (
    .b({\biu/bus_unit/n49 [40],open_n7576}),
    .c({\biu/paddress [107],_al_u3080_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3079_o}),
    .sr(rst_pad),
    .f({haddr_pad[43],open_n7594}),
    .q({open_n7598,\biu/paddress [107]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2798|biu/bus_unit/mmu/reg2_b42  (
    .b({\biu/bus_unit/n49 [39],open_n7601}),
    .c({\biu/paddress [106],_al_u3083_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3082_o}),
    .sr(rst_pad),
    .f({haddr_pad[42],open_n7615}),
    .q({open_n7619,\biu/paddress [106]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2799|biu/bus_unit/mmu/reg2_b41  (
    .b({\biu/bus_unit/n49 [38],open_n7622}),
    .c({\biu/paddress [105],_al_u3086_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3085_o}),
    .sr(rst_pad),
    .f({haddr_pad[41],open_n7636}),
    .q({open_n7640,\biu/paddress [105]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2800|biu/bus_unit/mmu/reg2_b40  (
    .b({\biu/bus_unit/n49 [37],open_n7643}),
    .c({\biu/paddress [104],_al_u3089_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3088_o}),
    .sr(rst_pad),
    .f({haddr_pad[40],open_n7661}),
    .q({open_n7665,\biu/paddress [104]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2802|biu/bus_unit/mmu/reg2_b39  (
    .b({\biu/bus_unit/n49 [36],open_n7668}),
    .c({\biu/paddress [103],_al_u3092_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3091_o}),
    .sr(rst_pad),
    .f({haddr_pad[39],open_n7686}),
    .q({open_n7690,\biu/paddress [103]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2803|biu/bus_unit/mmu/reg2_b38  (
    .b({\biu/bus_unit/n49 [35],open_n7693}),
    .c({\biu/paddress [102],_al_u3095_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3094_o}),
    .sr(rst_pad),
    .f({haddr_pad[38],open_n7707}),
    .q({open_n7711,\biu/paddress [102]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2804|biu/bus_unit/mmu/reg2_b37  (
    .b({\biu/bus_unit/n49 [34],open_n7714}),
    .c({\biu/paddress [101],_al_u3098_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3097_o}),
    .sr(rst_pad),
    .f({haddr_pad[37],open_n7728}),
    .q({open_n7732,\biu/paddress [101]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2805|biu/bus_unit/mmu/reg2_b36  (
    .b({\biu/bus_unit/n49 [33],open_n7735}),
    .c({\biu/paddress [100],_al_u3101_o}),
    .clk(clk_pad),
    .d({_al_u2705_o,_al_u3100_o}),
    .sr(rst_pad),
    .f({haddr_pad[36],open_n7753}),
    .q({open_n7757,\biu/paddress [100]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2806|biu/cache_ctrl_logic/reg6_b99  (
    .a({open_n7758,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [32],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [99],\biu/paddress [99]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [33]}),
    .mi({open_n7769,\biu/paddress [99]}),
    .sr(rst_pad),
    .f({haddr_pad[35],_al_u3104_o}),
    .q({open_n7773,\biu/cache_ctrl_logic/pa_temp [99]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2807|biu/cache_ctrl_logic/reg6_b98  (
    .a({open_n7774,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [31],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [98],\biu/paddress [98]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [32]}),
    .mi({open_n7785,\biu/paddress [98]}),
    .sr(rst_pad),
    .f({haddr_pad[34],_al_u3107_o}),
    .q({open_n7789,\biu/cache_ctrl_logic/pa_temp [98]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2808|biu/cache_ctrl_logic/reg6_b97  (
    .a({open_n7790,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [30],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [97],\biu/paddress [97]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [31]}),
    .mi({open_n7794,\biu/paddress [97]}),
    .sr(rst_pad),
    .f({haddr_pad[33],_al_u3110_o}),
    .q({open_n7809,\biu/cache_ctrl_logic/pa_temp [97]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2809|biu/cache_ctrl_logic/reg6_b96  (
    .a({open_n7810,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [29],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [96],\biu/paddress [96]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [30]}),
    .mi({open_n7814,\biu/paddress [96]}),
    .sr(rst_pad),
    .f({haddr_pad[32],_al_u3113_o}),
    .q({open_n7829,\biu/cache_ctrl_logic/pa_temp [96]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2810|biu/cache_ctrl_logic/reg6_b95  (
    .a({open_n7830,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [28],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [95],\biu/paddress [95]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [29]}),
    .mi({open_n7841,\biu/paddress [95]}),
    .sr(rst_pad),
    .f({haddr_pad[31],_al_u3116_o}),
    .q({open_n7845,\biu/cache_ctrl_logic/pa_temp [95]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2811|biu/cache_ctrl_logic/reg6_b94  (
    .a({open_n7846,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [27],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [94],\biu/paddress [94]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [28]}),
    .mi({open_n7857,\biu/paddress [94]}),
    .sr(rst_pad),
    .f({haddr_pad[30],_al_u3119_o}),
    .q({open_n7861,\biu/cache_ctrl_logic/pa_temp [94]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2813|biu/cache_ctrl_logic/reg6_b93  (
    .a({open_n7862,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [26],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [93],\biu/paddress [93]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [27]}),
    .mi({open_n7866,\biu/paddress [93]}),
    .sr(rst_pad),
    .f({haddr_pad[29],_al_u3122_o}),
    .q({open_n7881,\biu/cache_ctrl_logic/pa_temp [93]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2814|biu/cache_ctrl_logic/reg6_b92  (
    .a({open_n7882,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [25],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [92],\biu/paddress [92]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [26]}),
    .mi({open_n7886,\biu/paddress [92]}),
    .sr(rst_pad),
    .f({haddr_pad[28],_al_u3125_o}),
    .q({open_n7901,\biu/cache_ctrl_logic/pa_temp [92]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2815|biu/cache_ctrl_logic/reg6_b91  (
    .a({open_n7902,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [24],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [91],\biu/paddress [91]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [25]}),
    .mi({open_n7913,\biu/paddress [91]}),
    .sr(rst_pad),
    .f({haddr_pad[27],_al_u3128_o}),
    .q({open_n7917,\biu/cache_ctrl_logic/pa_temp [91]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2816|biu/cache_ctrl_logic/reg6_b90  (
    .a({open_n7918,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [23],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [90],\biu/paddress [90]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [24]}),
    .mi({open_n7929,\biu/paddress [90]}),
    .sr(rst_pad),
    .f({haddr_pad[26],_al_u3131_o}),
    .q({open_n7933,\biu/cache_ctrl_logic/pa_temp [90]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2817|biu/cache_ctrl_logic/reg6_b89  (
    .a({open_n7934,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [22],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [89],\biu/paddress [89]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [23]}),
    .mi({open_n7938,\biu/paddress [89]}),
    .sr(rst_pad),
    .f({haddr_pad[25],_al_u3134_o}),
    .q({open_n7953,\biu/cache_ctrl_logic/pa_temp [89]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2818|biu/cache_ctrl_logic/reg6_b88  (
    .a({open_n7954,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [21],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [88],\biu/paddress [88]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [22]}),
    .mi({open_n7958,\biu/paddress [88]}),
    .sr(rst_pad),
    .f({haddr_pad[24],_al_u3137_o}),
    .q({open_n7973,\biu/cache_ctrl_logic/pa_temp [88]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2819|biu/cache_ctrl_logic/reg6_b87  (
    .a({open_n7974,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [20],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [87],\biu/paddress [87]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [21]}),
    .mi({open_n7985,\biu/paddress [87]}),
    .sr(rst_pad),
    .f({haddr_pad[23],_al_u3140_o}),
    .q({open_n7989,\biu/cache_ctrl_logic/pa_temp [87]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2820|biu/cache_ctrl_logic/reg6_b86  (
    .a({open_n7990,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [19],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [86],\biu/paddress [86]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [20]}),
    .mi({open_n8001,\biu/paddress [86]}),
    .sr(rst_pad),
    .f({haddr_pad[22],_al_u3143_o}),
    .q({open_n8005,\biu/cache_ctrl_logic/pa_temp [86]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2821|biu/cache_ctrl_logic/reg6_b85  (
    .a({open_n8006,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [18],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [85],\biu/paddress [85]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [19]}),
    .mi({open_n8010,\biu/paddress [85]}),
    .sr(rst_pad),
    .f({haddr_pad[21],_al_u3146_o}),
    .q({open_n8025,\biu/cache_ctrl_logic/pa_temp [85]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2822|biu/cache_ctrl_logic/reg6_b84  (
    .a({open_n8026,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [17],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [84],\biu/paddress [84]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [18]}),
    .mi({open_n8030,\biu/paddress [84]}),
    .sr(rst_pad),
    .f({haddr_pad[20],_al_u3149_o}),
    .q({open_n8045,\biu/cache_ctrl_logic/pa_temp [84]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2823|biu/cache_ctrl_logic/reg6_b83  (
    .a({open_n8046,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [16],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [83],\biu/paddress [83]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [17]}),
    .mi({open_n8057,\biu/paddress [83]}),
    .sr(rst_pad),
    .f({haddr_pad[19],_al_u3153_o}),
    .q({open_n8061,\biu/cache_ctrl_logic/pa_temp [83]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2824|biu/cache_ctrl_logic/reg6_b82  (
    .a({open_n8062,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [15],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [82],\biu/paddress [82]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [16]}),
    .mi({open_n8073,\biu/paddress [82]}),
    .sr(rst_pad),
    .f({haddr_pad[18],_al_u3156_o}),
    .q({open_n8077,\biu/cache_ctrl_logic/pa_temp [82]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2825|biu/cache_ctrl_logic/reg6_b81  (
    .a({open_n8078,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [14],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [81],\biu/paddress [81]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [15]}),
    .mi({open_n8082,\biu/paddress [81]}),
    .sr(rst_pad),
    .f({haddr_pad[17],_al_u3159_o}),
    .q({open_n8097,\biu/cache_ctrl_logic/pa_temp [81]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2826|biu/cache_ctrl_logic/reg6_b80  (
    .a({open_n8098,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [13],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [80],\biu/paddress [80]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [14]}),
    .mi({open_n8102,\biu/paddress [80]}),
    .sr(rst_pad),
    .f({haddr_pad[16],_al_u3162_o}),
    .q({open_n8117,\biu/cache_ctrl_logic/pa_temp [80]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2827|biu/cache_ctrl_logic/reg6_b79  (
    .a({open_n8118,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [12],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [79],\biu/paddress [79]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [13]}),
    .mi({open_n8129,\biu/paddress [79]}),
    .sr(rst_pad),
    .f({haddr_pad[15],_al_u3165_o}),
    .q({open_n8133,\biu/cache_ctrl_logic/pa_temp [79]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000101000101),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2828|biu/cache_ctrl_logic/reg6_b78  (
    .a({open_n8134,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [11],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [78],\biu/paddress [78]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [12]}),
    .mi({open_n8145,\biu/paddress [78]}),
    .sr(rst_pad),
    .f({haddr_pad[14],_al_u3168_o}),
    .q({open_n8149,\biu/cache_ctrl_logic/pa_temp [78]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2829|biu/cache_ctrl_logic/reg6_b77  (
    .a({open_n8150,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [10],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [77],\biu/paddress [77]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [11]}),
    .mi({open_n8154,\biu/paddress [77]}),
    .sr(rst_pad),
    .f({haddr_pad[13],_al_u3171_o}),
    .q({open_n8169,\biu/cache_ctrl_logic/pa_temp [77]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000101000101),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000101000101),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2830|biu/cache_ctrl_logic/reg6_b76  (
    .a({open_n8170,_al_u2698_o}),
    .b({\biu/bus_unit/n49 [9],\biu/bus_unit/mmu/mux20_b0_sel_is_3_o }),
    .c({\biu/paddress [76],\biu/paddress [76]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u2705_o,\biu/bus_unit/mmu_hwdata [10]}),
    .mi({open_n8174,\biu/paddress [76]}),
    .sr(rst_pad),
    .f({haddr_pad[12],_al_u3174_o}),
    .q({open_n8189,\biu/cache_ctrl_logic/pa_temp [76]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2833|_al_u2705  (
    .c({\biu/bus_unit/statu [0],\biu/bus_unit/statu [0]}),
    .d({_al_u2704_o,_al_u2704_o}),
    .f({_al_u2833_o,_al_u2705_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~B*A)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~D*C*~B*A)"),
    //.LUTG1("(C*~B*D)"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2835|_al_u3223  (
    .a({open_n8214,\biu/cache_ctrl_logic/statu [1]}),
    .b(\biu/cache_ctrl_logic/statu [3:2]),
    .c(\biu/cache_ctrl_logic/statu [4:3]),
    .d({\biu/cache_ctrl_logic/statu [2],\biu/cache_ctrl_logic/statu [4]}),
    .f({_al_u2835_o,\biu/cache_ctrl_logic/n204_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2837|_al_u7160  (
    .b({open_n8241,_al_u2885_o}),
    .c({\biu/cache_ctrl_logic/statu [1],\biu/cache_ctrl_logic/statu [1]}),
    .d({\biu/cache_ctrl_logic/statu [0],_al_u7149_o}),
    .f({_al_u2837_o,_al_u7160_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*~A)"),
    //.LUT1("(C*~B*~D)"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"))
    \_al_u2838|_al_u2885  (
    .a({open_n8262,\biu/cache_ctrl_logic/statu [0]}),
    .b(\biu/cache_ctrl_logic/statu [3:2]),
    .c(\biu/cache_ctrl_logic/statu [4:3]),
    .d({\biu/cache_ctrl_logic/statu [2],\biu/cache_ctrl_logic/statu [4]}),
    .f({_al_u2838_o,_al_u2885_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*~D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~(~B*~D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000011000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000011000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2840|_al_u2842  (
    .b({open_n8285,1'b0}),
    .c({wb_valid,wb_valid}),
    .d(2'b00),
    .f({\cu_ru/m_s_status/n2 ,_al_u2842_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0101010000010000),
    .MODE("LOGIC"))
    \_al_u2845|_al_u6736  (
    .a({\cu_ru/m_s_status/n2 ,open_n8310}),
    .b({_al_u2844_o,_al_u2844_o}),
    .c({priv[1],\cu_ru/mtvec [2]}),
    .d({\cu_ru/mstatus [8],\cu_ru/trap_target_m }),
    .f({_al_u2845_o,_al_u6736_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(~D*C*B))"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(~A*~(~D*C*B))"),
    //.LUTG1("(~D*~C*~B*A)"),
    .INIT_LUTF0(16'b0101010100010101),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0101010100010101),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2848|_al_u3222  (
    .a({_al_u2847_o,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({\biu/cache_ctrl_logic/statu [2],_al_u2847_o}),
    .c({\biu/cache_ctrl_logic/statu [3],\biu/cache_ctrl_logic/statu [3]}),
    .d({\biu/cache_ctrl_logic/statu [4],\biu/cache_ctrl_logic/statu [4]}),
    .f({_al_u2848_o,_al_u3222_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~A*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0100010100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2850|cu_ru/m_s_status/reg1_b0  (
    .a({\cu_ru/m_s_status/n2 ,open_n8355}),
    .b({_al_u2844_o,open_n8356}),
    .c({priv[0],_al_u2850_o}),
    .clk(clk_pad),
    .d({\cu_ru/mstatus [8],_al_u2841_o}),
    .sr(rst_pad),
    .f({_al_u2850_o,open_n8370}),
    .q({open_n8374,priv[0]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u2853|_al_u2855  (
    .a({\exu/main_state [0],\exu/main_state [0]}),
    .b({\exu/main_state [1],\exu/main_state [1]}),
    .c({\exu/main_state [2],\exu/main_state [2]}),
    .d({\exu/main_state [3],\exu/main_state [3]}),
    .f({\exu/c_stb_lutinv ,_al_u2855_o}));
  // ../../RTL/CPU/EX/exu.v(290)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2856|exu/reg0_b7  (
    .b({\exu/shift_count [7],_al_u2856_o}),
    .c({\exu/n50 [7],op_count[7]}),
    .clk(clk_pad),
    .d({_al_u2855_o,\exu/n49 }),
    .sr(rst_pad),
    .f({_al_u2856_o,open_n8410}),
    .q({open_n8414,\exu/shift_count [7]}));  // ../../RTL/CPU/EX/exu.v(290)
  // ../../RTL/CPU/EX/exu.v(290)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2858|exu/reg0_b6  (
    .b({\exu/shift_count [6],_al_u2858_o}),
    .c({\exu/n50 [6],op_count[6]}),
    .clk(clk_pad),
    .d({_al_u2855_o,\exu/n49 }),
    .sr(rst_pad),
    .f({_al_u2858_o,open_n8430}),
    .q({open_n8434,\exu/shift_count [6]}));  // ../../RTL/CPU/EX/exu.v(290)
  // ../../RTL/CPU/EX/exu.v(290)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2860|exu/reg0_b5  (
    .b({\exu/shift_count [5],_al_u2860_o}),
    .c({\exu/n50 [5],op_count[5]}),
    .clk(clk_pad),
    .d({_al_u2855_o,\exu/n49 }),
    .sr(rst_pad),
    .f({_al_u2860_o,open_n8454}),
    .q({open_n8458,\exu/shift_count [5]}));  // ../../RTL/CPU/EX/exu.v(290)
  // ../../RTL/CPU/EX/exu.v(290)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2862|exu/reg0_b4  (
    .b({\exu/shift_count [4],_al_u2862_o}),
    .c({\exu/n50 [4],op_count[4]}),
    .clk(clk_pad),
    .d({_al_u2855_o,\exu/n49 }),
    .sr(rst_pad),
    .f({_al_u2862_o,open_n8478}),
    .q({open_n8482,\exu/shift_count [4]}));  // ../../RTL/CPU/EX/exu.v(290)
  // ../../RTL/CPU/EX/exu.v(290)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2864|exu/reg0_b3  (
    .b({\exu/shift_count [3],_al_u2864_o}),
    .c({\exu/n50 [3],op_count[3]}),
    .clk(clk_pad),
    .d({_al_u2855_o,\exu/n49 }),
    .sr(rst_pad),
    .f({_al_u2864_o,open_n8498}),
    .q({open_n8502,\exu/shift_count [3]}));  // ../../RTL/CPU/EX/exu.v(290)
  // ../../RTL/CPU/EX/exu.v(290)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2866|exu/reg0_b2  (
    .b({\exu/shift_count [2],_al_u2866_o}),
    .c({\exu/n50 [2],op_count[2]}),
    .clk(clk_pad),
    .d({_al_u2855_o,\exu/n49 }),
    .sr(rst_pad),
    .f({_al_u2866_o,open_n8518}),
    .q({open_n8522,\exu/shift_count [2]}));  // ../../RTL/CPU/EX/exu.v(290)
  // ../../RTL/CPU/EX/exu.v(290)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2868|exu/reg0_b1  (
    .b({\exu/shift_count [1],_al_u2868_o}),
    .c({\exu/n50 [1],op_count[1]}),
    .clk(clk_pad),
    .d({_al_u2855_o,\exu/n49 }),
    .sr(rst_pad),
    .f({_al_u2868_o,open_n8542}),
    .q({open_n8546,\exu/shift_count [1]}));  // ../../RTL/CPU/EX/exu.v(290)
  // ../../RTL/CPU/EX/exu.v(290)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2870|exu/reg0_b0  (
    .b({\exu/shift_count [0],_al_u2870_o}),
    .c({\exu/n50 [0],op_count[0]}),
    .clk(clk_pad),
    .d({_al_u2855_o,\exu/n49 }),
    .sr(rst_pad),
    .f({_al_u2870_o,open_n8566}),
    .q({open_n8570,\exu/shift_count [0]}));  // ../../RTL/CPU/EX/exu.v(290)
  // ../../RTL/CPU/BIU/mmu.v(154)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2872|biu/bus_unit/mmu/reg4_b3  (
    .a({open_n8571,_al_u7206_o}),
    .b({open_n8572,_al_u7208_o}),
    .c({rst_pad,_al_u2964_o}),
    .clk(clk_pad),
    .d({_al_u2697_o,hresp_pad}),
    .sr(\biu/bus_unit/mmu/mux18_b3_sel_is_2_o ),
    .f({\biu/bus_unit/mmu/mux18_b3_sel_is_2_o ,open_n8586}),
    .q({open_n8590,\biu/bus_unit/mmu/statu [3]}));  // ../../RTL/CPU/BIU/mmu.v(154)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u2873|_al_u2875  (
    .a({open_n8591,_al_u2873_o}),
    .b({\biu/bus_unit/addr_counter [7],_al_u2874_o}),
    .c({\biu/bus_unit/addr_counter [8],\biu/bus_unit/addr_counter [0]}),
    .d({\biu/bus_unit/addr_counter [6],\biu/bus_unit/addr_counter [1]}),
    .f({_al_u2873_o,\biu/bus_unit/n15_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u2874|_al_u2901  (
    .a({\biu/bus_unit/addr_counter [2],open_n8612}),
    .b({\biu/bus_unit/addr_counter [3],\biu/bus_unit/addr_counter [3]}),
    .c({\biu/bus_unit/addr_counter [4],\biu/bus_unit/last_addr [3]}),
    .d({\biu/bus_unit/addr_counter [5],_al_u2890_o}),
    .f({_al_u2874_o,_al_u2901_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2886|_al_u2913  (
    .c({\biu/cache_ctrl_logic/statu [1],\biu/cache_ctrl_logic/statu [1]}),
    .d({_al_u2885_o,_al_u2885_o}),
    .f({_al_u2886_o,\biu/bus_unit/mmu/n19_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*C*~B*A)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"))
    \_al_u2887|_al_u3947  (
    .a({_al_u2837_o,open_n8661}),
    .b({\biu/cache_ctrl_logic/statu [2],open_n8662}),
    .c({\biu/cache_ctrl_logic/statu [3],_al_u3944_o}),
    .d({\biu/cache_ctrl_logic/statu [4],_al_u2837_o}),
    .f({\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ,_al_u3947_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2890|_al_u2889  (
    .b({open_n8685,\biu/bus_unit/statu [1]}),
    .c({_al_u2889_o,\biu/bus_unit/statu [3]}),
    .d({_al_u2703_o,\biu/bus_unit/statu [0]}),
    .f({_al_u2890_o,_al_u2889_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"))
    \_al_u2891|_al_u2892  (
    .b({\biu/bus_unit/addr_counter [8],_al_u2891_o}),
    .c({\biu/bus_unit/last_addr [8],addr_ex[8]}),
    .d({_al_u2890_o,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .f({_al_u2891_o,\biu/l1d_addr [8]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2895|_al_u2896  (
    .b({\biu/bus_unit/addr_counter [6],_al_u2895_o}),
    .c({\biu/bus_unit/last_addr [6],addr_ex[6]}),
    .d({_al_u2890_o,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .f({_al_u2895_o,\biu/l1d_addr [6]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"))
    \_al_u2897|_al_u2898  (
    .b({\biu/bus_unit/addr_counter [5],_al_u2897_o}),
    .c({\biu/bus_unit/last_addr [5],addr_ex[5]}),
    .d({_al_u2890_o,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .f({_al_u2897_o,\biu/l1d_addr [5]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"))
    \_al_u2899|_al_u2900  (
    .b({\biu/bus_unit/addr_counter [4],_al_u2899_o}),
    .c({\biu/bus_unit/last_addr [4],addr_ex[4]}),
    .d({_al_u2890_o,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .f({_al_u2899_o,\biu/l1d_addr [4]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"))
    \_al_u2903|_al_u2904  (
    .b({\biu/bus_unit/addr_counter [2],_al_u2903_o}),
    .c({\biu/bus_unit/last_addr [2],addr_ex[2]}),
    .d({_al_u2890_o,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .f({_al_u2903_o,\biu/l1d_addr [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"))
    \_al_u2905|_al_u2906  (
    .b({\biu/bus_unit/addr_counter [1],_al_u2905_o}),
    .c({\biu/bus_unit/last_addr [1],addr_ex[1]}),
    .d({_al_u2890_o,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .f({_al_u2905_o,\biu/l1d_addr [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2907|_al_u2908  (
    .b({\biu/bus_unit/addr_counter [0],_al_u2907_o}),
    .c({\biu/bus_unit/last_addr [0],addr_ex[0]}),
    .d({_al_u2890_o,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .f({_al_u2907_o,\biu/l1d_addr [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2910|_al_u2909  (
    .b({open_n8870,\exu/main_state [1]}),
    .c({\exu/main_state [2],\exu/main_state [3]}),
    .d({_al_u2909_o,\exu/main_state [0]}),
    .f({_al_u2910_o,_al_u2909_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2916|_al_u2699  (
    .b({\biu/bus_unit/mmu/i [0],open_n8893}),
    .c({\biu/bus_unit/mmu/i [1],rst_pad}),
    .d({_al_u2915_o,_al_u2698_o}),
    .f({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/n58 }));
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0000001100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2929|ins_fetch/reg1_b4  (
    .a({ins_read[4],open_n8918}),
    .b({ins_read[36],ins_read[36]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[4]}),
    .sr(rst_pad),
    .f({_al_u2929_o,open_n8931}),
    .q({open_n8935,\ins_fetch/ins_hold [4]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0000001100000101),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0000001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2931|ins_fetch/reg1_b3  (
    .a({ins_read[3],open_n8936}),
    .b({ins_read[35],ins_read[35]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[3]}),
    .sr(rst_pad),
    .f({_al_u2931_o,open_n8953}),
    .q({open_n8957,\ins_fetch/ins_hold [3]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~(~D*~C)*~(~B*~A))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1110111011100000),
    .MODE("LOGIC"))
    \_al_u2933|_al_u2932  (
    .a({_al_u2929_o,open_n8958}),
    .b({_al_u2930_o,open_n8959}),
    .c({_al_u2931_o,\ins_fetch/ins_hold [3]}),
    .d({_al_u2932_o,1'b0}),
    .f({_al_u2933_o,_al_u2932_o}));
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0000001100000101),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2934|ins_dec/reg10_b0  (
    .a({ins_read[0],open_n8980}),
    .b({ins_read[32],_al_u2934_o}),
    .c({1'b0,_al_u2935_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins_pc[2],id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u2934_o,open_n8997}),
    .q({open_n9001,ex_exc_code[0]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2935|_al_u2937  (
    .c({\ins_fetch/ins_hold [0],\ins_fetch/ins_hold [1]}),
    .d(2'b00),
    .f({_al_u2935_o,_al_u2937_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0000001100000101),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0000001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2936|ins_fetch/reg1_b1  (
    .a({ins_read[1],open_n9030}),
    .b({ins_read[33],ins_read[33]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[1]}),
    .sr(rst_pad),
    .f({_al_u2936_o,open_n9047}),
    .q({open_n9051,\ins_fetch/ins_hold [1]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2938|ins_dec/reg10_b1  (
    .a({_al_u2934_o,open_n9052}),
    .b({_al_u2935_o,_al_u2936_o}),
    .c({_al_u2936_o,_al_u2937_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u2937_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u2938_o,open_n9065}),
    .q({open_n9069,ex_exc_code[1]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2939|ins_fetch/reg1_b2  (
    .b({1'b0,ins_read[34]}),
    .c({\ins_fetch/ins_hold [2],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({\ins_fetch/ins_shift [2],ins_read[2]}),
    .sr(rst_pad),
    .f({_al_u2939_o,\ins_fetch/ins_shift [2]}),
    .q({open_n9091,\ins_fetch/ins_hold [2]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0000001100000101),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0000001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2940|ins_fetch/reg1_b6  (
    .a({ins_read[6],open_n9092}),
    .b({ins_read[38],ins_read[38]}),
    .c({1'b0,id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({id_ins_pc[2],ins_read[6]}),
    .sr(rst_pad),
    .f({_al_u2940_o,open_n9109}),
    .q({open_n9113,\ins_fetch/ins_hold [6]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2943|ins_fetch/reg1_b5  (
    .b({open_n9116,ins_read[37]}),
    .c({\ins_fetch/ins_hold [5],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({1'b0,ins_read[5]}),
    .sr(rst_pad),
    .f({_al_u2943_o,open_n9133}),
    .q({open_n9137,\ins_fetch/ins_hold [5]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~D*~C*~(~B*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000101),
    .INIT_LUT1(16'b0000000000001110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2944|ins_dec/reg11_b2  (
    .a({_al_u2940_o,ins_read[5]}),
    .b({_al_u2941_o,ins_read[37]}),
    .c({_al_u2942_o,1'b0}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u2943_o,id_ins_pc[2]}),
    .mi({open_n9148,id_ins_pc[2]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u2944_o,_al_u2942_o}),
    .q({open_n9152,ex_ins_pc[2]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(~(~D*~C)*~(~B*~A))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(~(~D*~C)*~(~B*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b1110111011100000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1110111011100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2946|ins_dec/reg10_b6  (
    .a({_al_u2940_o,open_n9153}),
    .b({_al_u2941_o,_al_u2940_o}),
    .c({_al_u2942_o,_al_u2941_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u2943_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u2946_o,open_n9170}),
    .q({open_n9174,ex_exc_code[6]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~D*~C*~(~B*~A))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~D*~C*~(~B*~A))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000001110),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2948|_al_u2930  (
    .a({_al_u2929_o,open_n9175}),
    .b({_al_u2930_o,open_n9176}),
    .c({_al_u2931_o,\ins_fetch/ins_hold [4]}),
    .d({_al_u2932_o,1'b0}),
    .f({_al_u2948_o,_al_u2930_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(D*~C*B*A)"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2952|_al_u3403  (
    .a({_al_u2703_o,_al_u2703_o}),
    .b({\biu/bus_unit/statu [0],\biu/bus_unit/statu [0]}),
    .c({\biu/bus_unit/statu [1],\biu/bus_unit/statu [1]}),
    .d({\biu/bus_unit/statu [3],\biu/bus_unit/statu [3]}),
    .f({_al_u2952_o,_al_u3403_o}));
  // ../../RTL/CPU/BIU/bus_unit.v(177)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("~(~A*~(D*~(~C*~B)))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("~(~A*~(D*~(~C*~B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111010101010),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111111010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2953|biu/bus_unit/reg0_b4  (
    .a({\biu/bus_unit/n15_lutinv ,open_n9225}),
    .b({htrans_pad[0],open_n9226}),
    .c({_al_u2952_o,\biu/bus_unit/n39 [4]}),
    .ce(\biu/bus_unit/n39[0]_en ),
    .clk(clk_pad),
    .d({hready_pad,\biu/bus_unit/n15_lutinv }),
    .sr(\biu/bus_unit/n37 ),
    .f({\biu/bus_unit/n39[0]_en ,open_n9243}),
    .q({open_n9247,\biu/bus_unit/addr_counter [4]}));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~C*~B*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"))
    \_al_u2956|_al_u3404  (
    .b({\biu/bus_unit/statu [0],\biu/bus_unit/statu [0]}),
    .c({\biu/bus_unit/statu [1],\biu/bus_unit/statu [1]}),
    .d({_al_u2955_o,_al_u2955_o}),
    .f({_al_u2956_o,_al_u3404_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(~B*~(D*~C)))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0111010101110111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u2957|_al_u3220  (
    .a({open_n9270,_al_u2706_o}),
    .b({open_n9271,ex_size[0]}),
    .c({_al_u2956_o,ex_size[1]}),
    .d({_al_u2706_o,ex_size[2]}),
    .f({_al_u2957_o,hsize_pad[0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2959|_al_u2958  (
    .b({open_n9294,\biu/bus_unit/statu [0]}),
    .c({_al_u2958_o,\biu/bus_unit/statu [1]}),
    .d({_al_u2957_o,_al_u2703_o}),
    .f({\biu/bus_unit/mux15_b4_sel_is_2_o ,_al_u2958_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~D*~C*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1010101010100010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u2960|_al_u2954  (
    .a({open_n9315,_al_u2705_o}),
    .b({\biu/bus_unit/mux15_b4_sel_is_2_o ,\biu/bus_unit/mmu/statu [0]}),
    .c({htrans_pad[0],\biu/bus_unit/mmu/statu [1]}),
    .d({_al_u2954_o,\biu/bus_unit/mmu/statu [3]}),
    .f({htrans_pad[1],_al_u2954_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~C*~D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"))
    \_al_u2961|_al_u3417  (
    .c({_al_u2952_o,\biu/bus_unit/mux15_b4_sel_is_2_o }),
    .d({htrans_pad[0],\biu/bus_unit/n37 }),
    .f({hburst_pad[0],\biu/bus_unit/mux17_b4_sel_is_2_o }));
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(D*~C*~B*~A)"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100000000),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2962|cu_ru/csr_satp/reg1_b2  (
    .a({satp[60],\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({satp[61],\cu_ru/trap_target_m }),
    .c({satp[62],\cu_ru/mepc [62]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[63],data_csr[62]}),
    .mi({open_n9363,data_csr[62]}),
    .sr(rst_pad),
    .f({\biu/bus_unit/mmu/n31_lutinv ,_al_u6580_o}),
    .q({open_n9378,satp[62]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2965|_al_u5803  (
    .b({open_n9381,_al_u2705_o}),
    .c({hready_pad,\biu/bus_unit/mmu_hwdata [32]}),
    .d({_al_u2964_o,_al_u5802_o}),
    .f({\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ,hwdata_pad[32]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0011001100001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2966|biu/cache_ctrl_logic/reg7_b9  (
    .b({hrdata_pad[9],open_n9408}),
    .c({\biu/bus_unit/mmu_hwdata [9],hrdata_pad[9]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ,_al_u2705_o}),
    .sr(rst_pad),
    .f({_al_u2966_o,uncache_data[9]}),
    .q({open_n9424,\biu/cache_ctrl_logic/pte_temp [9]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(~D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0000000011001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2974|biu/bus_unit/mmu/reg3_b6  (
    .b({\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ,open_n9427}),
    .c({\biu/bus_unit/mmu_hwdata [6],_al_u2975_o}),
    .clk(clk_pad),
    .d({_al_u2963_o,_al_u2974_o}),
    .sr(rst_pad),
    .f({_al_u2974_o,open_n9441}),
    .q({open_n9445,\biu/bus_unit/mmu_hwdata [6]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2975|biu/cache_ctrl_logic/reg7_b6  (
    .b({_al_u2915_o,open_n9448}),
    .c({hrdata_pad[6],hrdata_pad[6]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ,_al_u2705_o}),
    .sr(rst_pad),
    .f({_al_u2975_o,uncache_data[6]}),
    .q({open_n9468,\biu/cache_ctrl_logic/pte_temp [6]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3033|biu/bus_unit/mmu/reg2_b13  (
    .c({\biu/bus_unit/mmu/n31_lutinv ,_al_u3171_o}),
    .clk(clk_pad),
    .d({_al_u2914_o,_al_u3170_o}),
    .sr(rst_pad),
    .f({_al_u3033_o,open_n9486}),
    .q({open_n9490,\biu/paddress [77]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000001111001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3034|biu/bus_unit/mmu/reg2_b58  (
    .b({_al_u2698_o,open_n9493}),
    .c({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/paddress [122]}),
    .clk(clk_pad),
    .d({_al_u3033_o,_al_u3034_o}),
    .sr(rst_pad),
    .f({_al_u3034_o,open_n9507}),
    .q({open_n9511,\biu/paddress [122]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3043|cu_ru/csr_satp/reg0_b43  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [119],\cu_ru/mepc [43]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[43],data_csr[43]}),
    .mi({open_n9522,data_csr[43]}),
    .sr(rst_pad),
    .f({_al_u3043_o,_al_u6622_o}),
    .q({open_n9526,satp[43]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3046|cu_ru/csr_satp/reg0_b42  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [118],\cu_ru/mepc [42]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[42],data_csr[42]}),
    .mi({open_n9530,data_csr[42]}),
    .sr(rst_pad),
    .f({_al_u3046_o,_al_u6624_o}),
    .q({open_n9545,satp[42]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3049|cu_ru/csr_satp/reg0_b41  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [117],\cu_ru/mepc [41]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[41],data_csr[41]}),
    .mi({open_n9549,data_csr[41]}),
    .sr(rst_pad),
    .f({_al_u3049_o,_al_u6626_o}),
    .q({open_n9564,satp[41]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3052|cu_ru/csr_satp/reg0_b40  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [116],\cu_ru/mepc [40]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[40],data_csr[40]}),
    .mi({open_n9575,data_csr[40]}),
    .sr(rst_pad),
    .f({_al_u3052_o,_al_u6628_o}),
    .q({open_n9579,satp[40]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3055|cu_ru/csr_satp/reg0_b39  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [115],\cu_ru/mepc [39]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[39],data_csr[39]}),
    .mi({open_n9590,data_csr[39]}),
    .sr(rst_pad),
    .f({_al_u3055_o,_al_u6632_o}),
    .q({open_n9594,satp[39]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3058|cu_ru/csr_satp/reg0_b38  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [114],\cu_ru/mepc [38]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[38],data_csr[38]}),
    .mi({open_n9598,data_csr[38]}),
    .sr(rst_pad),
    .f({_al_u3058_o,_al_u6634_o}),
    .q({open_n9613,satp[38]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3061|cu_ru/csr_satp/reg0_b37  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [113],\cu_ru/mepc [37]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[37],data_csr[37]}),
    .mi({open_n9617,data_csr[37]}),
    .sr(rst_pad),
    .f({_al_u3061_o,_al_u6636_o}),
    .q({open_n9632,satp[37]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3064|cu_ru/csr_satp/reg0_b36  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [112],\cu_ru/mepc [36]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[36],data_csr[36]}),
    .mi({open_n9643,data_csr[36]}),
    .sr(rst_pad),
    .f({_al_u3064_o,_al_u6638_o}),
    .q({open_n9647,satp[36]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3067|cu_ru/csr_satp/reg0_b35  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [111],\cu_ru/mepc [35]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[35],data_csr[35]}),
    .mi({open_n9658,data_csr[35]}),
    .sr(rst_pad),
    .f({_al_u3067_o,_al_u6640_o}),
    .q({open_n9662,satp[35]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3070|cu_ru/csr_satp/reg0_b34  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [110],\cu_ru/mepc [34]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[34],data_csr[34]}),
    .mi({open_n9666,data_csr[34]}),
    .sr(rst_pad),
    .f({_al_u3070_o,_al_u6642_o}),
    .q({open_n9681,satp[34]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3073|cu_ru/csr_satp/reg0_b33  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [109],\cu_ru/mepc [33]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[33],data_csr[33]}),
    .mi({open_n9685,data_csr[33]}),
    .sr(rst_pad),
    .f({_al_u3073_o,_al_u6644_o}),
    .q({open_n9700,satp[33]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3076|cu_ru/csr_satp/reg0_b32  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [108],\cu_ru/mepc [32]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[32],data_csr[32]}),
    .mi({open_n9711,data_csr[32]}),
    .sr(rst_pad),
    .f({_al_u3076_o,_al_u6646_o}),
    .q({open_n9715,satp[32]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3079|cu_ru/csr_satp/reg0_b31  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [107],\cu_ru/mepc [31]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[31],data_csr[31]}),
    .mi({open_n9726,data_csr[31]}),
    .sr(rst_pad),
    .f({_al_u3079_o,_al_u6648_o}),
    .q({open_n9730,satp[31]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3082|cu_ru/csr_satp/reg0_b30  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [106],\cu_ru/mepc [30]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[30],data_csr[30]}),
    .mi({open_n9734,data_csr[30]}),
    .sr(rst_pad),
    .f({_al_u3082_o,_al_u6650_o}),
    .q({open_n9749,satp[30]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3085|cu_ru/csr_satp/reg0_b29  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [105],\cu_ru/mepc [29]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[29],data_csr[29]}),
    .mi({open_n9753,data_csr[29]}),
    .sr(rst_pad),
    .f({_al_u3085_o,_al_u6654_o}),
    .q({open_n9768,satp[29]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3088|cu_ru/csr_satp/reg0_b28  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [104],\cu_ru/mepc [28]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[28],data_csr[28]}),
    .mi({open_n9779,data_csr[28]}),
    .sr(rst_pad),
    .f({_al_u3088_o,_al_u6656_o}),
    .q({open_n9783,satp[28]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3091|cu_ru/csr_satp/reg0_b27  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [103],\cu_ru/mepc [27]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[27],data_csr[27]}),
    .mi({open_n9794,data_csr[27]}),
    .sr(rst_pad),
    .f({_al_u3091_o,_al_u6658_o}),
    .q({open_n9798,satp[27]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3094|cu_ru/csr_satp/reg0_b26  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [102],\cu_ru/mepc [26]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[26],data_csr[26]}),
    .mi({open_n9802,data_csr[26]}),
    .sr(rst_pad),
    .f({_al_u3094_o,_al_u6660_o}),
    .q({open_n9817,satp[26]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3097|cu_ru/csr_satp/reg0_b25  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [101],\cu_ru/mepc [25]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[25],data_csr[25]}),
    .mi({open_n9821,data_csr[25]}),
    .sr(rst_pad),
    .f({_al_u3097_o,_al_u6662_o}),
    .q({open_n9836,satp[25]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3100|cu_ru/csr_satp/reg0_b24  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [100],\cu_ru/mepc [24]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[24],data_csr[24]}),
    .mi({open_n9847,data_csr[24]}),
    .sr(rst_pad),
    .f({_al_u3100_o,_al_u6664_o}),
    .q({open_n9851,satp[24]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3103|cu_ru/csr_satp/reg0_b23  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [99],\cu_ru/mepc [23]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[23],data_csr[23]}),
    .mi({open_n9862,data_csr[23]}),
    .sr(rst_pad),
    .f({_al_u3103_o,_al_u6666_o}),
    .q({open_n9866,satp[23]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3106|cu_ru/csr_satp/reg0_b22  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [98],\cu_ru/mepc [22]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[22],data_csr[22]}),
    .mi({open_n9870,data_csr[22]}),
    .sr(rst_pad),
    .f({_al_u3106_o,_al_u6668_o}),
    .q({open_n9885,satp[22]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3109|cu_ru/csr_satp/reg0_b21  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [97],\cu_ru/mepc [21]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[21],data_csr[21]}),
    .mi({open_n9889,data_csr[21]}),
    .sr(rst_pad),
    .f({_al_u3109_o,_al_u6670_o}),
    .q({open_n9904,satp[21]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3112|cu_ru/csr_satp/reg0_b20  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [96],\cu_ru/mepc [20]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[20],data_csr[20]}),
    .mi({open_n9915,data_csr[20]}),
    .sr(rst_pad),
    .f({_al_u3112_o,_al_u6672_o}),
    .q({open_n9919,satp[20]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3115|cu_ru/csr_satp/reg0_b19  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [95],\cu_ru/mepc [19]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[19],data_csr[19]}),
    .mi({open_n9930,data_csr[19]}),
    .sr(rst_pad),
    .f({_al_u3115_o,_al_u6676_o}),
    .q({open_n9934,satp[19]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3118|cu_ru/csr_satp/reg0_b18  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [94],\cu_ru/mepc [18]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[18],data_csr[18]}),
    .mi({open_n9938,data_csr[18]}),
    .sr(rst_pad),
    .f({_al_u3118_o,_al_u6678_o}),
    .q({open_n9953,satp[18]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3121|cu_ru/csr_satp/reg0_b17  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [93],\cu_ru/mepc [17]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[17],data_csr[17]}),
    .mi({open_n9957,data_csr[17]}),
    .sr(rst_pad),
    .f({_al_u3121_o,_al_u6680_o}),
    .q({open_n9972,satp[17]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3124|cu_ru/csr_satp/reg0_b16  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [92],\cu_ru/mepc [16]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[16],data_csr[16]}),
    .mi({open_n9976,data_csr[16]}),
    .sr(rst_pad),
    .f({_al_u3124_o,_al_u6682_o}),
    .q({open_n9991,satp[16]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3127|cu_ru/csr_satp/reg0_b15  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [91],\cu_ru/mepc [15]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[15],data_csr[15]}),
    .mi({open_n10002,data_csr[15]}),
    .sr(rst_pad),
    .f({_al_u3127_o,_al_u6684_o}),
    .q({open_n10006,satp[15]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3130|cu_ru/csr_satp/reg0_b14  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [90],\cu_ru/mepc [14]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[14],data_csr[14]}),
    .mi({open_n10010,data_csr[14]}),
    .sr(rst_pad),
    .f({_al_u3130_o,_al_u6686_o}),
    .q({open_n10025,satp[14]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3133|cu_ru/csr_satp/reg0_b13  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [89],\cu_ru/mepc [13]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[13],data_csr[13]}),
    .mi({open_n10036,data_csr[13]}),
    .sr(rst_pad),
    .f({_al_u3133_o,_al_u6688_o}),
    .q({open_n10040,satp[13]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3136|cu_ru/csr_satp/reg0_b12  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [88],\cu_ru/mepc [12]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[12],data_csr[12]}),
    .mi({open_n10044,data_csr[12]}),
    .sr(rst_pad),
    .f({_al_u3136_o,_al_u6690_o}),
    .q({open_n10059,satp[12]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3139|cu_ru/csr_satp/reg0_b11  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [87],\cu_ru/mepc [11]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[11],data_csr[11]}),
    .mi({open_n10063,data_csr[11]}),
    .sr(rst_pad),
    .f({_al_u3139_o,_al_u6692_o}),
    .q({open_n10078,satp[11]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3142|cu_ru/csr_satp/reg0_b10  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [86],\cu_ru/mepc [10]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[10],data_csr[10]}),
    .mi({open_n10089,data_csr[10]}),
    .sr(rst_pad),
    .f({_al_u3142_o,_al_u6694_o}),
    .q({open_n10093,satp[10]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3145|cu_ru/csr_satp/reg0_b9  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [85],\cu_ru/mepc [9]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[9],data_csr[9]}),
    .mi({open_n10097,data_csr[9]}),
    .sr(rst_pad),
    .f({_al_u3145_o,_al_u6570_o}),
    .q({open_n10112,satp[9]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3148|cu_ru/csr_satp/reg0_b8  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [84],\cu_ru/mepc [8]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[8],data_csr[8]}),
    .mi({open_n10123,data_csr[8]}),
    .sr(rst_pad),
    .f({_al_u3148_o,_al_u6572_o}),
    .q({open_n10127,satp[8]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3152|cu_ru/csr_satp/reg0_b7  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [83],\cu_ru/mepc [7]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[7],data_csr[7]}),
    .mi({open_n10138,data_csr[7]}),
    .sr(rst_pad),
    .f({_al_u3152_o,_al_u6574_o}),
    .q({open_n10142,satp[7]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3155|cu_ru/csr_satp/reg0_b6  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [82],\cu_ru/mepc [6]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[6],data_csr[6]}),
    .mi({open_n10153,data_csr[6]}),
    .sr(rst_pad),
    .f({_al_u3155_o,_al_u6576_o}),
    .q({open_n10157,satp[6]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3158|cu_ru/csr_satp/reg0_b5  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [81],\cu_ru/mepc [5]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[5],data_csr[5]}),
    .mi({open_n10161,data_csr[5]}),
    .sr(rst_pad),
    .f({_al_u3158_o,_al_u6586_o}),
    .q({open_n10176,satp[5]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3161|cu_ru/csr_satp/reg0_b4  (
    .a({_al_u3033_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2698_o,\cu_ru/trap_target_m }),
    .c({\biu/paddress [80],\cu_ru/mepc [4]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[4],data_csr[4]}),
    .mi({open_n10187,data_csr[4]}),
    .sr(rst_pad),
    .f({_al_u3161_o,_al_u6608_o}),
    .q({open_n10191,satp[4]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3164|cu_ru/csr_satp/reg0_b3  (
    .a({_al_u3033_o,open_n10192}),
    .b({_al_u2698_o,\cu_ru/scause [3]}),
    .c({\biu/paddress [79],data_csr[3]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[3],\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .mi({open_n10196,data_csr[3]}),
    .sr(rst_pad),
    .f({_al_u3164_o,_al_u6729_o}),
    .q({open_n10211,satp[3]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3167|cu_ru/csr_satp/reg0_b2  (
    .a({_al_u3033_o,open_n10212}),
    .b({_al_u2698_o,\cu_ru/mcause [2]}),
    .c({\biu/paddress [78],data_csr[2]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[2],\cu_ru/m_s_cause/mux4_b0_sel_is_2_o }),
    .mi({open_n10223,data_csr[2]}),
    .sr(rst_pad),
    .f({_al_u3167_o,_al_u6700_o}),
    .q({open_n10227,satp[2]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3170|cu_ru/csr_satp/reg0_b1  (
    .a({_al_u3033_o,open_n10228}),
    .b({_al_u2698_o,\cu_ru/scause [1]}),
    .c({\biu/paddress [77],data_csr[1]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({satp[1],\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .mi({open_n10239,data_csr[1]}),
    .sr(rst_pad),
    .f({_al_u3170_o,_al_u7337_o}),
    .q({open_n10243,satp[1]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3173|biu/bus_unit/mmu/reg2_b15  (
    .a({_al_u3033_o,open_n10244}),
    .b({_al_u2698_o,open_n10245}),
    .c({\biu/paddress [76],_al_u3165_o}),
    .clk(clk_pad),
    .d({satp[0],_al_u3164_o}),
    .sr(rst_pad),
    .f({_al_u3173_o,open_n10263}),
    .q({open_n10267,\biu/paddress [79]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1101110101010000),
    .MODE("LOGIC"))
    \_al_u3179|_al_u3178  (
    .a({\exu/lsu/n0_lutinv ,open_n10268}),
    .b({addr_ex[2],open_n10269}),
    .c({ex_size[2],addr_ex[1]}),
    .d({ex_size[3],addr_ex[0]}),
    .f({_al_u3179_o,\exu/lsu/n0_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~A*~(D*C*B))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010101010101),
    .MODE("LOGIC"))
    \_al_u3181|_al_u3180  (
    .a({_al_u3179_o,open_n10290}),
    .b({\exu/lsu/n8_lutinv ,open_n10291}),
    .c(addr_ex[2:1]),
    .d({ex_size[1],addr_ex[0]}),
    .f({_al_u3181_o,\exu/lsu/n8_lutinv }));
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3185|exu/csr_write_reg  (
    .a({_al_u3183_o,open_n10312}),
    .b({_al_u3184_o,open_n10313}),
    .c({csr_index[1],wb_valid}),
    .clk(clk_pad),
    .d({csr_index[2],wb_csr_write}),
    .mi({open_n10318,ex_csr_write}),
    .sr(rst_pad),
    .f({_al_u3185_o,_al_u3184_o}),
    .q({open_n10333,wb_csr_write}));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3187|cu_ru/csr_satp/reg0_b0  (
    .a({_al_u3186_o,open_n10334}),
    .b({csr_index[6],open_n10335}),
    .c({csr_index[7],_al_u3187_o}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({csr_index[8],_al_u3185_o}),
    .mi({open_n10339,data_csr[0]}),
    .sr(rst_pad),
    .f({_al_u3187_o,\cu_ru/csr_satp/n0 }),
    .q({open_n10354,satp[0]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~D)"),
    //.LUT1("(D*~C*B*A)"),
    .INIT_LUT0(16'b0000000011000000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"))
    \_al_u3191|_al_u5992  (
    .a({_al_u3183_o,open_n10355}),
    .b({_al_u3184_o,_al_u3190_o}),
    .c({csr_index[1],_al_u3184_o}),
    .d({csr_index[2],_al_u5157_o}),
    .f({_al_u3191_o,_al_u5992_o}));
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3195|exu/reg6_b8  (
    .a({open_n10376,_al_u3189_o}),
    .b({open_n10377,csr_index[6]}),
    .c({_al_u3194_o,csr_index[7]}),
    .clk(clk_pad),
    .d({_al_u3189_o,csr_index[8]}),
    .mi({open_n10382,ex_csr_index[8]}),
    .sr(rst_pad),
    .f({_al_u3195_o,_al_u3190_o}),
    .q({open_n10397,csr_index[8]}));  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*~C*B*A)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3201|_al_u3253  (
    .a({_al_u3184_o,open_n10398}),
    .b({_al_u3200_o,open_n10399}),
    .c({csr_index[1],_al_u3252_o}),
    .d({csr_index[2],_al_u3185_o}),
    .f({_al_u3201_o,_al_u3253_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3204|_al_u5159  (
    .b({csr_index[1],open_n10426}),
    .c({csr_index[2],_al_u3204_o}),
    .d({_al_u3200_o,_al_u5158_o}),
    .f({_al_u3204_o,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3208|_al_u9153  (
    .c({\exu/main_state [2],\exu/main_state [3]}),
    .d({_al_u2909_o,\exu/main_state [2]}),
    .f({\exu/c_fence_lutinv ,_al_u9153_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3209|_al_u2847  (
    .c({\biu/cache_ctrl_logic/statu [1],\biu/cache_ctrl_logic/statu [1]}),
    .d({\biu/cache_ctrl_logic/statu [0],\biu/cache_ctrl_logic/statu [0]}),
    .f({_al_u3209_o,_al_u2847_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~D*~C*~B*A)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"))
    \_al_u3210|_al_u3945  (
    .a({_al_u3209_o,open_n10503}),
    .b({\biu/cache_ctrl_logic/statu [2],open_n10504}),
    .c({\biu/cache_ctrl_logic/statu [3],_al_u3944_o}),
    .d({\biu/cache_ctrl_logic/statu [4],_al_u3209_o}),
    .f({\biu/cache_ctrl_logic/n55_lutinv ,_al_u3945_o}));
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3212|ins_dec/reg10_b5  (
    .a({_al_u2940_o,open_n10525}),
    .b({_al_u2941_o,_al_u2942_o}),
    .c({_al_u2942_o,_al_u2943_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u2943_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3212_o,open_n10538}),
    .q({open_n10542,ex_exc_code[5]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3213|ins_dec/reg10_b2  (
    .a({_al_u2933_o,open_n10543}),
    .b({_al_u2938_o,open_n10544}),
    .c({_al_u2939_o,_al_u2939_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3212_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3213_o,open_n10557}),
    .q({open_n10561,ex_exc_code[2]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3214|ins_dec/amo_reg  (
    .a({_al_u2938_o,_al_u2938_o}),
    .b({_al_u2939_o,_al_u2939_o}),
    .c({_al_u2948_o,_al_u2944_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3212_o,_al_u2948_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3214_o,\ins_dec/op_amo }),
    .q({open_n10581,amo}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3218|ins_dec/reg10_b13  (
    .c({_al_u3217_o,_al_u3217_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3216_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/n35_lutinv ,open_n10598}),
    .q({open_n10602,ex_exc_code[13]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3224|_al_u4403  (
    .c({\biu/cache_ctrl_logic/statu [0],\biu/cache_ctrl_logic/n204_lutinv }),
    .d({\biu/cache_ctrl_logic/n204_lutinv ,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .f({_al_u3224_o,_al_u4403_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*D))"),
    //.LUTF1("(C*~(~B*D))"),
    //.LUTG0("(C*~(~B*D))"),
    //.LUTG1("(C*~(~B*D))"),
    .INIT_LUTF0(16'b1100000011110000),
    .INIT_LUTF1(16'b1100000011110000),
    .INIT_LUTG0(16'b1100000011110000),
    .INIT_LUTG1(16'b1100000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3225|_al_u3235  (
    .b({_al_u3224_o,_al_u3224_o}),
    .c({addr_ex[9],addr_ex[1]}),
    .d({_al_u3222_o,_al_u3222_o}),
    .f({\biu/cache_ctrl_logic/off [9],\biu/cache_ctrl_logic/off [1]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~B*D))"),
    //.LUT1("(C*~(~B*D))"),
    .INIT_LUT0(16'b1100000011110000),
    .INIT_LUT1(16'b1100000011110000),
    .MODE("LOGIC"))
    \_al_u3226|_al_u3236  (
    .b({_al_u3224_o,_al_u3224_o}),
    .c({addr_ex[8],addr_ex[0]}),
    .d({_al_u3222_o,_al_u3222_o}),
    .f({\biu/cache_ctrl_logic/off [8],\biu/cache_ctrl_logic/off [0]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(C*~(~B*D))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(C*~(~B*D))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100000011110000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3227|_al_u5787  (
    .b({_al_u3224_o,_al_u2705_o}),
    .c({addr_ex[7],\biu/bus_unit/mmu_hwdata [36]}),
    .d({_al_u3222_o,_al_u5786_o}),
    .f({\biu/cache_ctrl_logic/off [7],hwdata_pad[36]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(C*~(~B*D))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1100000011110000),
    .MODE("LOGIC"))
    \_al_u3228|_al_u5783  (
    .b({_al_u3224_o,_al_u2705_o}),
    .c({addr_ex[6],\biu/bus_unit/mmu_hwdata [37]}),
    .d({_al_u3222_o,_al_u5782_o}),
    .f({\biu/cache_ctrl_logic/off [6],hwdata_pad[37]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(C*~(~B*D))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1100000011110000),
    .MODE("LOGIC"))
    \_al_u3229|_al_u5771  (
    .b({_al_u3224_o,_al_u2705_o}),
    .c({addr_ex[5],\biu/bus_unit/mmu_hwdata [40]}),
    .d({_al_u3222_o,_al_u5770_o}),
    .f({\biu/cache_ctrl_logic/off [5],hwdata_pad[40]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(C*~(~B*D))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(C*~(~B*D))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100000011110000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3230|_al_u5767  (
    .b({_al_u3224_o,_al_u2705_o}),
    .c({addr_ex[4],\biu/bus_unit/mmu_hwdata [41]}),
    .d({_al_u3222_o,_al_u5766_o}),
    .f({\biu/cache_ctrl_logic/off [4],hwdata_pad[41]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(C*~(~B*D))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(C*~(~B*D))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100000011110000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3231|_al_u5763  (
    .b({_al_u3224_o,_al_u2705_o}),
    .c({addr_ex[3],\biu/bus_unit/mmu_hwdata [42]}),
    .d({_al_u3222_o,_al_u5762_o}),
    .f({\biu/cache_ctrl_logic/off [3],hwdata_pad[42]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(C*~(~B*D))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1100000011110000),
    .MODE("LOGIC"))
    \_al_u3232|_al_u5759  (
    .b({_al_u3224_o,_al_u2705_o}),
    .c({addr_ex[2],\biu/bus_unit/mmu_hwdata [43]}),
    .d({_al_u3222_o,_al_u5758_o}),
    .f({\biu/cache_ctrl_logic/off [2],hwdata_pad[43]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(C*~(~B*D))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1100000011110000),
    .MODE("LOGIC"))
    \_al_u3233|_al_u5755  (
    .b({_al_u3224_o,_al_u2705_o}),
    .c({addr_ex[11],\biu/bus_unit/mmu_hwdata [44]}),
    .d({_al_u3222_o,_al_u5754_o}),
    .f({\biu/cache_ctrl_logic/off [11],hwdata_pad[44]}));
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*~(~B*D))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*~(~B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1100000011110000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1100000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3234|exu/reg5_b10  (
    .b({_al_u3224_o,addr_ex[10]}),
    .c({addr_ex[10],ex_exc_code[10]}),
    .clk(clk_pad),
    .d({_al_u3222_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\biu/cache_ctrl_logic/off [10],open_n10864}),
    .q({open_n10868,wb_exc_code[10]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3237|cu_ru/m_s_ie/mtie_reg  (
    .b({\cu_ru/m_sip [7],\cu_ru/sepc [7]}),
    .c({\cu_ru/mie ,data_csr[7]}),
    .ce(\cu_ru/m_s_ie/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_sie [7],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n10874,data_csr[7]}),
    .sr(rst_pad),
    .f({_al_u3237_o,_al_u5365_o}),
    .q({open_n10889,\cu_ru/m_sie [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3238|cu_ru/m_s_ie/msie_reg  (
    .a({open_n10890,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/m_sip [3],\cu_ru/trap_target_m }),
    .c({\cu_ru/mie ,\cu_ru/mepc [3]}),
    .ce(\cu_ru/m_s_ie/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_sie [3],data_csr[3]}),
    .mi({open_n10901,data_csr[3]}),
    .sr(rst_pad),
    .f({_al_u3238_o,_al_u6630_o}),
    .q({open_n10905,\cu_ru/m_sie [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3239|_al_u4140  (
    .a({open_n10906,_al_u4132_o}),
    .b({open_n10907,_al_u4138_o}),
    .c({_al_u3238_o,_al_u3238_o}),
    .d({_al_u3237_o,_al_u4139_o}),
    .f({\cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ,_al_u4140_o}));
  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(~D*C*B))"),
    //.LUTF1("(A*~(~D*C*B))"),
    //.LUTG0("(~A*~(~D*C*B))"),
    //.LUTG1("(A*~(~D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010100010101),
    .INIT_LUTF1(16'b1010101000101010),
    .INIT_LUTG0(16'b0101010100010101),
    .INIT_LUTG1(16'b1010101000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3240|cu_ru/mideleg_int_ctrl/dsti_reg  (
    .a({\cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ,\cu_ru/mideleg_int_ctrl/sti_ack_s }),
    .b({\cu_ru/m_sip [5],\cu_ru/m_sip [5]}),
    .c({\cu_ru/mie ,\cu_ru/mie }),
    .ce(\cu_ru/mideleg_int_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mideleg [5],\cu_ru/mideleg [5]}),
    .mi({open_n10935,data_csr[5]}),
    .sr(rst_pad),
    .f({_al_u3240_o,_al_u4131_o}),
    .q({open_n10950,\cu_ru/mideleg [5]}));  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~D*C*~(~B*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000011100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3241|cu_ru/mideleg_int_ctrl/dsei_reg  (
    .a({s_ext_int_pad,open_n10951}),
    .b({\cu_ru/m_s_ip/seip ,_al_u3204_o}),
    .c({\cu_ru/mie ,_al_u3184_o}),
    .ce(\cu_ru/mideleg_int_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mideleg [9],_al_u3195_o}),
    .mi({open_n10962,data_csr[9]}),
    .sr(rst_pad),
    .f({\cu_ru/mideleg_int_ctrl/sei_ack_m ,\cu_ru/mideleg_int_ctrl/n0 }),
    .q({open_n10966,\cu_ru/mideleg [9]}));  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~A*~(~D*C*B))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~A*~(~D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0101010100010101),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0101010100010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3242|cu_ru/mideleg_int_ctrl/dssi_reg  (
    .a({\cu_ru/mideleg_int_ctrl/sei_ack_m ,_al_u6763_o}),
    .b({\cu_ru/m_sip [1],\cu_ru/read_mideleg_sel_lutinv }),
    .c({\cu_ru/mie ,\cu_ru/minstret [1]}),
    .ce(\cu_ru/mideleg_int_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mideleg [1],\cu_ru/mideleg [1]}),
    .mi({open_n10970,data_csr[1]}),
    .sr(rst_pad),
    .f({_al_u3242_o,_al_u7869_o}),
    .q({open_n10985,\cu_ru/mideleg [1]}));  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3243|_al_u4130  (
    .c({_al_u3242_o,_al_u3242_o}),
    .d({_al_u3240_o,\cu_ru/mideleg_int_ctrl/n29_lutinv }),
    .f({\cu_ru/mideleg_int_ctrl/n28_lutinv ,\cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*A)"),
    //.LUTF1("(D*B*~(~C*~A))"),
    //.LUTG0("~(~D*~C*B*A)"),
    //.LUTG1("(D*B*~(~C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110111),
    .INIT_LUTF1(16'b1100100000000000),
    .INIT_LUTG0(16'b1111111111110111),
    .INIT_LUTG1(16'b1100100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3244|cu_ru/m_s_ie/seie_reg  (
    .a({s_ext_int_pad,_al_u3191_o}),
    .b({\cu_ru/m_sie [9],_al_u3194_o}),
    .c({\cu_ru/m_s_ip/seip ,csr_index[10]}),
    .ce(\cu_ru/m_s_ie/u11_sel_is_0_o ),
    .clk(clk_pad),
    .d({\cu_ru/mideleg [9],csr_index[11]}),
    .mi({open_n11013,data_csr[9]}),
    .sr(rst_pad),
    .f({_al_u3244_o,\cu_ru/m_s_ie/u11_sel_is_0_o }),
    .q({open_n11028,\cu_ru/m_sie [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~A*~(D*C*B))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~A*~(D*C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001010101010101),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3245|cu_ru/m_s_ie/ssie_reg  (
    .a({_al_u3244_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/m_sie [1],\cu_ru/trap_target_m }),
    .c({\cu_ru/m_sip [1],\cu_ru/mepc [1]}),
    .ce(\cu_ru/m_s_ie/u11_sel_is_0_o ),
    .clk(clk_pad),
    .d({\cu_ru/mideleg [1],data_csr[1]}),
    .mi({open_n11032,data_csr[1]}),
    .sr(rst_pad),
    .f({_al_u3245_o,_al_u6674_o}),
    .q({open_n11047,\cu_ru/m_sie [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*~B*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"))
    \_al_u3247|_al_u6940  (
    .b({\cu_ru/m_s_status/n5 [1],open_n11050}),
    .c({\cu_ru/mstatus [1],\cu_ru/mstatus [1]}),
    .d({_al_u3245_o,\cu_ru/m_s_status/n2 }),
    .f({\cu_ru/mideleg_int_ctrl/n29_lutinv ,_al_u6940_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3248|cu_ru/m_s_ie/stie_reg  (
    .b({\cu_ru/m_sip [5],\cu_ru/sepc [5]}),
    .c({\cu_ru/mideleg [5],data_csr[5]}),
    .ce(\cu_ru/m_s_ie/u11_sel_is_0_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_sie [5],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n11076,data_csr[5]}),
    .sr(rst_pad),
    .f({_al_u3248_o,_al_u5429_o}),
    .q({open_n11091,\cu_ru/m_sie [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*B*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3249|_al_u6750  (
    .b({_al_u3248_o,open_n11094}),
    .c({\cu_ru/mstatus [1],priv[3]}),
    .d({\cu_ru/m_s_status/n5 [1],\cu_ru/m_s_status/n5 [1]}),
    .f({\cu_ru/mideleg_int_ctrl/sti_ack_s ,_al_u6750_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3254|cu_ru/m_cycle_event/reg1_b9  (
    .b({\cu_ru/mcountinhibit ,_al_u3254_o}),
    .c({\cu_ru/mcycle [9],data_csr[9]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [9],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3254_o,open_n11138}),
    .q({open_n11142,\cu_ru/mcycle [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3256|cu_ru/m_cycle_event/reg1_b8  (
    .b({\cu_ru/mcountinhibit ,_al_u3256_o}),
    .c({\cu_ru/mcycle [8],data_csr[8]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [8],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3256_o,open_n11158}),
    .q({open_n11162,\cu_ru/mcycle [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3258|cu_ru/m_cycle_event/reg1_b7  (
    .b({\cu_ru/mcountinhibit ,_al_u3258_o}),
    .c({\cu_ru/mcycle [7],data_csr[7]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [7],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3258_o,open_n11182}),
    .q({open_n11186,\cu_ru/mcycle [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~B)*~(D*~A))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~(C*~B)*~(D*~A))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000101011001111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1000101011001111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3260|cu_ru/m_cycle_event/reg0_b63  (
    .a({open_n11187,_al_u6788_o}),
    .b({\cu_ru/mcountinhibit ,_al_u6763_o}),
    .c({\cu_ru/mcycle [63],\cu_ru/minstret [63]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [63],\cu_ru/mcycle [63]}),
    .mi({open_n11191,\cu_ru/m_cycle_event/n4 [63]}),
    .sr(rst_pad),
    .f({_al_u3260_o,_al_u6954_o}),
    .q({open_n11206,\cu_ru/minstret [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3262|cu_ru/m_cycle_event/reg1_b62  (
    .b({\cu_ru/mcountinhibit ,_al_u3262_o}),
    .c({\cu_ru/mcycle [62],data_csr[62]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [62],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3262_o,open_n11226}),
    .q({open_n11230,\cu_ru/mcycle [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3264|cu_ru/m_cycle_event/reg1_b61  (
    .b({\cu_ru/mcountinhibit ,_al_u3264_o}),
    .c({\cu_ru/mcycle [61],data_csr[61]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [61],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3264_o,open_n11250}),
    .q({open_n11254,\cu_ru/mcycle [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3266|cu_ru/m_cycle_event/reg1_b60  (
    .b({\cu_ru/mcountinhibit ,_al_u3266_o}),
    .c({\cu_ru/mcycle [60],data_csr[60]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [60],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3266_o,open_n11270}),
    .q({open_n11274,\cu_ru/mcycle [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3268|cu_ru/m_cycle_event/reg1_b6  (
    .b({\cu_ru/mcountinhibit ,_al_u3268_o}),
    .c({\cu_ru/mcycle [6],data_csr[6]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [6],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3268_o,open_n11290}),
    .q({open_n11294,\cu_ru/mcycle [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3270|cu_ru/m_cycle_event/reg1_b59  (
    .b({\cu_ru/mcountinhibit ,_al_u3270_o}),
    .c({\cu_ru/mcycle [59],data_csr[59]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [59],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3270_o,open_n11314}),
    .q({open_n11318,\cu_ru/mcycle [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3272|cu_ru/m_cycle_event/reg1_b58  (
    .b({\cu_ru/mcountinhibit ,_al_u3272_o}),
    .c({\cu_ru/mcycle [58],data_csr[58]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [58],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3272_o,open_n11334}),
    .q({open_n11338,\cu_ru/mcycle [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3274|cu_ru/m_cycle_event/reg1_b57  (
    .b({\cu_ru/mcountinhibit ,_al_u3274_o}),
    .c({\cu_ru/mcycle [57],data_csr[57]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [57],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3274_o,open_n11354}),
    .q({open_n11358,\cu_ru/mcycle [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3276|cu_ru/m_cycle_event/reg1_b56  (
    .b({\cu_ru/mcountinhibit ,_al_u3276_o}),
    .c({\cu_ru/mcycle [56],data_csr[56]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [56],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3276_o,open_n11374}),
    .q({open_n11378,\cu_ru/mcycle [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3278|cu_ru/m_cycle_event/reg1_b55  (
    .b({\cu_ru/mcountinhibit ,_al_u3278_o}),
    .c({\cu_ru/mcycle [55],data_csr[55]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [55],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3278_o,open_n11398}),
    .q({open_n11402,\cu_ru/mcycle [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3280|cu_ru/m_cycle_event/reg1_b54  (
    .b({\cu_ru/mcountinhibit ,_al_u3280_o}),
    .c({\cu_ru/mcycle [54],data_csr[54]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [54],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3280_o,open_n11422}),
    .q({open_n11426,\cu_ru/mcycle [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3282|cu_ru/m_cycle_event/reg1_b53  (
    .b({\cu_ru/mcountinhibit ,_al_u3282_o}),
    .c({\cu_ru/mcycle [53],data_csr[53]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [53],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3282_o,open_n11446}),
    .q({open_n11450,\cu_ru/mcycle [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3284|cu_ru/m_cycle_event/reg1_b52  (
    .b({\cu_ru/mcountinhibit ,_al_u3284_o}),
    .c({\cu_ru/mcycle [52],data_csr[52]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [52],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3284_o,open_n11470}),
    .q({open_n11474,\cu_ru/mcycle [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3286|cu_ru/m_cycle_event/reg1_b51  (
    .b({\cu_ru/mcountinhibit ,_al_u3286_o}),
    .c({\cu_ru/mcycle [51],data_csr[51]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [51],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3286_o,open_n11490}),
    .q({open_n11494,\cu_ru/mcycle [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3288|cu_ru/m_cycle_event/reg1_b50  (
    .b({\cu_ru/mcountinhibit ,_al_u3288_o}),
    .c({\cu_ru/mcycle [50],data_csr[50]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [50],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3288_o,open_n11510}),
    .q({open_n11514,\cu_ru/mcycle [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3290|cu_ru/m_cycle_event/reg1_b5  (
    .b({\cu_ru/mcountinhibit ,_al_u3290_o}),
    .c({\cu_ru/mcycle [5],data_csr[5]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [5],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3290_o,open_n11530}),
    .q({open_n11534,\cu_ru/mcycle [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3292|cu_ru/m_cycle_event/reg1_b49  (
    .b({\cu_ru/mcountinhibit ,_al_u3292_o}),
    .c({\cu_ru/mcycle [49],data_csr[49]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [49],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3292_o,open_n11554}),
    .q({open_n11558,\cu_ru/mcycle [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3294|cu_ru/m_cycle_event/reg1_b48  (
    .b({\cu_ru/mcountinhibit ,_al_u3294_o}),
    .c({\cu_ru/mcycle [48],data_csr[48]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [48],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3294_o,open_n11574}),
    .q({open_n11578,\cu_ru/mcycle [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3296|cu_ru/m_cycle_event/reg1_b47  (
    .b({\cu_ru/mcountinhibit ,_al_u3296_o}),
    .c({\cu_ru/mcycle [47],data_csr[47]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [47],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3296_o,open_n11594}),
    .q({open_n11598,\cu_ru/mcycle [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3298|cu_ru/m_cycle_event/reg1_b46  (
    .b({\cu_ru/mcountinhibit ,_al_u3298_o}),
    .c({\cu_ru/mcycle [46],data_csr[46]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [46],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3298_o,open_n11618}),
    .q({open_n11622,\cu_ru/mcycle [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3300|cu_ru/m_cycle_event/reg1_b45  (
    .b({\cu_ru/mcountinhibit ,_al_u3300_o}),
    .c({\cu_ru/mcycle [45],data_csr[45]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [45],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3300_o,open_n11642}),
    .q({open_n11646,\cu_ru/mcycle [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3302|cu_ru/m_cycle_event/reg1_b44  (
    .b({\cu_ru/mcountinhibit ,_al_u3302_o}),
    .c({\cu_ru/mcycle [44],data_csr[44]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [44],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3302_o,open_n11662}),
    .q({open_n11666,\cu_ru/mcycle [44]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~B)*~(D*~A))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~(C*~B)*~(D*~A))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000101011001111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1000101011001111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3304|cu_ru/m_cycle_event/reg0_b43  (
    .a({open_n11667,_al_u6788_o}),
    .b({\cu_ru/mcountinhibit ,_al_u6763_o}),
    .c({\cu_ru/mcycle [43],\cu_ru/minstret [43]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [43],\cu_ru/mcycle [43]}),
    .mi({open_n11671,\cu_ru/m_cycle_event/n4 [43]}),
    .sr(rst_pad),
    .f({_al_u3304_o,_al_u6994_o}),
    .q({open_n11686,\cu_ru/minstret [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3306|cu_ru/m_cycle_event/reg1_b42  (
    .b({\cu_ru/mcountinhibit ,_al_u3306_o}),
    .c({\cu_ru/mcycle [42],data_csr[42]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [42],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3306_o,open_n11702}),
    .q({open_n11706,\cu_ru/mcycle [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3308|cu_ru/m_cycle_event/reg1_b41  (
    .b({\cu_ru/mcountinhibit ,_al_u3308_o}),
    .c({\cu_ru/mcycle [41],data_csr[41]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [41],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3308_o,open_n11722}),
    .q({open_n11726,\cu_ru/mcycle [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3310|cu_ru/m_cycle_event/reg1_b40  (
    .b({\cu_ru/mcountinhibit ,_al_u3310_o}),
    .c({\cu_ru/mcycle [40],data_csr[40]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [40],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3310_o,open_n11746}),
    .q({open_n11750,\cu_ru/mcycle [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3312|cu_ru/m_cycle_event/reg1_b4  (
    .b({\cu_ru/mcountinhibit ,_al_u3312_o}),
    .c({\cu_ru/mcycle [4],data_csr[4]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [4],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3312_o,open_n11770}),
    .q({open_n11774,\cu_ru/mcycle [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3314|cu_ru/m_cycle_event/reg1_b39  (
    .b({\cu_ru/mcountinhibit ,_al_u3314_o}),
    .c({\cu_ru/mcycle [39],data_csr[39]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [39],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3314_o,open_n11794}),
    .q({open_n11798,\cu_ru/mcycle [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3316|cu_ru/m_cycle_event/reg1_b38  (
    .b({\cu_ru/mcountinhibit ,_al_u3316_o}),
    .c({\cu_ru/mcycle [38],data_csr[38]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [38],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3316_o,open_n11814}),
    .q({open_n11818,\cu_ru/mcycle [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3318|cu_ru/m_cycle_event/reg1_b37  (
    .b({\cu_ru/mcountinhibit ,_al_u3318_o}),
    .c({\cu_ru/mcycle [37],data_csr[37]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [37],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3318_o,open_n11834}),
    .q({open_n11838,\cu_ru/mcycle [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3320|cu_ru/m_cycle_event/reg1_b36  (
    .b({\cu_ru/mcountinhibit ,_al_u3320_o}),
    .c({\cu_ru/mcycle [36],data_csr[36]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [36],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3320_o,open_n11858}),
    .q({open_n11862,\cu_ru/mcycle [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3322|cu_ru/m_cycle_event/reg1_b35  (
    .b({\cu_ru/mcountinhibit ,_al_u3322_o}),
    .c({\cu_ru/mcycle [35],data_csr[35]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [35],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3322_o,open_n11882}),
    .q({open_n11886,\cu_ru/mcycle [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3324|cu_ru/m_cycle_event/reg1_b34  (
    .b({\cu_ru/mcountinhibit ,_al_u3324_o}),
    .c({\cu_ru/mcycle [34],data_csr[34]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [34],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3324_o,open_n11902}),
    .q({open_n11906,\cu_ru/mcycle [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3326|cu_ru/m_cycle_event/reg1_b33  (
    .b({\cu_ru/mcountinhibit ,_al_u3326_o}),
    .c({\cu_ru/mcycle [33],data_csr[33]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [33],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3326_o,open_n11922}),
    .q({open_n11926,\cu_ru/mcycle [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3328|cu_ru/m_cycle_event/reg1_b32  (
    .b({\cu_ru/mcountinhibit ,_al_u3328_o}),
    .c({\cu_ru/mcycle [32],data_csr[32]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [32],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3328_o,open_n11946}),
    .q({open_n11950,\cu_ru/mcycle [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3330|cu_ru/m_cycle_event/reg1_b31  (
    .b({\cu_ru/mcountinhibit ,_al_u3330_o}),
    .c({\cu_ru/mcycle [31],data_csr[31]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [31],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3330_o,open_n11966}),
    .q({open_n11970,\cu_ru/mcycle [31]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3332|cu_ru/m_cycle_event/reg1_b30  (
    .b({\cu_ru/mcountinhibit ,_al_u3332_o}),
    .c({\cu_ru/mcycle [30],data_csr[30]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [30],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3332_o,open_n11990}),
    .q({open_n11994,\cu_ru/mcycle [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3334|cu_ru/m_cycle_event/reg1_b3  (
    .b({\cu_ru/mcountinhibit ,_al_u3334_o}),
    .c({\cu_ru/mcycle [3],data_csr[3]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [3],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3334_o,open_n12010}),
    .q({open_n12014,\cu_ru/mcycle [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3336|cu_ru/m_cycle_event/reg1_b29  (
    .b({\cu_ru/mcountinhibit ,_al_u3336_o}),
    .c({\cu_ru/mcycle [29],data_csr[29]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [29],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3336_o,open_n12034}),
    .q({open_n12038,\cu_ru/mcycle [29]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3338|cu_ru/m_cycle_event/reg1_b28  (
    .b({\cu_ru/mcountinhibit ,_al_u3338_o}),
    .c({\cu_ru/mcycle [28],data_csr[28]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [28],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3338_o,open_n12054}),
    .q({open_n12058,\cu_ru/mcycle [28]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3340|cu_ru/m_cycle_event/reg1_b27  (
    .b({\cu_ru/mcountinhibit ,_al_u3340_o}),
    .c({\cu_ru/mcycle [27],data_csr[27]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [27],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3340_o,open_n12078}),
    .q({open_n12082,\cu_ru/mcycle [27]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3342|cu_ru/m_cycle_event/reg1_b26  (
    .b({\cu_ru/mcountinhibit ,_al_u3342_o}),
    .c({\cu_ru/mcycle [26],data_csr[26]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [26],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3342_o,open_n12098}),
    .q({open_n12102,\cu_ru/mcycle [26]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3344|cu_ru/m_cycle_event/reg1_b25  (
    .b({\cu_ru/mcountinhibit ,_al_u3344_o}),
    .c({\cu_ru/mcycle [25],data_csr[25]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [25],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3344_o,open_n12118}),
    .q({open_n12122,\cu_ru/mcycle [25]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3346|cu_ru/m_cycle_event/reg1_b24  (
    .b({\cu_ru/mcountinhibit ,_al_u3346_o}),
    .c({\cu_ru/mcycle [24],data_csr[24]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [24],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3346_o,open_n12142}),
    .q({open_n12146,\cu_ru/mcycle [24]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3348|cu_ru/m_cycle_event/reg1_b23  (
    .b({\cu_ru/mcountinhibit ,_al_u3348_o}),
    .c({\cu_ru/mcycle [23],data_csr[23]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [23],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3348_o,open_n12166}),
    .q({open_n12170,\cu_ru/mcycle [23]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3350|cu_ru/m_cycle_event/reg1_b22  (
    .b({\cu_ru/mcountinhibit ,_al_u3350_o}),
    .c({\cu_ru/mcycle [22],data_csr[22]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [22],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3350_o,open_n12190}),
    .q({open_n12194,\cu_ru/mcycle [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3352|cu_ru/m_cycle_event/reg1_b21  (
    .b({\cu_ru/mcountinhibit ,_al_u3352_o}),
    .c({\cu_ru/mcycle [21],data_csr[21]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [21],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3352_o,open_n12210}),
    .q({open_n12214,\cu_ru/mcycle [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3354|cu_ru/m_cycle_event/reg1_b20  (
    .b({\cu_ru/mcountinhibit ,_al_u3354_o}),
    .c({\cu_ru/mcycle [20],data_csr[20]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [20],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3354_o,open_n12230}),
    .q({open_n12234,\cu_ru/mcycle [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3356|cu_ru/m_cycle_event/reg1_b2  (
    .b({\cu_ru/mcountinhibit ,_al_u3356_o}),
    .c({\cu_ru/mcycle [2],data_csr[2]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [2],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3356_o,open_n12250}),
    .q({open_n12254,\cu_ru/mcycle [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3358|cu_ru/m_cycle_event/reg1_b19  (
    .b({\cu_ru/mcountinhibit ,_al_u3358_o}),
    .c({\cu_ru/mcycle [19],data_csr[19]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [19],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3358_o,open_n12274}),
    .q({open_n12278,\cu_ru/mcycle [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3360|cu_ru/m_cycle_event/reg1_b18  (
    .b({\cu_ru/mcountinhibit ,_al_u3360_o}),
    .c({\cu_ru/mcycle [18],data_csr[18]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [18],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3360_o,open_n12298}),
    .q({open_n12302,\cu_ru/mcycle [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3362|cu_ru/m_cycle_event/reg1_b17  (
    .b({\cu_ru/mcountinhibit ,_al_u3362_o}),
    .c({\cu_ru/mcycle [17],data_csr[17]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [17],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3362_o,open_n12318}),
    .q({open_n12322,\cu_ru/mcycle [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3364|cu_ru/m_cycle_event/reg1_b16  (
    .b({\cu_ru/mcountinhibit ,_al_u3364_o}),
    .c({\cu_ru/mcycle [16],data_csr[16]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [16],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3364_o,open_n12338}),
    .q({open_n12342,\cu_ru/mcycle [16]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3366|cu_ru/m_cycle_event/reg1_b15  (
    .b({\cu_ru/mcountinhibit ,_al_u3366_o}),
    .c({\cu_ru/mcycle [15],data_csr[15]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [15],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3366_o,open_n12358}),
    .q({open_n12362,\cu_ru/mcycle [15]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3368|cu_ru/m_cycle_event/reg1_b14  (
    .b({\cu_ru/mcountinhibit ,_al_u3368_o}),
    .c({\cu_ru/mcycle [14],data_csr[14]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [14],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3368_o,open_n12378}),
    .q({open_n12382,\cu_ru/mcycle [14]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3370|cu_ru/m_cycle_event/reg1_b13  (
    .b({\cu_ru/mcountinhibit ,_al_u3370_o}),
    .c({\cu_ru/mcycle [13],data_csr[13]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [13],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3370_o,open_n12402}),
    .q({open_n12406,\cu_ru/mcycle [13]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3372|cu_ru/m_cycle_event/reg1_b12  (
    .b({\cu_ru/mcountinhibit ,_al_u3372_o}),
    .c({\cu_ru/mcycle [12],data_csr[12]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [12],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3372_o,open_n12426}),
    .q({open_n12430,\cu_ru/mcycle [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3374|cu_ru/m_cycle_event/reg1_b11  (
    .b({\cu_ru/mcountinhibit ,_al_u3374_o}),
    .c({\cu_ru/mcycle [11],data_csr[11]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [11],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3374_o,open_n12450}),
    .q({open_n12454,\cu_ru/mcycle [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3376|cu_ru/m_cycle_event/reg1_b10  (
    .b({\cu_ru/mcountinhibit ,_al_u3376_o}),
    .c({\cu_ru/mcycle [10],data_csr[10]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [10],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3376_o,open_n12474}),
    .q({open_n12478,\cu_ru/mcycle [10]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3378|cu_ru/m_cycle_event/reg1_b1  (
    .b({\cu_ru/mcountinhibit ,_al_u3378_o}),
    .c({\cu_ru/mcycle [1],data_csr[1]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [1],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3378_o,open_n12494}),
    .q({open_n12498,\cu_ru/mcycle [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3380|cu_ru/m_cycle_event/reg1_b0  (
    .b({\cu_ru/mcountinhibit ,_al_u3380_o}),
    .c({\cu_ru/mcycle [0],data_csr[0]}),
    .clk(clk_pad),
    .d({\cu_ru/m_cycle_event/n2 [0],_al_u3253_o}),
    .sr(rst_pad),
    .f({_al_u3380_o,open_n12518}),
    .q({open_n12522,\cu_ru/mcycle [0]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3382|ins_dec/id_jmp_reg  (
    .b({_al_u2938_o,open_n12525}),
    .c({_al_u3212_o,_al_u3382_o}),
    .ce(\ins_dec/u461_sel_is_0_o ),
    .clk(clk_pad),
    .d({_al_u2933_o,_al_u3214_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3382_o,\ins_dec/n302 }),
    .q({open_n12541,ex_jmp}));  // ../../RTL/CPU/ID/ins_dec.v(830)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3386|ins_dec/reg1_b9  (
    .b({open_n12544,1'b0}),
    .c({id_ins[28],\ins_fetch/ins_hold [29]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[29],\ins_fetch/ins_shift [29]}),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/n80_lutinv ,id_ins[29]}),
    .q({open_n12560,ex_csr_index[9]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(~D*~C)*~(~B*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1110111011100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3387|ins_dec/reg1_b7  (
    .a({_al_u2667_o,open_n12561}),
    .b({_al_u2668_o,open_n12562}),
    .c({_al_u2670_o,_al_u2668_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u2671_o,_al_u2667_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3387_o,id_ins[27]}),
    .q({open_n12578,ex_csr_index[7]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(~(~D*~C)*~(~B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b1110111011100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3388|exu/reg6_b11  (
    .a({_al_u2659_o,open_n12579}),
    .b({_al_u2660_o,csr_index[11]}),
    .c({_al_u2662_o,csr_index[9]}),
    .clk(clk_pad),
    .d({_al_u2663_o,csr_index[10]}),
    .mi({open_n12591,ex_csr_index[11]}),
    .sr(rst_pad),
    .f({_al_u3388_o,_al_u3189_o}),
    .q({open_n12595,csr_index[11]}));  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3389|_al_u2668  (
    .b({_al_u3387_o,open_n12598}),
    .c({_al_u3388_o,\ins_fetch/ins_hold [27]}),
    .d({\ins_dec/n80_lutinv ,1'b0}),
    .f({\ins_dec/funct6_0_lutinv ,_al_u2668_o}));
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3390|ins_dec/reg10_b12  (
    .c({_al_u3384_o,_al_u3384_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/n35_lutinv ,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/funct3_0_lutinv ,open_n12643}),
    .q({open_n12647,ex_exc_code[12]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(~D*~C)*~(~B*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1110111011100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3392|ins_dec/reg1_b4  (
    .a({_al_u2674_o,open_n12648}),
    .b({_al_u2675_o,open_n12649}),
    .c({_al_u2677_o,_al_u2675_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u2678_o,_al_u2674_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3392_o,id_ins[24]}),
    .q({open_n12665,ex_csr_index[4]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3393|ins_dec/reg1_b5  (
    .b({open_n12668,1'b0}),
    .c({_al_u3392_o,\ins_fetch/ins_hold [25]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[25],\ins_fetch/ins_shift [25]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3393_o,id_ins[25]}),
    .q({open_n12684,ex_csr_index[5]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(~D*~C)*~(~B*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1110111011100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3394|ins_dec/reg1_b2  (
    .a({_al_u2680_o,open_n12685}),
    .b({_al_u2681_o,open_n12686}),
    .c({_al_u2683_o,_al_u2681_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u2684_o,_al_u2680_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3394_o,id_ins[22]}),
    .q({open_n12702,ex_csr_index[2]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3395|ins_dec/reg1_b0  (
    .b({id_ins[20],1'b0}),
    .c({_al_u3394_o,\ins_fetch/ins_hold [20]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3393_o,\ins_fetch/ins_shift [20]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3395_o,id_ins[20]}),
    .q({open_n12724,ex_csr_index[0]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*C*~B*~A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3397|ins_dec/reg10_b20  (
    .a({id_ins[25],open_n12725}),
    .b({id_ins[20],open_n12726}),
    .c({_al_u3394_o,id_ins[20]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3392_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3397_o,open_n12743}),
    .q({open_n12747,ex_exc_code[20]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3399|ins_dec/reg10_b29  (
    .c({_al_u3388_o,id_ins[29]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[29],id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3399_o,open_n12768}),
    .q({open_n12772,ex_exc_code[29]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3400|ins_dec/reg1_b8  (
    .b({open_n12775,1'b0}),
    .c({_al_u3387_o,\ins_fetch/ins_hold [28]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[28],\ins_fetch/ins_shift [28]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3400_o,id_ins[28]}),
    .q({open_n12795,ex_csr_index[8]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3401|ins_dec/reg10_b25  (
    .a({id_system,open_n12796}),
    .b({_al_u3399_o,open_n12797}),
    .c({_al_u3400_o,id_ins[25]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[25],id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/ins_sfencevma ,open_n12810}),
    .q({open_n12814,ex_exc_code[25]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u3405|_al_u4765  (
    .c({_al_u3404_o,\biu/bus_unit/mux11_b4_sel_is_2_o }),
    .d({_al_u3403_o,hresp_pad}),
    .f({\biu/bus_unit/mux10_b3_sel_is_0_o ,_al_u4765_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(A*~(D*C*B))"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(A*~(D*C*B))"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0010101010101010),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3406|_al_u6322  (
    .a({\biu/bus_unit/mux10_b3_sel_is_0_o ,_al_u2703_o}),
    .b({_al_u2703_o,hready_pad}),
    .c({\biu/bus_unit/statu [1],\biu/bus_unit/statu [1]}),
    .d({\biu/bus_unit/statu [3],\biu/bus_unit/statu [3]}),
    .f({\biu/bus_unit/mux11_b4_sel_is_2_o ,\biu/cache_write_lutinv }));
  // ../../RTL/CPU/BIU/bus_unit.v(163)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111001001010000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0111001001010000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u3407|biu/bus_unit/reg1_b4  (
    .a({open_n12863,\biu/bus_unit/mux11_b4_sel_is_2_o }),
    .b({\biu/bus_unit/statu [2],_al_u3407_o}),
    .c({\biu/bus_unit/statu [4],hresp_pad}),
    .clk(clk_pad),
    .d({_al_u2889_o,\biu/bus_unit/statu [4]}),
    .sr(\biu/bus_unit/mux17_b4_sel_is_2_o ),
    .f({_al_u3407_o,open_n12881}),
    .q({open_n12885,\biu/bus_unit/statu [4]}));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  EG_PHY_LSLICE #(
    //.LUTF0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0010111000111111),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0010111000111111),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3410|_al_u3412  (
    .a({open_n12886,_al_u3410_o}),
    .b({_al_u2890_o,_al_u2705_o}),
    .c({\biu/bus_unit/n45_lutinv ,_al_u3411_o}),
    .d({\biu/bus_unit/mux10_b3_sel_is_0_o ,hready_pad}),
    .f({_al_u3410_o,\biu/cache_ctrl_logic/n100 [4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*~A)"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~D*C*B*~A)"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b0000000001000000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000001000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3411|_al_u7204  (
    .a({\biu/bus_unit/mmu/statu [0],\biu/bus_unit/mmu/statu [0]}),
    .b({\biu/bus_unit/mmu/statu [1],\biu/bus_unit/mmu/statu [1]}),
    .c({\biu/bus_unit/mmu/statu [2],\biu/bus_unit/mmu/statu [2]}),
    .d({\biu/bus_unit/mmu/statu [3],\biu/bus_unit/mmu/statu [3]}),
    .f({_al_u3411_o,\biu/bus_unit/mmu/n45_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3413|_al_u3942  (
    .c({\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ,_al_u2914_o}),
    .d({\biu/cache_ctrl_logic/n100 [4],\biu/cache_ctrl_logic/n100 [4]}),
    .f({\biu/cache_ctrl_logic/n149 ,\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*C)*~(~B*~A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1110111000001110),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u3415|_al_u7913  (
    .a({open_n12963,_al_u7908_o}),
    .b({open_n12964,_al_u7911_o}),
    .c({ex_size[1],_al_u7912_o}),
    .d({ex_size[0],ex_size[1]}),
    .f({_al_u3415_o,_al_u7913_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("~(~C*D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b1111000011111111),
    .MODE("LOGIC"))
    \_al_u3416|_al_u6324  (
    .b({open_n12987,ex_size[2]}),
    .c({_al_u3415_o,ex_size[3]}),
    .d({_al_u2706_o,_al_u3415_o}),
    .f({hsize_pad[1],\biu/cache_ctrl_logic/n176_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3427|cu_ru/m_s_tvec/reg0_b0  (
    .b({_al_u3186_o,_al_u3186_o}),
    .c({_al_u3194_o,_al_u3194_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u3185_o,_al_u3201_o}),
    .mi({open_n13013,csr_data[0]}),
    .sr(rst_pad),
    .f({_al_u3427_o,\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o }),
    .q({open_n13028,\cu_ru/stvec [0]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTF1("(~D*(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C))"),
    //.LUTG0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTG1("(~D*(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011110011),
    .INIT_LUTF1(16'b0000000010110010),
    .INIT_LUTG0(16'b1100000011110011),
    .INIT_LUTG1(16'b0000000010110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3429|ins_dec/reg5_b63  (
    .a({\exu/alu_au/n12 ,open_n13029}),
    .b({ds1[63],\ins_dec/op_lui_lutinv }),
    .c({ds2[63],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({unsign,_al_u7512_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n15 ,open_n13046}),
    .q({open_n13050,ds1[63]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3431|exu/reg2_b9  (
    .a({_al_u3430_o,\exu/alu_au/n53 [9]}),
    .b({mem_csr_data_max,_al_u3434_o}),
    .c({ds1[9],\exu/alu_au/n55 [9]}),
    .clk(clk_pad),
    .d({ds2[9],\exu/alu_au/n47 [9]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [9],\exu/alu_data_mem_csr [9]}),
    .q({open_n13067,data_csr[9]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3433|_al_u7925  (
    .a({_al_u3432_o,\exu/alu_au/sub_64 [9]}),
    .b({mem_csr_data_or,rd_data_ds1}),
    .c({ds1[9],rd_data_sub}),
    .d({ds2[9],ds1[9]}),
    .f({_al_u3433_o,_al_u7925_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3434|_al_u3436  (
    .a({_al_u3433_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[9],ds1[9]}),
    .d({ds2[9],ds2[9]}),
    .f({_al_u3434_o,\exu/alu_au/n55 [9]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010101010001110),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010101010001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3435|_al_u3461  (
    .a({\exu/alu_au/n5 ,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({ds1[63],mem_csr_data_min}),
    .c({ds2[63],ds1[63]}),
    .d({unsign,ds2[63]}),
    .f({\exu/alu_au/ds1_light_than_ds2_lutinv ,\exu/alu_au/n55 [63]}));
  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3438|ins_dec/mem_csr_data_and_reg  (
    .c({mem_csr_data_and,\ins_dec/n71 }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\exu/alu_au/alu_and [9],_al_u3969_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n47 [9],open_n13156}),
    .q({open_n13160,mem_csr_data_and}));  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3440|exu/reg2_b8  (
    .a({_al_u3430_o,\exu/alu_au/n53 [8]}),
    .b({mem_csr_data_max,_al_u3443_o}),
    .c({ds1[8],\exu/alu_au/n55 [8]}),
    .clk(clk_pad),
    .d({ds2[8],\exu/alu_au/n47 [8]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [8],\exu/alu_data_mem_csr [8]}),
    .q({open_n13177,data_csr[8]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3442|_al_u7946  (
    .a({_al_u3441_o,\exu/alu_au/sub_64 [8]}),
    .b({mem_csr_data_or,rd_data_ds1}),
    .c({ds1[8],rd_data_sub}),
    .d({ds2[8],ds1[8]}),
    .f({_al_u3442_o,_al_u7946_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3443|_al_u3444  (
    .a({_al_u3442_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[8],ds1[8]}),
    .d({ds2[8],ds2[8]}),
    .f({_al_u3443_o,\exu/alu_au/n55 [8]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(C@D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*(C@D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000110011000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000110011000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3446|_al_u3445  (
    .b({open_n13220,ds1[8]}),
    .c({mem_csr_data_and,ds2[8]}),
    .d({\exu/alu_au/alu_and [8],and_clr}),
    .f({\exu/alu_au/n47 [8],\exu/alu_au/alu_and [8]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3448|exu/reg2_b7  (
    .a({_al_u3430_o,\exu/alu_au/n53 [7]}),
    .b({mem_csr_data_max,_al_u3451_o}),
    .c({ds1[7],\exu/alu_au/n55 [7]}),
    .clk(clk_pad),
    .d({ds2[7],\exu/alu_au/n47 [7]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [7],\exu/alu_data_mem_csr [7]}),
    .q({open_n13261,data_csr[7]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3450|_al_u3453  (
    .a({_al_u3449_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[7],ds1[7]}),
    .d({ds2[7],ds2[7]}),
    .f({_al_u3450_o,\exu/alu_au/n47 [7]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3451|_al_u7959  (
    .a({_al_u3450_o,\exu/alu_au/sub_64 [7]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[7],rd_data_sub}),
    .d({ds2[7],ds1[7]}),
    .f({_al_u3451_o,_al_u7959_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001000100111111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001000100111111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3457|_al_u3456  (
    .a({_al_u3456_o,mem_csr_data_ds2}),
    .b({mem_csr_data_xor,mem_csr_data_or}),
    .c({ds1[63],ds1[63]}),
    .d({ds2[63],ds2[63]}),
    .f({_al_u3457_o,_al_u3456_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3459|_al_u3728  (
    .b({\exu/alu_au/add_64 [63],\exu/alu_au/add_64 [32]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3459_o,_al_u3728_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*A*~(D*~C))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010000000100010),
    .MODE("LOGIC"))
    \_al_u3460|_al_u3458  (
    .a({_al_u3457_o,and_clr}),
    .b({\exu/alu_au/n47 [63],mem_csr_data_and}),
    .c({_al_u3459_o,ds1[63]}),
    .d({mem_csr_data_add,ds2[63]}),
    .f({_al_u3460_o,\exu/alu_au/n47 [63]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011110011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1100000011110011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3463|ins_dec/reg5_b62  (
    .a({_al_u3430_o,open_n13372}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[62],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[62],_al_u7516_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [62],open_n13389}),
    .q({open_n13393,ds1[62]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3465|_al_u3469  (
    .a({_al_u3464_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[62],ds1[62]}),
    .d({ds2[62],ds2[62]}),
    .f({_al_u3465_o,\exu/alu_au/n55 [62]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u3467|_al_u3720  (
    .b({\exu/alu_au/add_64 [62],\exu/alu_au/add_64 [33]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3467_o,_al_u3720_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3468|_al_u3466  (
    .a({_al_u3465_o,and_clr}),
    .b({\exu/alu_au/n47 [62],mem_csr_data_and}),
    .c({_al_u3467_o,ds1[62]}),
    .d({mem_csr_data_add,ds2[62]}),
    .f({_al_u3468_o,\exu/alu_au/n47 [62]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011110011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3471|ins_dec/reg5_b61  (
    .a({_al_u3430_o,open_n13464}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[61],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[61],_al_u7520_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [61],open_n13477}),
    .q({open_n13481,ds1[61]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3473|_al_u3477  (
    .a({_al_u3472_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[61],ds1[61]}),
    .d({ds2[61],ds2[61]}),
    .f({_al_u3473_o,\exu/alu_au/n55 [61]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3475|_al_u3712  (
    .b({\exu/alu_au/add_64 [61],\exu/alu_au/add_64 [34]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3475_o,_al_u3712_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3476|_al_u3474  (
    .a({_al_u3473_o,and_clr}),
    .b({\exu/alu_au/n47 [61],mem_csr_data_and}),
    .c({_al_u3475_o,ds1[61]}),
    .d({mem_csr_data_add,ds2[61]}),
    .f({_al_u3476_o,\exu/alu_au/n47 [61]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011110011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3479|ins_dec/reg5_b60  (
    .a({_al_u3430_o,open_n13552}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[60],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[60],_al_u7524_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [60],open_n13565}),
    .q({open_n13569,ds1[60]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3481|_al_u3485  (
    .a({_al_u3480_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[60],ds1[60]}),
    .d({ds2[60],ds2[60]}),
    .f({_al_u3481_o,\exu/alu_au/n55 [60]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u3483|_al_u3704  (
    .b({\exu/alu_au/add_64 [60],\exu/alu_au/add_64 [35]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3483_o,_al_u3704_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"))
    \_al_u3484|_al_u3482  (
    .a({_al_u3481_o,and_clr}),
    .b({\exu/alu_au/n47 [60],mem_csr_data_and}),
    .c({_al_u3483_o,ds1[60]}),
    .d({mem_csr_data_add,ds2[60]}),
    .f({_al_u3484_o,\exu/alu_au/n47 [60]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3487|exu/reg2_b6  (
    .a({_al_u3430_o,\exu/alu_au/n53 [6]}),
    .b({mem_csr_data_max,_al_u3490_o}),
    .c({ds1[6],\exu/alu_au/n55 [6]}),
    .clk(clk_pad),
    .d({ds2[6],\exu/alu_au/n47 [6]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [6],\exu/alu_data_mem_csr [6]}),
    .q({open_n13652,data_csr[6]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3489|_al_u3492  (
    .a({_al_u3488_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[6],ds1[6]}),
    .d({ds2[6],ds2[6]}),
    .f({_al_u3489_o,\exu/alu_au/n47 [6]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3490|_al_u8914  (
    .a({_al_u3489_o,\exu/alu_au/sub_64 [6]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[6],rd_data_sub}),
    .d({ds2[6],ds1[6]}),
    .f({_al_u3490_o,_al_u8914_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3494|ins_dec/reg5_b59  (
    .a({_al_u3430_o,open_n13697}),
    .b({mem_csr_data_max,open_n13698}),
    .c({ds1[59],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[59],_al_u7352_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [59],open_n13711}),
    .q({open_n13715,ds1[59]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3496|_al_u3500  (
    .a({_al_u3495_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[59],ds1[59]}),
    .d({ds2[59],ds2[59]}),
    .f({_al_u3496_o,\exu/alu_au/n55 [59]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3498|_al_u3696  (
    .b({\exu/alu_au/add_64 [59],\exu/alu_au/add_64 [36]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3498_o,_al_u3696_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"))
    \_al_u3499|_al_u3497  (
    .a({_al_u3496_o,and_clr}),
    .b({\exu/alu_au/n47 [59],mem_csr_data_and}),
    .c({_al_u3498_o,ds1[59]}),
    .d({mem_csr_data_add,ds2[59]}),
    .f({_al_u3499_o,\exu/alu_au/n47 [59]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3502|ins_dec/reg5_b58  (
    .a({_al_u3430_o,open_n13786}),
    .b({mem_csr_data_max,open_n13787}),
    .c({ds1[58],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[58],_al_u7356_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [58],open_n13800}),
    .q({open_n13804,ds1[58]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3504|_al_u3508  (
    .a({_al_u3503_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[58],ds1[58]}),
    .d({ds2[58],ds2[58]}),
    .f({_al_u3504_o,\exu/alu_au/n55 [58]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u3506|_al_u3688  (
    .b({\exu/alu_au/add_64 [58],\exu/alu_au/add_64 [37]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3506_o,_al_u3688_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3507|_al_u3505  (
    .a({_al_u3504_o,and_clr}),
    .b({\exu/alu_au/n47 [58],mem_csr_data_and}),
    .c({_al_u3506_o,ds1[58]}),
    .d({mem_csr_data_add,ds2[58]}),
    .f({_al_u3507_o,\exu/alu_au/n47 [58]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3510|ins_dec/reg5_b57  (
    .a({_al_u3430_o,open_n13875}),
    .b({mem_csr_data_max,open_n13876}),
    .c({ds1[57],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[57],_al_u7359_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [57],open_n13893}),
    .q({open_n13897,ds1[57]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3512|_al_u3516  (
    .a({_al_u3511_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[57],ds1[57]}),
    .d({ds2[57],ds2[57]}),
    .f({_al_u3512_o,\exu/alu_au/n55 [57]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3514|_al_u3680  (
    .b({\exu/alu_au/add_64 [57],\exu/alu_au/add_64 [38]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3514_o,_al_u3680_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3515|_al_u3513  (
    .a({_al_u3512_o,and_clr}),
    .b({\exu/alu_au/n47 [57],mem_csr_data_and}),
    .c({_al_u3514_o,ds1[57]}),
    .d({mem_csr_data_add,ds2[57]}),
    .f({_al_u3515_o,\exu/alu_au/n47 [57]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3518|ins_dec/reg5_b56  (
    .a({_al_u3430_o,open_n13968}),
    .b({mem_csr_data_max,open_n13969}),
    .c({ds1[56],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[56],_al_u7362_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [56],open_n13986}),
    .q({open_n13990,ds1[56]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3520|_al_u3524  (
    .a({_al_u3519_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[56],ds1[56]}),
    .d({ds2[56],ds2[56]}),
    .f({_al_u3520_o,\exu/alu_au/n55 [56]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u3522|_al_u3672  (
    .b({\exu/alu_au/add_64 [56],\exu/alu_au/add_64 [39]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3522_o,_al_u3672_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"))
    \_al_u3523|_al_u3521  (
    .a({_al_u3520_o,and_clr}),
    .b({\exu/alu_au/n47 [56],mem_csr_data_and}),
    .c({_al_u3522_o,ds1[56]}),
    .d({mem_csr_data_add,ds2[56]}),
    .f({_al_u3523_o,\exu/alu_au/n47 [56]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3526|ins_dec/reg5_b55  (
    .a({_al_u3430_o,open_n14053}),
    .b({mem_csr_data_max,open_n14054}),
    .c({ds1[55],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[55],_al_u7365_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [55],open_n14067}),
    .q({open_n14071,ds1[55]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3528|_al_u3529  (
    .a({_al_u3527_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[55],ds1[55]}),
    .d({ds2[55],ds2[55]}),
    .f({_al_u3528_o,\exu/alu_au/n47 [55]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3530|_al_u3657  (
    .b({\exu/alu_au/add_64 [55],\exu/alu_au/add_64 [40]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3530_o,_al_u3657_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3531|exu/reg2_b55  (
    .a({_al_u3528_o,open_n14118}),
    .b({\exu/alu_au/n47 [55],_al_u3531_o}),
    .c({_al_u3530_o,\exu/alu_au/n55 [55]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [55]}),
    .sr(rst_pad),
    .f({_al_u3531_o,\exu/alu_data_mem_csr [55]}),
    .q({open_n14135,data_csr[55]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3534|ins_dec/reg5_b54  (
    .a({_al_u3430_o,open_n14136}),
    .b({mem_csr_data_max,open_n14137}),
    .c({ds1[54],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[54],_al_u7368_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [54],open_n14150}),
    .q({open_n14154,ds1[54]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3536|_al_u3537  (
    .a({_al_u3535_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[54],ds1[54]}),
    .d({ds2[54],ds2[54]}),
    .f({_al_u3536_o,\exu/alu_au/n47 [54]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u3538|_al_u3649  (
    .b({\exu/alu_au/add_64 [54],\exu/alu_au/add_64 [41]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3538_o,_al_u3649_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3539|exu/reg2_b54  (
    .a({_al_u3536_o,open_n14201}),
    .b({\exu/alu_au/n47 [54],_al_u3539_o}),
    .c({_al_u3538_o,\exu/alu_au/n55 [54]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [54]}),
    .sr(rst_pad),
    .f({_al_u3539_o,\exu/alu_data_mem_csr [54]}),
    .q({open_n14218,data_csr[54]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3542|ins_dec/reg5_b53  (
    .a({_al_u3430_o,open_n14219}),
    .b({mem_csr_data_max,open_n14220}),
    .c({ds1[53],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[53],_al_u7371_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [53],open_n14237}),
    .q({open_n14241,ds1[53]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3544|_al_u3545  (
    .a({_al_u3543_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[53],ds1[53]}),
    .d({ds2[53],ds2[53]}),
    .f({_al_u3544_o,\exu/alu_au/n47 [53]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3546|_al_u3641  (
    .b({\exu/alu_au/add_64 [53],\exu/alu_au/add_64 [42]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3546_o,_al_u3641_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3547|exu/reg2_b53  (
    .a({_al_u3544_o,open_n14292}),
    .b({\exu/alu_au/n47 [53],_al_u3547_o}),
    .c({_al_u3546_o,\exu/alu_au/n55 [53]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [53]}),
    .sr(rst_pad),
    .f({_al_u3547_o,\exu/alu_data_mem_csr [53]}),
    .q({open_n14313,data_csr[53]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3550|ins_dec/reg5_b52  (
    .a({_al_u3430_o,open_n14314}),
    .b({mem_csr_data_max,open_n14315}),
    .c({ds1[52],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[52],_al_u7374_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [52],open_n14332}),
    .q({open_n14336,ds1[52]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3552|_al_u3553  (
    .a({_al_u3551_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[52],ds1[52]}),
    .d({ds2[52],ds2[52]}),
    .f({_al_u3552_o,\exu/alu_au/n47 [52]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u3554|_al_u3633  (
    .b({\exu/alu_au/add_64 [52],\exu/alu_au/add_64 [43]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3554_o,_al_u3633_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3555|exu/reg2_b52  (
    .a({_al_u3552_o,open_n14379}),
    .b({\exu/alu_au/n47 [52],_al_u3555_o}),
    .c({_al_u3554_o,\exu/alu_au/n55 [52]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [52]}),
    .sr(rst_pad),
    .f({_al_u3555_o,\exu/alu_data_mem_csr [52]}),
    .q({open_n14400,data_csr[52]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3558|ins_dec/reg5_b51  (
    .a({_al_u3430_o,open_n14401}),
    .b({mem_csr_data_max,open_n14402}),
    .c({ds1[51],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[51],_al_u7377_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [51],open_n14415}),
    .q({open_n14419,ds1[51]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3560|_al_u3561  (
    .a({_al_u3559_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[51],ds1[51]}),
    .d({ds2[51],ds2[51]}),
    .f({_al_u3560_o,\exu/alu_au/n47 [51]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3562|_al_u3625  (
    .b({\exu/alu_au/add_64 [51],\exu/alu_au/add_64 [44]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3562_o,_al_u3625_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3563|exu/reg2_b51  (
    .a({_al_u3560_o,open_n14466}),
    .b({\exu/alu_au/n47 [51],_al_u3563_o}),
    .c({_al_u3562_o,\exu/alu_au/n55 [51]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [51]}),
    .sr(rst_pad),
    .f({_al_u3563_o,\exu/alu_data_mem_csr [51]}),
    .q({open_n14483,data_csr[51]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3566|ins_dec/reg5_b50  (
    .a({_al_u3430_o,open_n14484}),
    .b({mem_csr_data_max,open_n14485}),
    .c({ds1[50],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[50],_al_u7380_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [50],open_n14498}),
    .q({open_n14502,ds1[50]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3568|_al_u3569  (
    .a({_al_u3567_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[50],ds1[50]}),
    .d({ds2[50],ds2[50]}),
    .f({_al_u3568_o,\exu/alu_au/n47 [50]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u3570|_al_u3617  (
    .b({\exu/alu_au/add_64 [50],\exu/alu_au/add_64 [45]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3570_o,_al_u3617_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3571|exu/reg2_b50  (
    .a({_al_u3568_o,open_n14549}),
    .b({\exu/alu_au/n47 [50],_al_u3571_o}),
    .c({_al_u3570_o,\exu/alu_au/n55 [50]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [50]}),
    .sr(rst_pad),
    .f({_al_u3571_o,\exu/alu_data_mem_csr [50]}),
    .q({open_n14566,data_csr[50]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3574|exu/reg2_b5  (
    .a({_al_u3430_o,\exu/alu_au/n53 [5]}),
    .b({mem_csr_data_max,_al_u3577_o}),
    .c({ds1[5],\exu/alu_au/n55 [5]}),
    .clk(clk_pad),
    .d({ds2[5],\exu/alu_au/n47 [5]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [5],\exu/alu_data_mem_csr [5]}),
    .q({open_n14583,data_csr[5]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3576|_al_u3579  (
    .a({_al_u3575_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[5],ds1[5]}),
    .d({ds2[5],ds2[5]}),
    .f({_al_u3576_o,\exu/alu_au/n47 [5]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3577|_al_u8951  (
    .a({_al_u3576_o,\exu/alu_au/sub_64 [5]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[5],rd_data_sub}),
    .d({ds2[5],ds1[5]}),
    .f({_al_u3577_o,_al_u8951_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3581|ins_dec/reg5_b49  (
    .a({_al_u3430_o,open_n14632}),
    .b({mem_csr_data_max,open_n14633}),
    .c({ds1[49],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[49],_al_u7383_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [49],open_n14650}),
    .q({open_n14654,ds1[49]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3583|_al_u3584  (
    .a({_al_u3582_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[49],ds1[49]}),
    .d({ds2[49],ds2[49]}),
    .f({_al_u3583_o,\exu/alu_au/n47 [49]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3585|_al_u3609  (
    .b({\exu/alu_au/add_64 [49],\exu/alu_au/add_64 [46]}),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3585_o,_al_u3609_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3586|exu/reg2_b49  (
    .a({_al_u3583_o,open_n14705}),
    .b({\exu/alu_au/n47 [49],_al_u3586_o}),
    .c({_al_u3585_o,\exu/alu_au/n55 [49]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [49]}),
    .sr(rst_pad),
    .f({_al_u3586_o,\exu/alu_data_mem_csr [49]}),
    .q({open_n14726,data_csr[49]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3589|ins_dec/reg5_b48  (
    .a({_al_u3430_o,open_n14727}),
    .b({mem_csr_data_max,open_n14728}),
    .c({ds1[48],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[48],_al_u7386_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [48],open_n14745}),
    .q({open_n14749,ds1[48]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3591|_al_u3592  (
    .a({_al_u3590_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[48],ds1[48]}),
    .d({ds2[48],ds2[48]}),
    .f({_al_u3591_o,\exu/alu_au/n47 [48]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3593|_al_u3601  (
    .b(\exu/alu_au/add_64 [48:47]),
    .c({ex_size[2],ex_size[2]}),
    .d({\exu/alu_au/add_64 [31],\exu/alu_au/add_64 [31]}),
    .f({_al_u3593_o,_al_u3601_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3594|exu/reg2_b48  (
    .a({_al_u3591_o,open_n14796}),
    .b({\exu/alu_au/n47 [48],_al_u3594_o}),
    .c({_al_u3593_o,\exu/alu_au/n55 [48]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [48]}),
    .sr(rst_pad),
    .f({_al_u3594_o,\exu/alu_data_mem_csr [48]}),
    .q({open_n14817,data_csr[48]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3597|ins_dec/reg5_b47  (
    .a({_al_u3430_o,open_n14818}),
    .b({mem_csr_data_max,open_n14819}),
    .c({ds1[47],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[47],_al_u7389_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [47],open_n14832}),
    .q({open_n14836,ds1[47]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3599|_al_u3600  (
    .a({_al_u3598_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[47],ds1[47]}),
    .d({ds2[47],ds2[47]}),
    .f({_al_u3599_o,\exu/alu_au/n47 [47]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3602|exu/reg2_b47  (
    .a({_al_u3599_o,open_n14857}),
    .b({\exu/alu_au/n47 [47],_al_u3602_o}),
    .c({_al_u3601_o,\exu/alu_au/n55 [47]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [47]}),
    .sr(rst_pad),
    .f({_al_u3602_o,\exu/alu_data_mem_csr [47]}),
    .q({open_n14874,data_csr[47]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT_LUT0(16'b1111001101011111),
    .INIT_LUT1(16'b1100010010000000),
    .MODE("LOGIC"))
    \_al_u3603|_al_u4236  (
    .a({\exu/alu_au/ds1_light_than_ds2_lutinv ,\exu/alu_data_mem_csr [55]}),
    .b({mem_csr_data_min,\exu/alu_data_mem_csr [47]}),
    .c({ds1[47],addr_ex[0]}),
    .d({ds2[47],addr_ex[1]}),
    .f({\exu/alu_au/n55 [47],_al_u4236_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3605|ins_dec/reg5_b46  (
    .a({_al_u3430_o,open_n14895}),
    .b({mem_csr_data_max,open_n14896}),
    .c({ds1[46],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[46],_al_u7392_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [46],open_n14909}),
    .q({open_n14913,ds1[46]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3607|_al_u3608  (
    .a({_al_u3606_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[46],ds1[46]}),
    .d({ds2[46],ds2[46]}),
    .f({_al_u3607_o,\exu/alu_au/n47 [46]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3610|exu/reg2_b46  (
    .a({_al_u3607_o,open_n14938}),
    .b({\exu/alu_au/n47 [46],_al_u3610_o}),
    .c({_al_u3609_o,\exu/alu_au/n55 [46]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [46]}),
    .sr(rst_pad),
    .f({_al_u3610_o,\exu/alu_data_mem_csr [46]}),
    .q({open_n14959,data_csr[46]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3613|ins_dec/reg5_b45  (
    .a({_al_u3430_o,open_n14960}),
    .b({mem_csr_data_max,open_n14961}),
    .c({ds1[45],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[45],_al_u7395_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [45],open_n14978}),
    .q({open_n14982,ds1[45]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3615|_al_u3616  (
    .a({_al_u3614_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[45],ds1[45]}),
    .d({ds2[45],ds2[45]}),
    .f({_al_u3615_o,\exu/alu_au/n47 [45]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3618|exu/reg2_b45  (
    .a({_al_u3615_o,open_n15007}),
    .b({\exu/alu_au/n47 [45],_al_u3618_o}),
    .c({_al_u3617_o,\exu/alu_au/n55 [45]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [45]}),
    .sr(rst_pad),
    .f({_al_u3618_o,\exu/alu_data_mem_csr [45]}),
    .q({open_n15028,data_csr[45]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3621|ins_dec/reg5_b44  (
    .a({_al_u3430_o,open_n15029}),
    .b({mem_csr_data_max,open_n15030}),
    .c({ds1[44],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[44],_al_u7398_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [44],open_n15047}),
    .q({open_n15051,ds1[44]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3623|_al_u3624  (
    .a({_al_u3622_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[44],ds1[44]}),
    .d({ds2[44],ds2[44]}),
    .f({_al_u3623_o,\exu/alu_au/n47 [44]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3626|exu/reg2_b44  (
    .a({_al_u3623_o,open_n15072}),
    .b({\exu/alu_au/n47 [44],_al_u3626_o}),
    .c({_al_u3625_o,\exu/alu_au/n55 [44]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [44]}),
    .sr(rst_pad),
    .f({_al_u3626_o,\exu/alu_data_mem_csr [44]}),
    .q({open_n15089,data_csr[44]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011110011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1100000011110011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3629|ins_dec/reg5_b43  (
    .a({_al_u3430_o,open_n15090}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[43],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[43],_al_u7528_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [43],open_n15107}),
    .q({open_n15111,ds1[43]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3631|_al_u3635  (
    .a({_al_u3630_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[43],ds1[43]}),
    .d({ds2[43],ds2[43]}),
    .f({_al_u3631_o,\exu/alu_au/n55 [43]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"))
    \_al_u3634|_al_u3632  (
    .a({_al_u3631_o,and_clr}),
    .b({\exu/alu_au/n47 [43],mem_csr_data_and}),
    .c({_al_u3633_o,ds1[43]}),
    .d({mem_csr_data_add,ds2[43]}),
    .f({_al_u3634_o,\exu/alu_au/n47 [43]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3637|_al_u3640  (
    .a({_al_u3430_o,and_clr}),
    .b({mem_csr_data_max,mem_csr_data_and}),
    .c({ds1[42],ds1[42]}),
    .d({ds2[42],ds2[42]}),
    .f({\exu/alu_au/n53 [42],\exu/alu_au/n47 [42]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3639|_al_u3643  (
    .a({_al_u3638_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[42],ds1[42]}),
    .d({ds2[42],ds2[42]}),
    .f({_al_u3639_o,\exu/alu_au/n55 [42]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3642|exu/reg2_b42  (
    .a({_al_u3639_o,open_n15200}),
    .b({\exu/alu_au/n47 [42],_al_u3642_o}),
    .c({_al_u3641_o,\exu/alu_au/n55 [42]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [42]}),
    .sr(rst_pad),
    .f({_al_u3642_o,\exu/alu_data_mem_csr [42]}),
    .q({open_n15217,data_csr[42]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011110011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1100000011110011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3645|ins_dec/reg5_b41  (
    .a({_al_u3430_o,open_n15218}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[41],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[41],_al_u7535_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [41],open_n15235}),
    .q({open_n15239,ds1[41]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3647|_al_u3648  (
    .a({_al_u3646_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[41],ds1[41]}),
    .d({ds2[41],ds2[41]}),
    .f({_al_u3647_o,\exu/alu_au/n47 [41]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3650|exu/reg2_b41  (
    .a({_al_u3647_o,open_n15264}),
    .b({\exu/alu_au/n47 [41],_al_u3650_o}),
    .c({_al_u3649_o,\exu/alu_au/n55 [41]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [41]}),
    .sr(rst_pad),
    .f({_al_u3650_o,\exu/alu_data_mem_csr [41]}),
    .q({open_n15285,data_csr[41]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011110011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3653|ins_dec/reg5_b40  (
    .a({_al_u3430_o,open_n15286}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[40],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[40],_al_u7539_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [40],open_n15299}),
    .q({open_n15303,ds1[40]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3655|_al_u3656  (
    .a({_al_u3654_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[40],ds1[40]}),
    .d({ds2[40],ds2[40]}),
    .f({_al_u3655_o,\exu/alu_au/n47 [40]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3658|exu/reg2_b40  (
    .a({_al_u3655_o,open_n15324}),
    .b({\exu/alu_au/n47 [40],_al_u3658_o}),
    .c({_al_u3657_o,\exu/alu_au/n55 [40]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [40]}),
    .sr(rst_pad),
    .f({_al_u3658_o,\exu/alu_data_mem_csr [40]}),
    .q({open_n15345,data_csr[40]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3661|exu/reg2_b4  (
    .a({_al_u3430_o,\exu/alu_au/n53 [4]}),
    .b({mem_csr_data_max,_al_u3664_o}),
    .c({ds1[4],\exu/alu_au/n55 [4]}),
    .clk(clk_pad),
    .d({ds2[4],\exu/alu_au/n47 [4]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [4],\exu/alu_data_mem_csr [4]}),
    .q({open_n15366,data_csr[4]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3663|_al_u3666  (
    .a({_al_u3662_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[4],ds1[4]}),
    .d({ds2[4],ds2[4]}),
    .f({_al_u3663_o,\exu/alu_au/n47 [4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3664|_al_u8986  (
    .a({_al_u3663_o,\exu/alu_au/sub_64 [4]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[4],rd_data_sub}),
    .d({ds2[4],ds1[4]}),
    .f({_al_u3664_o,_al_u8986_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011110011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3668|ins_dec/reg5_b39  (
    .a({_al_u3430_o,open_n15411}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[39],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[39],_al_u7555_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [39],open_n15424}),
    .q({open_n15428,ds1[39]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3670|_al_u3671  (
    .a({_al_u3669_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[39],ds1[39]}),
    .d({ds2[39],ds2[39]}),
    .f({_al_u3670_o,\exu/alu_au/n47 [39]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3673|exu/reg2_b39  (
    .a({_al_u3670_o,open_n15449}),
    .b({\exu/alu_au/n47 [39],_al_u3673_o}),
    .c({_al_u3672_o,\exu/alu_au/n55 [39]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [39]}),
    .sr(rst_pad),
    .f({_al_u3673_o,\exu/alu_data_mem_csr [39]}),
    .q({open_n15466,data_csr[39]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011110011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1100000011110011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3676|ins_dec/reg5_b38  (
    .a({_al_u3430_o,open_n15467}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[38],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[38],_al_u7559_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [38],open_n15484}),
    .q({open_n15488,ds1[38]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3678|_al_u3679  (
    .a({_al_u3677_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[38],ds1[38]}),
    .d({ds2[38],ds2[38]}),
    .f({_al_u3678_o,\exu/alu_au/n47 [38]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3681|exu/reg2_b38  (
    .a({_al_u3678_o,open_n15513}),
    .b({\exu/alu_au/n47 [38],_al_u3681_o}),
    .c({_al_u3680_o,\exu/alu_au/n55 [38]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [38]}),
    .sr(rst_pad),
    .f({_al_u3681_o,\exu/alu_data_mem_csr [38]}),
    .q({open_n15534,data_csr[38]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011110011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1100000011110011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3684|ins_dec/reg5_b37  (
    .a({_al_u3430_o,open_n15535}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[37],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[37],_al_u7563_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [37],open_n15552}),
    .q({open_n15556,ds1[37]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3686|_al_u3687  (
    .a({_al_u3685_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[37],ds1[37]}),
    .d({ds2[37],ds2[37]}),
    .f({_al_u3686_o,\exu/alu_au/n47 [37]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3689|exu/reg2_b37  (
    .a({_al_u3686_o,open_n15581}),
    .b({\exu/alu_au/n47 [37],_al_u3689_o}),
    .c({_al_u3688_o,\exu/alu_au/n55 [37]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [37]}),
    .sr(rst_pad),
    .f({_al_u3689_o,\exu/alu_data_mem_csr [37]}),
    .q({open_n15602,data_csr[37]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011110011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3692|ins_dec/reg5_b36  (
    .a({_al_u3430_o,open_n15603}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[36],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[36],_al_u7567_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [36],open_n15616}),
    .q({open_n15620,ds1[36]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3694|_al_u3695  (
    .a({_al_u3693_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[36],ds1[36]}),
    .d({ds2[36],ds2[36]}),
    .f({_al_u3694_o,\exu/alu_au/n47 [36]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3697|exu/reg2_b36  (
    .a({_al_u3694_o,open_n15641}),
    .b({\exu/alu_au/n47 [36],_al_u3697_o}),
    .c({_al_u3696_o,\exu/alu_au/n55 [36]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [36]}),
    .sr(rst_pad),
    .f({_al_u3697_o,\exu/alu_data_mem_csr [36]}),
    .q({open_n15658,data_csr[36]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3700|ins_dec/reg5_b35  (
    .a({_al_u3430_o,open_n15659}),
    .b({mem_csr_data_max,open_n15660}),
    .c({ds1[35],_al_u7353_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[35],_al_u7679_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [35],open_n15673}),
    .q({open_n15677,ds1[35]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3702|_al_u3703  (
    .a({_al_u3701_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[35],ds1[35]}),
    .d({ds2[35],ds2[35]}),
    .f({_al_u3702_o,\exu/alu_au/n47 [35]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3705|exu/reg2_b35  (
    .a({_al_u3702_o,open_n15698}),
    .b({\exu/alu_au/n47 [35],_al_u3705_o}),
    .c({_al_u3704_o,\exu/alu_au/n55 [35]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [35]}),
    .sr(rst_pad),
    .f({_al_u3705_o,\exu/alu_data_mem_csr [35]}),
    .q({open_n15715,data_csr[35]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011110011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3708|ins_dec/reg5_b34  (
    .a({_al_u3430_o,open_n15716}),
    .b({mem_csr_data_max,\ins_dec/op_lui_lutinv }),
    .c({ds1[34],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[34],_al_u7683_o}),
    .sr(\ins_dec/n107 ),
    .f({\exu/alu_au/n53 [34],open_n15729}),
    .q({open_n15733,ds1[34]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3710|_al_u3711  (
    .a({_al_u3709_o,and_clr}),
    .b({mem_csr_data_xor,mem_csr_data_and}),
    .c({ds1[34],ds1[34]}),
    .d({ds2[34],ds2[34]}),
    .f({_al_u3710_o,\exu/alu_au/n47 [34]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3713|exu/reg2_b34  (
    .a({_al_u3710_o,open_n15758}),
    .b({\exu/alu_au/n47 [34],_al_u3713_o}),
    .c({_al_u3712_o,\exu/alu_au/n55 [34]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [34]}),
    .sr(rst_pad),
    .f({_al_u3713_o,\exu/alu_data_mem_csr [34]}),
    .q({open_n15779,data_csr[34]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3716|_al_u3719  (
    .a({_al_u3430_o,and_clr}),
    .b({mem_csr_data_max,mem_csr_data_and}),
    .c({ds1[33],ds1[33]}),
    .d({ds2[33],ds2[33]}),
    .f({\exu/alu_au/n53 [33],\exu/alu_au/n47 [33]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3718|_al_u3722  (
    .a({_al_u3717_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[33],ds1[33]}),
    .d({ds2[33],ds2[33]}),
    .f({_al_u3718_o,\exu/alu_au/n55 [33]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~B*~A*~(D*~C))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0001000000010001),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0001000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3721|exu/reg2_b33  (
    .a({_al_u3718_o,open_n15828}),
    .b({\exu/alu_au/n47 [33],_al_u3721_o}),
    .c({_al_u3720_o,\exu/alu_au/n55 [33]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [33]}),
    .sr(rst_pad),
    .f({_al_u3721_o,\exu/alu_data_mem_csr [33]}),
    .q({open_n15849,data_csr[33]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"))
    \_al_u3724|_al_u3727  (
    .a({_al_u3430_o,and_clr}),
    .b({mem_csr_data_max,mem_csr_data_and}),
    .c({ds1[32],ds1[32]}),
    .d({ds2[32],ds2[32]}),
    .f({\exu/alu_au/n53 [32],\exu/alu_au/n47 [32]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u3726|_al_u3730  (
    .a({_al_u3725_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[32],ds1[32]}),
    .d({ds2[32],ds2[32]}),
    .f({_al_u3726_o,\exu/alu_au/n55 [32]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~B*~A*~(D*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0001000000010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3729|exu/reg2_b32  (
    .a({_al_u3726_o,open_n15890}),
    .b({\exu/alu_au/n47 [32],_al_u3729_o}),
    .c({_al_u3728_o,\exu/alu_au/n55 [32]}),
    .clk(clk_pad),
    .d({mem_csr_data_add,\exu/alu_au/n53 [32]}),
    .sr(rst_pad),
    .f({_al_u3729_o,\exu/alu_data_mem_csr [32]}),
    .q({open_n15907,data_csr[32]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3732|exu/reg2_b31  (
    .a({_al_u3430_o,\exu/alu_au/n53 [31]}),
    .b({mem_csr_data_max,_al_u3735_o}),
    .c({ds1[31],\exu/alu_au/n55 [31]}),
    .clk(clk_pad),
    .d({ds2[31],\exu/alu_au/n47 [31]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [31],\exu/alu_data_mem_csr [31]}),
    .q({open_n15928,data_csr[31]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011110011),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b1100000011110011),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3734|ins_dec/reg5_b31  (
    .a({_al_u3733_o,open_n15929}),
    .b({mem_csr_data_or,\ins_dec/op_lui_lutinv }),
    .c({ds1[31],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({ds2[31],_al_u7571_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3734_o,open_n15946}),
    .q({open_n15950,ds1[31]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3735|_al_u8595  (
    .a({_al_u3734_o,\exu/c_stb_lutinv }),
    .b({mem_csr_data_xor,rd_data_or}),
    .c({ds1[31],ds1[31]}),
    .d({ds2[31],ds2[31]}),
    .f({_al_u3735_o,_al_u8595_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b1100010010000000),
    .MODE("LOGIC"))
    \_al_u3736|_al_u3737  (
    .a({\exu/alu_au/ds1_light_than_ds2_lutinv ,and_clr}),
    .b({mem_csr_data_min,mem_csr_data_and}),
    .c({ds1[31],ds1[31]}),
    .d({ds2[31],ds2[31]}),
    .f({\exu/alu_au/n55 [31],\exu/alu_au/n47 [31]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3739|exu/reg2_b30  (
    .a({_al_u3430_o,\exu/alu_au/n53 [30]}),
    .b({mem_csr_data_max,_al_u3742_o}),
    .c({ds1[30],\exu/alu_au/n55 [30]}),
    .clk(clk_pad),
    .d({ds2[30],\exu/alu_au/n47 [30]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [30],\exu/alu_data_mem_csr [30]}),
    .q({open_n16007,data_csr[30]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3741|_al_u3744  (
    .a({_al_u3740_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[30],ds1[30]}),
    .d({ds2[30],ds2[30]}),
    .f({_al_u3741_o,\exu/alu_au/n47 [30]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3742|_al_u8616  (
    .a({_al_u3741_o,\exu/alu_au/sub_64 [30]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[30],rd_data_sub}),
    .d({ds2[30],ds1[30]}),
    .f({_al_u3742_o,_al_u8616_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3746|exu/reg2_b3  (
    .a({_al_u3430_o,\exu/alu_au/n53 [3]}),
    .b({mem_csr_data_max,_al_u3749_o}),
    .c({ds1[3],\exu/alu_au/n55 [3]}),
    .clk(clk_pad),
    .d({ds2[3],\exu/alu_au/n47 [3]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [3],\exu/alu_data_mem_csr [3]}),
    .q({open_n16072,data_csr[3]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3748|_al_u3751  (
    .a({_al_u3747_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[3],ds1[3]}),
    .d({ds2[3],ds2[3]}),
    .f({_al_u3748_o,\exu/alu_au/n47 [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3749|_al_u9021  (
    .a({_al_u3748_o,\exu/alu_au/sub_64 [3]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[3],rd_data_sub}),
    .d({ds2[3],ds1[3]}),
    .f({_al_u3749_o,_al_u9021_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3753|exu/reg2_b29  (
    .a({_al_u3430_o,\exu/alu_au/n53 [29]}),
    .b({mem_csr_data_max,_al_u3756_o}),
    .c({ds1[29],\exu/alu_au/n55 [29]}),
    .clk(clk_pad),
    .d({ds2[29],\exu/alu_au/n47 [29]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [29],\exu/alu_data_mem_csr [29]}),
    .q({open_n16133,data_csr[29]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3755|_al_u3758  (
    .a({_al_u3754_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[29],ds1[29]}),
    .d({ds2[29],ds2[29]}),
    .f({_al_u3755_o,\exu/alu_au/n47 [29]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3756|_al_u8636  (
    .a({_al_u3755_o,\exu/alu_au/sub_64 [29]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[29],rd_data_sub}),
    .d({ds2[29],ds1[29]}),
    .f({_al_u3756_o,_al_u8636_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3760|exu/reg2_b28  (
    .a({_al_u3430_o,\exu/alu_au/n53 [28]}),
    .b({mem_csr_data_max,_al_u3763_o}),
    .c({ds1[28],\exu/alu_au/n55 [28]}),
    .clk(clk_pad),
    .d({ds2[28],\exu/alu_au/n47 [28]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [28],\exu/alu_data_mem_csr [28]}),
    .q({open_n16198,data_csr[28]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3762|_al_u3765  (
    .a({_al_u3761_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[28],ds1[28]}),
    .d({ds2[28],ds2[28]}),
    .f({_al_u3762_o,\exu/alu_au/n47 [28]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3763|_al_u8656  (
    .a({_al_u3762_o,\exu/alu_au/sub_64 [28]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[28],rd_data_sub}),
    .d({ds2[28],ds1[28]}),
    .f({_al_u3763_o,_al_u8656_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3767|exu/reg2_b27  (
    .a({_al_u3430_o,\exu/alu_au/n53 [27]}),
    .b({mem_csr_data_max,_al_u3770_o}),
    .c({ds1[27],\exu/alu_au/n55 [27]}),
    .clk(clk_pad),
    .d({ds2[27],\exu/alu_au/n47 [27]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [27],\exu/alu_data_mem_csr [27]}),
    .q({open_n16263,data_csr[27]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3769|_al_u3772  (
    .a({_al_u3768_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[27],ds1[27]}),
    .d({ds2[27],ds2[27]}),
    .f({_al_u3769_o,\exu/alu_au/n47 [27]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3770|_al_u8675  (
    .a({_al_u3769_o,\exu/alu_au/sub_64 [27]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[27],rd_data_sub}),
    .d({ds2[27],ds1[27]}),
    .f({_al_u3770_o,_al_u8675_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3774|exu/reg2_b26  (
    .a({_al_u3430_o,\exu/alu_au/n53 [26]}),
    .b({mem_csr_data_max,_al_u3777_o}),
    .c({ds1[26],\exu/alu_au/n55 [26]}),
    .clk(clk_pad),
    .d({ds2[26],\exu/alu_au/n47 [26]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [26],\exu/alu_data_mem_csr [26]}),
    .q({open_n16324,data_csr[26]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3776|_al_u3779  (
    .a({_al_u3775_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[26],ds1[26]}),
    .d({ds2[26],ds2[26]}),
    .f({_al_u3776_o,\exu/alu_au/n47 [26]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3777|_al_u8694  (
    .a({_al_u3776_o,\exu/alu_au/sub_64 [26]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[26],rd_data_sub}),
    .d({ds2[26],ds1[26]}),
    .f({_al_u3777_o,_al_u8694_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3781|exu/reg2_b25  (
    .a({_al_u3430_o,\exu/alu_au/n53 [25]}),
    .b({mem_csr_data_max,_al_u3784_o}),
    .c({ds1[25],\exu/alu_au/n55 [25]}),
    .clk(clk_pad),
    .d({ds2[25],\exu/alu_au/n47 [25]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [25],\exu/alu_data_mem_csr [25]}),
    .q({open_n16385,data_csr[25]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3783|_al_u3786  (
    .a({_al_u3782_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[25],ds1[25]}),
    .d({ds2[25],ds2[25]}),
    .f({_al_u3783_o,\exu/alu_au/n47 [25]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3784|_al_u8712  (
    .a({_al_u3783_o,\exu/alu_au/sub_64 [25]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[25],rd_data_sub}),
    .d({ds2[25],ds1[25]}),
    .f({_al_u3784_o,_al_u8712_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3788|exu/reg2_b24  (
    .a({_al_u3430_o,\exu/alu_au/n53 [24]}),
    .b({mem_csr_data_max,_al_u3791_o}),
    .c({ds1[24],\exu/alu_au/n55 [24]}),
    .clk(clk_pad),
    .d({ds2[24],\exu/alu_au/n47 [24]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [24],\exu/alu_data_mem_csr [24]}),
    .q({open_n16450,data_csr[24]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3790|_al_u3793  (
    .a({_al_u3789_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[24],ds1[24]}),
    .d({ds2[24],ds2[24]}),
    .f({_al_u3790_o,\exu/alu_au/n47 [24]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3791|_al_u8730  (
    .a({_al_u3790_o,\exu/alu_au/sub_64 [24]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[24],rd_data_sub}),
    .d({ds2[24],ds1[24]}),
    .f({_al_u3791_o,_al_u8730_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3795|exu/reg2_b23  (
    .a({_al_u3430_o,\exu/alu_au/n53 [23]}),
    .b({mem_csr_data_max,_al_u3798_o}),
    .c({ds1[23],\exu/alu_au/n55 [23]}),
    .clk(clk_pad),
    .d({ds2[23],\exu/alu_au/n47 [23]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [23],\exu/alu_data_mem_csr [23]}),
    .q({open_n16515,data_csr[23]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3797|_al_u3800  (
    .a({_al_u3796_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[23],ds1[23]}),
    .d({ds2[23],ds2[23]}),
    .f({_al_u3797_o,\exu/alu_au/n47 [23]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3798|_al_u8751  (
    .a({_al_u3797_o,\exu/alu_au/sub_64 [23]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[23],rd_data_sub}),
    .d({ds2[23],ds1[23]}),
    .f({_al_u3798_o,_al_u8751_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3802|exu/reg2_b22  (
    .a({_al_u3430_o,\exu/alu_au/n53 [22]}),
    .b({mem_csr_data_max,_al_u3805_o}),
    .c({ds1[22],\exu/alu_au/n55 [22]}),
    .clk(clk_pad),
    .d({ds2[22],\exu/alu_au/n47 [22]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [22],\exu/alu_data_mem_csr [22]}),
    .q({open_n16576,data_csr[22]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3804|_al_u3807  (
    .a({_al_u3803_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[22],ds1[22]}),
    .d({ds2[22],ds2[22]}),
    .f({_al_u3804_o,\exu/alu_au/n47 [22]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3805|_al_u8770  (
    .a({_al_u3804_o,\exu/alu_au/sub_64 [22]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[22],rd_data_sub}),
    .d({ds2[22],ds1[22]}),
    .f({_al_u3805_o,_al_u8770_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUT1("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT_LUT0(16'b0011111111110101),
    .INIT_LUT1(16'b1100010010000000),
    .MODE("LOGIC"))
    \_al_u3806|_al_u4305  (
    .a({\exu/alu_au/ds1_light_than_ds2_lutinv ,\exu/alu_data_mem_csr [46]}),
    .b({mem_csr_data_min,\exu/alu_data_mem_csr [22]}),
    .c({ds1[22],addr_ex[0]}),
    .d({ds2[22],addr_ex[1]}),
    .f({\exu/alu_au/n55 [22],_al_u4305_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3809|exu/reg2_b21  (
    .a({_al_u3430_o,\exu/alu_au/n53 [21]}),
    .b({mem_csr_data_max,_al_u3812_o}),
    .c({ds1[21],\exu/alu_au/n55 [21]}),
    .clk(clk_pad),
    .d({ds2[21],\exu/alu_au/n47 [21]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [21],\exu/alu_data_mem_csr [21]}),
    .q({open_n16657,data_csr[21]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3811|_al_u3814  (
    .a({_al_u3810_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[21],ds1[21]}),
    .d({ds2[21],ds2[21]}),
    .f({_al_u3811_o,\exu/alu_au/n47 [21]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3812|_al_u8789  (
    .a({_al_u3811_o,\exu/alu_au/sub_64 [21]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[21],rd_data_sub}),
    .d({ds2[21],ds1[21]}),
    .f({_al_u3812_o,_al_u8789_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3816|exu/reg2_b20  (
    .a({_al_u3430_o,\exu/alu_au/n53 [20]}),
    .b({mem_csr_data_max,_al_u3819_o}),
    .c({ds1[20],\exu/alu_au/n55 [20]}),
    .clk(clk_pad),
    .d({ds2[20],\exu/alu_au/n47 [20]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [20],\exu/alu_data_mem_csr [20]}),
    .q({open_n16722,data_csr[20]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3818|_al_u3821  (
    .a({_al_u3817_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[20],ds1[20]}),
    .d({ds2[20],ds2[20]}),
    .f({_al_u3818_o,\exu/alu_au/n47 [20]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3819|_al_u8808  (
    .a({_al_u3818_o,\exu/alu_au/sub_64 [20]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[20],rd_data_sub}),
    .d({ds2[20],ds1[20]}),
    .f({_al_u3819_o,_al_u8808_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3823|exu/reg2_b2  (
    .a({_al_u3430_o,\exu/alu_au/n53 [2]}),
    .b({mem_csr_data_max,_al_u3826_o}),
    .c({ds1[2],\exu/alu_au/n55 [2]}),
    .clk(clk_pad),
    .d({ds2[2],\exu/alu_au/n47 [2]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [2],\exu/alu_data_mem_csr [2]}),
    .q({open_n16787,data_csr[2]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3825|_al_u3828  (
    .a({_al_u3824_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[2],ds1[2]}),
    .d({ds2[2],ds2[2]}),
    .f({_al_u3825_o,\exu/alu_au/n47 [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3826|_al_u9058  (
    .a({_al_u3825_o,\exu/alu_au/sub_64 [2]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[2],rd_data_sub}),
    .d({ds2[2],ds1[2]}),
    .f({_al_u3826_o,_al_u9058_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3830|exu/reg2_b19  (
    .a({_al_u3430_o,\exu/alu_au/n53 [19]}),
    .b({mem_csr_data_max,_al_u3833_o}),
    .c({ds1[19],\exu/alu_au/n55 [19]}),
    .clk(clk_pad),
    .d({ds2[19],\exu/alu_au/n47 [19]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [19],\exu/alu_data_mem_csr [19]}),
    .q({open_n16852,data_csr[19]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3832|_al_u3835  (
    .a({_al_u3831_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[19],ds1[19]}),
    .d({ds2[19],ds2[19]}),
    .f({_al_u3832_o,\exu/alu_au/n47 [19]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3833|_al_u8827  (
    .a({_al_u3832_o,\exu/alu_au/sub_64 [19]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[19],rd_data_sub}),
    .d({ds2[19],ds1[19]}),
    .f({_al_u3833_o,_al_u8827_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3837|exu/reg2_b18  (
    .a({_al_u3430_o,\exu/alu_au/n53 [18]}),
    .b({mem_csr_data_max,_al_u3840_o}),
    .c({ds1[18],\exu/alu_au/n55 [18]}),
    .clk(clk_pad),
    .d({ds2[18],\exu/alu_au/n47 [18]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [18],\exu/alu_data_mem_csr [18]}),
    .q({open_n16913,data_csr[18]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3839|_al_u3842  (
    .a({_al_u3838_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[18],ds1[18]}),
    .d({ds2[18],ds2[18]}),
    .f({_al_u3839_o,\exu/alu_au/n47 [18]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3840|_al_u8846  (
    .a({_al_u3839_o,\exu/alu_au/sub_64 [18]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[18],rd_data_sub}),
    .d({ds2[18],ds1[18]}),
    .f({_al_u3840_o,_al_u8846_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3844|exu/reg2_b17  (
    .a({_al_u3430_o,\exu/alu_au/n53 [17]}),
    .b({mem_csr_data_max,_al_u3847_o}),
    .c({ds1[17],\exu/alu_au/n55 [17]}),
    .clk(clk_pad),
    .d({ds2[17],\exu/alu_au/n47 [17]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [17],\exu/alu_data_mem_csr [17]}),
    .q({open_n16970,data_csr[17]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3846|_al_u3849  (
    .a({_al_u3845_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[17],ds1[17]}),
    .d({ds2[17],ds2[17]}),
    .f({_al_u3846_o,\exu/alu_au/n47 [17]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3847|_al_u8864  (
    .a({_al_u3846_o,\exu/alu_au/sub_64 [17]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[17],rd_data_sub}),
    .d({ds2[17],ds1[17]}),
    .f({_al_u3847_o,_al_u8864_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3851|exu/reg2_b16  (
    .a({_al_u3430_o,\exu/alu_au/n53 [16]}),
    .b({mem_csr_data_max,_al_u3854_o}),
    .c({ds1[16],\exu/alu_au/n55 [16]}),
    .clk(clk_pad),
    .d({ds2[16],\exu/alu_au/n47 [16]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [16],\exu/alu_data_mem_csr [16]}),
    .q({open_n17031,data_csr[16]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3853|_al_u3856  (
    .a({_al_u3852_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[16],ds1[16]}),
    .d({ds2[16],ds2[16]}),
    .f({_al_u3853_o,\exu/alu_au/n47 [16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3854|_al_u8882  (
    .a({_al_u3853_o,\exu/alu_au/sub_64 [16]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[16],rd_data_sub}),
    .d({ds2[16],ds1[16]}),
    .f({_al_u3854_o,_al_u8882_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3858|exu/reg2_b15  (
    .a({_al_u3430_o,\exu/alu_au/n53 [15]}),
    .b({mem_csr_data_max,_al_u3861_o}),
    .c({ds1[15],\exu/alu_au/n55 [15]}),
    .clk(clk_pad),
    .d({ds2[15],\exu/alu_au/n47 [15]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [15],\exu/alu_data_mem_csr [15]}),
    .q({open_n17100,data_csr[15]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3860|_al_u3863  (
    .a({_al_u3859_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[15],ds1[15]}),
    .d({ds2[15],ds2[15]}),
    .f({_al_u3860_o,\exu/alu_au/n47 [15]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3861|_al_u8896  (
    .a({_al_u3860_o,\exu/alu_au/sub_64 [15]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[15],rd_data_sub}),
    .d({ds2[15],ds1[15]}),
    .f({_al_u3861_o,_al_u8896_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3865|exu/reg2_b14  (
    .a({_al_u3430_o,\exu/alu_au/n53 [14]}),
    .b({mem_csr_data_max,_al_u3868_o}),
    .c({ds1[14],\exu/alu_au/n55 [14]}),
    .clk(clk_pad),
    .d({ds2[14],\exu/alu_au/n47 [14]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [14],\exu/alu_data_mem_csr [14]}),
    .q({open_n17161,data_csr[14]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3867|_al_u8932  (
    .a({_al_u3866_o,\exu/alu_au/sub_64 [14]}),
    .b({mem_csr_data_or,rd_data_ds1}),
    .c({ds1[14],rd_data_sub}),
    .d({ds2[14],ds1[14]}),
    .f({_al_u3867_o,_al_u8932_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3868|_al_u3869  (
    .a({_al_u3867_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[14],ds1[14]}),
    .d({ds2[14],ds2[14]}),
    .f({_al_u3868_o,\exu/alu_au/n55 [14]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(C@D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*(C@D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000110011000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000110011000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3871|_al_u3870  (
    .b({open_n17204,ds1[14]}),
    .c({mem_csr_data_and,ds2[14]}),
    .d({\exu/alu_au/alu_and [14],and_clr}),
    .f({\exu/alu_au/n47 [14],\exu/alu_au/alu_and [14]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3873|exu/reg2_b13  (
    .a({_al_u3430_o,\exu/alu_au/n53 [13]}),
    .b({mem_csr_data_max,_al_u3876_o}),
    .c({ds1[13],\exu/alu_au/n55 [13]}),
    .clk(clk_pad),
    .d({ds2[13],\exu/alu_au/n47 [13]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [13],\exu/alu_data_mem_csr [13]}),
    .q({open_n17249,data_csr[13]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3875|_al_u8969  (
    .a({_al_u3874_o,\exu/alu_au/sub_64 [13]}),
    .b({mem_csr_data_or,rd_data_ds1}),
    .c({ds1[13],rd_data_sub}),
    .d({ds2[13],ds1[13]}),
    .f({_al_u3875_o,_al_u8969_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3876|_al_u3877  (
    .a({_al_u3875_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[13],ds1[13]}),
    .d({ds2[13],ds2[13]}),
    .f({_al_u3876_o,\exu/alu_au/n55 [13]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(C@D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*(C@D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000110011000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000110011000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3879|_al_u3878  (
    .b({open_n17300,ds1[13]}),
    .c({mem_csr_data_and,ds2[13]}),
    .d({\exu/alu_au/alu_and [13],and_clr}),
    .f({\exu/alu_au/n47 [13],\exu/alu_au/alu_and [13]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3881|exu/reg2_b12  (
    .a({_al_u3430_o,\exu/alu_au/n53 [12]}),
    .b({mem_csr_data_max,_al_u3884_o}),
    .c({ds1[12],\exu/alu_au/n55 [12]}),
    .clk(clk_pad),
    .d({ds2[12],\exu/alu_au/n47 [12]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [12],\exu/alu_data_mem_csr [12]}),
    .q({open_n17345,data_csr[12]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*~(~D*~C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*~(~D*~C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3883|_al_u9004  (
    .a({_al_u3882_o,\exu/alu_au/sub_64 [12]}),
    .b({mem_csr_data_or,rd_data_ds1}),
    .c({ds1[12],rd_data_sub}),
    .d({ds2[12],ds1[12]}),
    .f({_al_u3883_o,_al_u9004_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3884|_al_u3885  (
    .a({_al_u3883_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[12],ds1[12]}),
    .d({ds2[12],ds2[12]}),
    .f({_al_u3884_o,\exu/alu_au/n55 [12]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(C@D))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000110011000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3887|_al_u3886  (
    .b({open_n17396,ds1[12]}),
    .c({mem_csr_data_and,ds2[12]}),
    .d({\exu/alu_au/alu_and [12],and_clr}),
    .f({\exu/alu_au/n47 [12],\exu/alu_au/alu_and [12]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3889|exu/reg2_b11  (
    .a({_al_u3430_o,\exu/alu_au/n53 [11]}),
    .b({mem_csr_data_max,_al_u3892_o}),
    .c({ds1[11],\exu/alu_au/n55 [11]}),
    .clk(clk_pad),
    .d({ds2[11],\exu/alu_au/n47 [11]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [11],\exu/alu_data_mem_csr [11]}),
    .q({open_n17433,data_csr[11]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3891|_al_u9039  (
    .a({_al_u3890_o,\exu/alu_au/sub_64 [11]}),
    .b({mem_csr_data_or,rd_data_ds1}),
    .c({ds1[11],rd_data_sub}),
    .d({ds2[11],ds1[11]}),
    .f({_al_u3891_o,_al_u9039_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3892|_al_u3893  (
    .a({_al_u3891_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[11],ds1[11]}),
    .d({ds2[11],ds2[11]}),
    .f({_al_u3892_o,\exu/alu_au/n55 [11]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(C@D))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000110011000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u3895|_al_u3894  (
    .b({open_n17476,ds1[11]}),
    .c({mem_csr_data_and,ds2[11]}),
    .d({\exu/alu_au/alu_and [11],and_clr}),
    .f({\exu/alu_au/n47 [11],\exu/alu_au/alu_and [11]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~C*B*~A)"),
    //.LUTF1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(~D*~C*B*~A)"),
    //.LUTG1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111011),
    .INIT_LUTF1(16'b1100100001000000),
    .INIT_LUTG0(16'b1111111111111011),
    .INIT_LUTG1(16'b1100100001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3897|exu/reg2_b10  (
    .a({_al_u3430_o,\exu/alu_au/n53 [10]}),
    .b({mem_csr_data_max,_al_u3900_o}),
    .c({ds1[10],\exu/alu_au/n55 [10]}),
    .clk(clk_pad),
    .d({ds2[10],\exu/alu_au/n47 [10]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [10],\exu/alu_data_mem_csr [10]}),
    .q({open_n17517,data_csr[10]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3899|_al_u9076  (
    .a({_al_u3898_o,\exu/alu_au/sub_64 [10]}),
    .b({mem_csr_data_or,rd_data_ds1}),
    .c({ds1[10],rd_data_sub}),
    .d({ds2[10],ds1[10]}),
    .f({_al_u3899_o,_al_u9076_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u3900|_al_u3901  (
    .a({_al_u3899_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[10],ds1[10]}),
    .d({ds2[10],ds2[10]}),
    .f({_al_u3900_o,\exu/alu_au/n55 [10]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(C@D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*(C@D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000110011000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000110011000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3903|_al_u3902  (
    .b({open_n17560,ds1[10]}),
    .c({mem_csr_data_and,ds2[10]}),
    .d({\exu/alu_au/alu_and [10],and_clr}),
    .f({\exu/alu_au/n47 [10],\exu/alu_au/alu_and [10]}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3905|exu/reg2_b1  (
    .a({_al_u3430_o,\exu/alu_au/n53 [1]}),
    .b({mem_csr_data_max,_al_u3908_o}),
    .c({ds1[1],\exu/alu_au/n55 [1]}),
    .clk(clk_pad),
    .d({ds2[1],\exu/alu_au/n47 [1]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [1],\exu/alu_data_mem_csr [1]}),
    .q({open_n17601,data_csr[1]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3907|_al_u3910  (
    .a({_al_u3906_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[1],ds1[1]}),
    .d({ds2[1],ds2[1]}),
    .f({_al_u3907_o,\exu/alu_au/n47 [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3908|_al_u9094  (
    .a({_al_u3907_o,\exu/alu_au/sub_64 [1]}),
    .b({mem_csr_data_xor,rd_data_ds1}),
    .c({ds1[1],rd_data_sub}),
    .d({ds2[1],ds1[1]}),
    .f({_al_u3908_o,_al_u9094_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*B*~A)"),
    //.LUT1("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111011),
    .INIT_LUT1(16'b1100100001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3912|exu/reg2_b0  (
    .a({_al_u3430_o,\exu/alu_au/n53 [0]}),
    .b({mem_csr_data_max,_al_u3915_o}),
    .c({ds1[0],\exu/alu_au/n55 [0]}),
    .clk(clk_pad),
    .d({ds2[0],\exu/alu_au/n47 [0]}),
    .sr(rst_pad),
    .f({\exu/alu_au/n53 [0],\exu/alu_data_mem_csr [0]}),
    .q({open_n17662,data_csr[0]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*C)*~(B*A))"),
    //.LUT1("(~(D*C)*~(B*A))"),
    .INIT_LUT0(16'b0000011101110111),
    .INIT_LUT1(16'b0000011101110111),
    .MODE("LOGIC"))
    \_al_u3913|_al_u9112  (
    .a({\exu/alu_au/add_64 [0],\exu/alu_au/add_64 [0]}),
    .b({mem_csr_data_add,rd_data_add}),
    .c({mem_csr_data_ds2,rd_data_ds1}),
    .d({ds2[0],ds1[0]}),
    .f({_al_u3913_o,_al_u9112_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(A*~(B*~(~D*~C)))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0010001000101010),
    .MODE("LOGIC"))
    \_al_u3914|_al_u3917  (
    .a({_al_u3913_o,and_clr}),
    .b({mem_csr_data_or,mem_csr_data_and}),
    .c({ds1[0],ds1[0]}),
    .d({ds2[0],ds2[0]}),
    .f({_al_u3914_o,\exu/alu_au/n47 [0]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3915|_al_u3916  (
    .a({_al_u3914_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({mem_csr_data_xor,mem_csr_data_min}),
    .c({ds1[0],ds1[0]}),
    .d({ds2[0],ds2[0]}),
    .f({_al_u3915_o,\exu/alu_au/n55 [0]}));
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~B*~(~C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3919|ins_dec/reg10_b14  (
    .b({\ins_dec/op_load ,open_n17729}),
    .c({_al_u3216_o,_al_u3216_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/op_store ,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3919_o,open_n17746}),
    .q({open_n17750,ex_exc_code[14]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3922|_al_u3391  (
    .b({open_n17753,\ins_dec/funct3_0_lutinv }),
    .c({id_ins[25],id_system}),
    .d({\ins_dec/funct6_0_lutinv ,\ins_dec/funct6_0_lutinv }),
    .f({\ins_dec/funct7_0_lutinv ,_al_u3391_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(~B*~A*~(~D*~C))"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(~B*~A*~(~D*~C))"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0001000100010000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0001000100010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3923|_al_u3954  (
    .a({_al_u2929_o,_al_u2938_o}),
    .b({_al_u2930_o,_al_u2939_o}),
    .c({_al_u2931_o,_al_u2944_o}),
    .d({_al_u2932_o,_al_u3923_o}),
    .f({_al_u3923_o,\ins_dec/op_lui_lutinv }));
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3924|ins_dec/reg10_b4  (
    .c({_al_u2930_o,_al_u3924_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u2929_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3924_o,open_n17818}),
    .q({open_n17822,ex_exc_code[4]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(D*~C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3925|ins_dec/store_reg  (
    .a({_al_u3924_o,_al_u2933_o}),
    .b({_al_u2938_o,_al_u2938_o}),
    .c({_al_u2939_o,_al_u2939_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u2944_o,_al_u2944_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3925_o,\ins_dec/op_store }),
    .q({open_n17838,store}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3926|_al_u7141  (
    .b({_al_u3923_o,_al_u3925_o}),
    .c({_al_u3925_o,_al_u4064_o}),
    .d({\ins_dec/funct7_0_lutinv ,_al_u3927_o}),
    .f({_al_u3926_o,_al_u7141_o}));
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(D*~C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3927|ins_dec/load_reg  (
    .a({_al_u3924_o,_al_u2933_o}),
    .b({_al_u2938_o,_al_u2938_o}),
    .c({_al_u2939_o,_al_u2939_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u2946_o,_al_u2946_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3927_o,\ins_dec/op_load }),
    .q({open_n17884,load}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3929|ins_dec/reg10_b3  (
    .b({_al_u3927_o,open_n17887}),
    .c({_al_u3928_o,_al_u3928_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3926_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3929_o,open_n17904}),
    .q({open_n17908,ex_exc_code[3]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*C*B*~A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*C*B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3932|ins_dec/reg10_b31  (
    .a({id_ins[31],open_n17909}),
    .b({id_ins[30],open_n17910}),
    .c({id_ins[28],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[26],id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3932_o,open_n17927}),
    .q({open_n17931,ex_exc_code[31]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("(D*C*~B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b0010000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3933|ins_dec/reg8_b16  (
    .a({_al_u3932_o,open_n17932}),
    .b({id_ins[29],_al_u3214_o}),
    .c({id_ins[27],id_ins[27]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[25],_al_u4055_o}),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/funct7_32_lutinv ,open_n17945}),
    .q({open_n17949,as2[16]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3937|_al_u3936  (
    .b({\ins_dec/funct3_0_lutinv ,open_n17952}),
    .c({\ins_dec/op_32_reg_lutinv ,_al_u3928_o}),
    .d({\ins_dec/funct7_0_lutinv ,_al_u3925_o}),
    .f({\ins_dec/ins_addw ,\ins_dec/op_32_reg_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("(C*~B*D)"),
    .INIT_LUT0(16'b1111001111000000),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"))
    \_al_u3938|_al_u3217  (
    .b({_al_u3216_o,1'b0}),
    .c({_al_u3217_o,\ins_fetch/ins_hold [13]}),
    .d({\ins_dec/op_amo ,\ins_fetch/ins_shift [13]}),
    .f({_al_u3938_o,_al_u3217_o}));
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3939|ins_dec/reg10_b28  (
    .b({id_ins[28],open_n18001}),
    .c({id_ins[27],id_ins[28]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3938_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3939_o,open_n18018}),
    .q({open_n18022,ex_exc_code[28]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~B*A)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(~D*C*~B*A)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3944|_al_u4834  (
    .a({open_n18023,_al_u2847_o}),
    .b(\biu/cache_ctrl_logic/statu [3:2]),
    .c(\biu/cache_ctrl_logic/statu [4:3]),
    .d({\biu/cache_ctrl_logic/statu [2],\biu/cache_ctrl_logic/statu [4]}),
    .f({_al_u3944_o,_al_u4834_o}));
  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3955|ins_dec/id_system_reg  (
    .a({_al_u2938_o,_al_u2938_o}),
    .b({_al_u2939_o,_al_u2939_o}),
    .c({_al_u2946_o,_al_u2946_o}),
    .ce(\ins_dec/u461_sel_is_0_o ),
    .clk(clk_pad),
    .d({_al_u3923_o,_al_u2948_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3955_o,id_system}),
    .q({open_n18063,ex_system}));  // ../../RTL/CPU/ID/ins_dec.v(830)
  // ../../RTL/CPU/ID/ins_dec.v(674)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3956|ins_dec/jmp_reg  (
    .a({_al_u3213_o,open_n18064}),
    .b({_al_u3214_o,open_n18065}),
    .c({\ins_dec/op_lui_lutinv ,_al_u3214_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3955_o,_al_u3213_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3956_o,\ins_dec/n59 }),
    .q({open_n18081,jmp}));  // ../../RTL/CPU/ID/ins_dec.v(674)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3957|ins_fetch/reg1_b19  (
    .b({1'b0,ins_read[51]}),
    .c({\ins_fetch/ins_hold [19],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({\ins_fetch/ins_shift [19],ins_read[19]}),
    .sr(rst_pad),
    .f({id_ins[19],\ins_fetch/ins_shift [19]}),
    .q({open_n18103,\ins_fetch/ins_hold [19]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3958|ins_dec/reg10_b19  (
    .c({id_ins[19],id_ins[19]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3956_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({id_rs1_index[4],open_n18120}),
    .q({open_n18124,ex_exc_code[19]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1111001111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3959|ins_fetch/reg1_b18  (
    .b({1'b0,ins_read[50]}),
    .c({\ins_fetch/ins_hold [18],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({\ins_fetch/ins_shift [18],ins_read[18]}),
    .sr(rst_pad),
    .f({id_ins[18],\ins_fetch/ins_shift [18]}),
    .q({open_n18142,\ins_fetch/ins_hold [18]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3960|ins_dec/reg10_b18  (
    .c({id_ins[18],id_ins[18]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3956_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({id_rs1_index[3],open_n18159}),
    .q({open_n18163,ex_exc_code[18]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1111001111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3961|ins_fetch/reg1_b17  (
    .b({1'b0,ins_read[49]}),
    .c({\ins_fetch/ins_hold [17],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({\ins_fetch/ins_shift [17],ins_read[17]}),
    .sr(rst_pad),
    .f({id_ins[17],\ins_fetch/ins_shift [17]}),
    .q({open_n18181,\ins_fetch/ins_hold [17]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3962|ins_dec/reg10_b17  (
    .c({id_ins[17],id_ins[17]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3956_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({id_rs1_index[2],open_n18198}),
    .q({open_n18202,ex_exc_code[17]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3963|ins_fetch/reg1_b16  (
    .b({1'b0,ins_read[48]}),
    .c({\ins_fetch/ins_hold [16],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({\ins_fetch/ins_shift [16],ins_read[16]}),
    .sr(rst_pad),
    .f({id_ins[16],\ins_fetch/ins_shift [16]}),
    .q({open_n18224,\ins_fetch/ins_hold [16]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3964|ins_dec/reg10_b16  (
    .c({id_ins[16],id_ins[16]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3956_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({id_rs1_index[1],open_n18241}),
    .q({open_n18245,ex_exc_code[16]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3966|ins_dec/reg10_b15  (
    .c({id_ins[15],id_ins[15]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3956_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({id_rs1_index[0],open_n18266}),
    .q({open_n18270,ex_exc_code[15]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u3967|_al_u7142  (
    .c({\ins_dec/op_load ,id_system}),
    .d({\ins_dec/op_store ,\ins_dec/op_load }),
    .f({\ins_dec/mux24_b10_sel_is_0_o ,_al_u7142_o}));
  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(D*C*~B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3969|ins_dec/mem_csr_data_min_reg  (
    .a({_al_u3939_o,open_n18295}),
    .b({id_ins[31],id_ins[31]}),
    .c(id_ins[30:29]),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[29],_al_u3939_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3969_o,open_n18312}),
    .q({open_n18316,mem_csr_data_min}));  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b1111001111000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u3971|_al_u3384  (
    .b({_al_u3217_o,1'b0}),
    .c({_al_u3384_o,\ins_fetch/ins_hold [12]}),
    .d({id_system,\ins_fetch/ins_shift [12]}),
    .f({\ins_dec/n149_lutinv ,_al_u3384_o}));
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3972|ins_dec/reg10_b30  (
    .b({id_ins[30],open_n18341}),
    .c({id_ins[29],id_ins[30]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[31],id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u3972_o,open_n18358}),
    .q({open_n18362,ex_exc_code[30]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*~B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u3973|ins_dec/reg10_b27  (
    .b({id_ins[28],open_n18365}),
    .c({id_ins[27],id_ins[27]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3972_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/funct5_8_lutinv ,open_n18378}),
    .q({open_n18382,ex_exc_code[27]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4039|_al_u7983  (
    .c({\exu/lsu/n0_lutinv ,unsign}),
    .d({\exu/alu_data_mem_csr [7],\exu/lsu/n0_lutinv }),
    .f({\exu/lsu/n1 [7],\exu/lsu/mux27_b56_sel_is_3_o }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u4040|_al_u3943  (
    .b({uncache_data[7],open_n18413}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[7]}),
    .d({\exu/lsu/n1 [7],_al_u2705_o}),
    .f({\biu/l1i_in [7],uncache_data[7]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4041|_al_u4223  (
    .b({open_n18436,\exu/alu_data_mem_csr [19]}),
    .c({\exu/lsu/n0_lutinv ,\exu/lsu/n0_lutinv }),
    .d({\exu/alu_data_mem_csr [6],_al_u4222_o}),
    .f({\exu/lsu/n1 [6],_al_u4223_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0011111111110101),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0011111111110101),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4042|_al_u8910  (
    .a({open_n18457,uncache_data[6]}),
    .b({uncache_data[6],uncache_data[30]}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,addr_ex[0]}),
    .d({\exu/lsu/n1 [6],addr_ex[1]}),
    .f({\biu/l1i_in [6],_al_u8910_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4043|_al_u4211  (
    .b({open_n18484,\exu/alu_data_mem_csr [23]}),
    .c({\exu/lsu/n0_lutinv ,\exu/lsu/n0_lutinv }),
    .d({\exu/alu_data_mem_csr [5],_al_u4210_o}),
    .f({\exu/lsu/n1 [5],_al_u4211_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4044|biu/cache_ctrl_logic/reg7_b5  (
    .b({uncache_data[5],open_n18507}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[5]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n1 [5],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [5],uncache_data[5]}),
    .q({open_n18527,\biu/cache_ctrl_logic/pte_temp [5]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4045|_al_u7989  (
    .c({\exu/lsu/n0_lutinv ,\exu/lsu/n0_lutinv }),
    .d({\exu/alu_data_mem_csr [4],uncache_data[15]}),
    .f({\exu/lsu/n1 [4],\exu/lsu/n22 [15]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4046|biu/cache_ctrl_logic/reg7_b4  (
    .b({uncache_data[4],open_n18554}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[4]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n1 [4],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [4],uncache_data[4]}),
    .q({open_n18570,\biu/cache_ctrl_logic/pte_temp [4]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4047|_al_u4051  (
    .c({\exu/lsu/n0_lutinv ,\exu/lsu/n0_lutinv }),
    .d({\exu/alu_data_mem_csr [3],\exu/alu_data_mem_csr [1]}),
    .f({\exu/lsu/n1 [3],\exu/lsu/n1 [1]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4048|biu/cache_ctrl_logic/reg7_b3  (
    .b({uncache_data[3],open_n18601}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[3]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n1 [3],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [3],uncache_data[3]}),
    .q({open_n18617,\biu/cache_ctrl_logic/pte_temp [3]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4050|biu/cache_ctrl_logic/reg7_b2  (
    .b({uncache_data[2],open_n18620}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[2]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n1 [2],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [2],uncache_data[2]}),
    .q({open_n18640,\biu/cache_ctrl_logic/pte_temp [2]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4052|biu/cache_ctrl_logic/reg7_b1  (
    .b({uncache_data[1],open_n18643}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[1]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n1 [1],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [1],uncache_data[1]}),
    .q({open_n18663,\biu/cache_ctrl_logic/pte_temp [1]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000110000001010),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000110000001010),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4053|_al_u4207  (
    .a({open_n18664,\exu/alu_data_mem_csr [16]}),
    .b({open_n18665,\exu/alu_data_mem_csr [0]}),
    .c({\exu/lsu/n0_lutinv ,addr_ex[0]}),
    .d({\exu/alu_data_mem_csr [0],addr_ex[1]}),
    .f({\exu/lsu/n1 [0],_al_u4207_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4054|biu/cache_ctrl_logic/reg7_b0  (
    .b({uncache_data[0],hrdata_pad[0]}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,\biu/bus_unit/mmu_hwdata [0]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n1 [0],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [0],uncache_data[0]}),
    .q({open_n18711,\biu/cache_ctrl_logic/pte_temp [0]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("(C*~(~B*D))"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("(C*~(~B*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b1100000011110000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b1100000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4055|ins_dec/reg8_b20  (
    .b({_al_u3382_o,\ins_dec/mux24_b10_sel_is_0_o }),
    .c({id_ins[31],id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/mux24_b10_sel_is_0_o ,\ins_dec/n302 }),
    .sr(\ins_dec/n107 ),
    .f({_al_u4055_o,open_n18730}),
    .q({open_n18734,as2[20]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(D*~C*B*A)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"))
    \_al_u4064|_al_u2941  (
    .a({_al_u2933_o,open_n18735}),
    .b({_al_u2938_o,open_n18736}),
    .c({_al_u2939_o,\ins_fetch/ins_hold [6]}),
    .d({_al_u3212_o,1'b0}),
    .f({_al_u4064_o,_al_u2941_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4065|_al_u4875  (
    .c({_al_u4064_o,_al_u4064_o}),
    .d({_al_u3213_o,_al_u3214_o}),
    .f({\ins_dec/mux27_b12_sel_is_0_o ,_al_u4875_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4066|ins_dec/reg8_b4  (
    .b({_al_u3214_o,open_n18787}),
    .c({id_ins[15],_al_u4069_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/mux27_b12_sel_is_0_o ,_al_u4067_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4066_o,open_n18804}),
    .q({open_n18808,as2[4]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(B*~(~A*~(~D*C)))"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(B*~(~A*~(~D*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1000100011001000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1000100011001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4067|ins_dec/reg4_b4  (
    .a({\ins_dec/mux24_b10_sel_is_0_o ,open_n18809}),
    .b({_al_u4066_o,1'b0}),
    .c({\ins_dec/op_store ,\ins_fetch/ins_hold [11]}),
    .ce(\ins_dec/mux13_b0_sel_is_0_o ),
    .clk(clk_pad),
    .d({id_ins[11],\ins_fetch/ins_shift [11]}),
    .f({_al_u4067_o,id_ins[11]}),
    .q({open_n18830,ex_rd_index[4]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4068|ins_dec/reg8_b56  (
    .b({_al_u3214_o,open_n18833}),
    .c({_al_u4064_o,id_ins[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/op_store ,\ins_dec/mux27_b56_sel_is_0_o }),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/mux27_b56_sel_is_0_o ,open_n18846}),
    .q({open_n18850,as2[56]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111000000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4069|ins_dec/reg4_b3  (
    .a({\ins_dec/mux27_b56_sel_is_0_o ,open_n18851}),
    .b({_al_u4064_o,1'b0}),
    .c({id_ins[24],\ins_fetch/ins_hold [10]}),
    .ce(\ins_dec/mux13_b0_sel_is_0_o ),
    .clk(clk_pad),
    .d({id_ins[10],\ins_fetch/ins_shift [10]}),
    .f({_al_u4069_o,id_ins[10]}),
    .q({open_n18868,ex_rd_index[3]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4071|_al_u3216  (
    .b({_al_u3214_o,1'b0}),
    .c({_al_u3216_o,\ins_fetch/ins_hold [14]}),
    .d({\ins_dec/mux27_b12_sel_is_0_o ,\ins_fetch/ins_shift [14]}),
    .f({_al_u4071_o,_al_u3216_o}));
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~(~A*~(~D*C)))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~(~A*~(~D*C)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000100011001000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000100011001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4072|ins_dec/reg10_b10  (
    .a({\ins_dec/mux24_b10_sel_is_0_o ,open_n18895}),
    .b({_al_u4071_o,open_n18896}),
    .c({\ins_dec/op_store ,id_ins[10]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[10],id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4072_o,open_n18913}),
    .q({open_n18917,ex_exc_code[10]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4073|ins_dec/reg4_b2  (
    .a({\ins_dec/mux27_b56_sel_is_0_o ,open_n18918}),
    .b({_al_u4064_o,1'b0}),
    .c({id_ins[9],\ins_fetch/ins_hold [9]}),
    .ce(\ins_dec/mux13_b0_sel_is_0_o ),
    .clk(clk_pad),
    .d({id_ins[23],\ins_fetch/ins_shift [9]}),
    .f({_al_u4073_o,id_ins[9]}),
    .q({open_n18939,ex_rd_index[2]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4075|_al_u4079  (
    .b({_al_u3214_o,_al_u3214_o}),
    .c({_al_u3217_o,_al_u3384_o}),
    .d({\ins_dec/mux27_b12_sel_is_0_o ,\ins_dec/mux27_b12_sel_is_0_o }),
    .f({_al_u4075_o,_al_u4079_o}));
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*~(~A*~(~D*C)))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*~(~A*~(~D*C)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000100011001000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000100011001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4076|ins_dec/reg10_b9  (
    .a({\ins_dec/mux24_b10_sel_is_0_o ,open_n18966}),
    .b({_al_u4075_o,open_n18967}),
    .c({\ins_dec/op_store ,id_ins[9]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[9],id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4076_o,open_n18984}),
    .q({open_n18988,ex_exc_code[9]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111000000),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4077|ins_dec/reg4_b1  (
    .a({\ins_dec/mux27_b56_sel_is_0_o ,open_n18989}),
    .b({_al_u4064_o,1'b0}),
    .c({id_ins[8],\ins_fetch/ins_hold [8]}),
    .ce(\ins_dec/mux13_b0_sel_is_0_o ),
    .clk(clk_pad),
    .d({id_ins[22],\ins_fetch/ins_shift [8]}),
    .f({_al_u4077_o,id_ins[8]}),
    .q({open_n19006,ex_rd_index[1]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~(~A*~(~D*C)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000100011001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4080|ins_dec/reg10_b8  (
    .a({\ins_dec/mux24_b10_sel_is_0_o ,open_n19007}),
    .b({_al_u4079_o,open_n19008}),
    .c({\ins_dec/op_store ,id_ins[8]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[8],id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4080_o,open_n19021}),
    .q({open_n19025,ex_exc_code[8]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u4081|ins_dec/reg4_b0  (
    .a({\ins_dec/mux27_b56_sel_is_0_o ,open_n19026}),
    .b({_al_u4064_o,1'b0}),
    .c({id_ins[7],\ins_fetch/ins_hold [7]}),
    .ce(\ins_dec/mux13_b0_sel_is_0_o ),
    .clk(clk_pad),
    .d({id_ins[21],\ins_fetch/ins_shift [7]}),
    .f({_al_u4081_o,id_ins[7]}),
    .q({open_n19047,ex_rd_index[0]}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4083|ins_dec/reg10_b7  (
    .c({id_ins[7],id_ins[7]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/op_store ,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4083_o,open_n19064}),
    .q({open_n19068,ex_exc_code[7]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("~(~D*~(C*~B))"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100110000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111111100110000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4084|ins_dec/reg8_b0  (
    .b({open_n19071,_al_u4084_o}),
    .c({_al_u3213_o,id_ins[20]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/op_load ,_al_u4083_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4084_o,open_n19088}),
    .q({open_n19092,as2[0]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4086|ins_dec/gpr_write_reg  (
    .a({\ins_dec/op_store ,open_n19093}),
    .b({\ins_dec/op_amo ,\ins_dec/op_store }),
    .c({_al_u3925_o,_al_u4064_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4064_o,\ins_dec/ins_fence }),
    .sr(\ins_dec/n107 ),
    .f({_al_u4086_o,open_n19110}),
    .q({open_n19114,ex_gpr_write}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4087|ins_dec/reg10_b24  (
    .c({id_ins[24],id_ins[24]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4086_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({id_rs2_index[4],open_n19135}),
    .q({open_n19139,ex_exc_code[24]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4088|ins_dec/reg10_b23  (
    .c({id_ins[23],id_ins[23]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4086_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({id_rs2_index[3],open_n19160}),
    .q({open_n19164,ex_exc_code[23]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4089|ins_dec/reg10_b22  (
    .c({id_ins[22],id_ins[22]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4086_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({id_rs2_index[2],open_n19181}),
    .q({open_n19185,ex_exc_code[22]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4090|ins_dec/reg10_b21  (
    .c({id_ins[21],id_ins[21]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4086_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({id_rs2_index[1],open_n19206}),
    .q({open_n19210,ex_exc_code[21]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u4091|_al_u6211  (
    .b({open_n19213,_al_u3927_o}),
    .c({id_ins[20],id_ins[20]}),
    .d({_al_u4086_o,_al_u4086_o}),
    .f({id_rs2_index[0],_al_u6211_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4092|_al_u6065  (
    .b({_al_u3927_o,open_n19236}),
    .c({_al_u3928_o,id_ins[31]}),
    .d({\ins_dec/funct6_0_lutinv ,_al_u3927_o}),
    .f({_al_u4092_o,_al_u6065_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4093|_al_u4094  (
    .b({\ins_dec/n35_lutinv ,\ins_dec/n35_lutinv }),
    .c({_al_u3384_o,_al_u3384_o}),
    .d({_al_u4092_o,\ins_dec/funct7_0_lutinv }),
    .f({\ins_dec/ins_slli ,_al_u4094_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4095|_al_u4805  (
    .a({open_n19287,\ins_dec/funct5_8_lutinv }),
    .b({open_n19288,_al_u3927_o}),
    .c({_al_u3928_o,_al_u4804_o}),
    .d({_al_u3927_o,_al_u3928_o}),
    .f({\ins_dec/op_32_imm_lutinv ,\ins_dec/ins_srai }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4099|_al_u7495  (
    .b({open_n19315,hready_pad}),
    .c({hresp_pad,hresp_pad}),
    .d({hready_pad,_al_u2964_o}),
    .f({_al_u4099_o,_al_u7495_o}));
  // ../../RTL/CPU/BIU/bus_unit.v(163)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)"),
    //.LUTG0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b1100110000001111),
    .INIT_LUTG0(16'b0011001100001111),
    .INIT_LUTG1(16'b1100110000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4101|biu/bus_unit/reg1_b3  (
    .b({_al_u4100_o,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .c({hresp_pad,_al_u4101_o}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mux10_b3_sel_is_0_o ,_al_u2833_o}),
    .sr(rst_pad),
    .f({_al_u4101_o,open_n19359}),
    .q({open_n19363,\biu/bus_unit/statu [3]}));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000000011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4103|cu_ru/medeleg_exc_ctrl/dspf_reg  (
    .a({open_n19364,\cu_ru/read_mcycle_sel_lutinv }),
    .b({\cu_ru/medeleg [15],\cu_ru/read_medeleg_sel_lutinv }),
    .c({wb_st_page_fault,\cu_ru/mcycle [15]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n5 [1],\cu_ru/medeleg [15]}),
    .mi({open_n19375,data_csr[15]}),
    .sr(rst_pad),
    .f({\cu_ru/medeleg_exc_ctrl/spf_target_s ,_al_u7266_o}),
    .q({open_n19379,\cu_ru/medeleg [15]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4105|_al_u4104  (
    .b({open_n19382,\cu_ru/medeleg [15]}),
    .c({\cu_ru/medeleg_exc_ctrl/spf_target_m_lutinv ,wb_st_page_fault}),
    .d({\cu_ru/medeleg_exc_ctrl/spf_target_s ,priv[3]}),
    .f({\cu_ru/medeleg_exc_ctrl/n85_neg_lutinv ,\cu_ru/medeleg_exc_ctrl/spf_target_m_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(D*~(C*~B*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(D*~(C*~B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b1101111100000000),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b1101111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4106|cu_ru/medeleg_exc_ctrl/dlpf_reg  (
    .a({\cu_ru/m_s_status/n5 [1],open_n19403}),
    .b({priv[3],\cu_ru/stval [13]}),
    .c({\cu_ru/medeleg [13],data_csr[13]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({wb_ld_page_fault,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n19407,data_csr[13]}),
    .sr(rst_pad),
    .f({_al_u4106_o,_al_u5335_o}),
    .q({open_n19422,\cu_ru/medeleg [13]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4107|_al_u4116  (
    .c({_al_u4106_o,\cu_ru/medeleg_exc_ctrl/iam_target_m_lutinv }),
    .d({\cu_ru/medeleg_exc_ctrl/n85_neg_lutinv ,\cu_ru/medeleg_exc_ctrl/iam_target_s }),
    .f({_al_u4107_o,\cu_ru/medeleg_exc_ctrl/n80_neg_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4108|cu_ru/medeleg_exc_ctrl/dsaf_reg  (
    .a({open_n19451,\cu_ru/read_scause_sel_lutinv }),
    .b({open_n19452,\cu_ru/read_medeleg_sel_lutinv }),
    .c({wb_st_acc_fault,\cu_ru/scause [7]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/medeleg [7],\cu_ru/medeleg [7]}),
    .mi({open_n19456,data_csr[7]}),
    .sr(rst_pad),
    .f({_al_u4108_o,_al_u7502_o}),
    .q({open_n19471,\cu_ru/medeleg [7]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("(~C*~(B*~D))"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("(~C*~(B*~D))"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000111100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4110|_al_u4109  (
    .b({_al_u4108_o,\cu_ru/medeleg [7]}),
    .c({\cu_ru/medeleg_exc_ctrl/saf_target_m_lutinv ,wb_st_acc_fault}),
    .d({\cu_ru/m_s_status/n5 [1],priv[3]}),
    .f({\cu_ru/medeleg_exc_ctrl/n87_neg_lutinv ,\cu_ru/medeleg_exc_ctrl/saf_target_m_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000000011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4111|cu_ru/medeleg_exc_ctrl/dlaf_reg  (
    .a({open_n19498,\cu_ru/read_medeleg_sel_lutinv }),
    .b({\cu_ru/medeleg [5],\cu_ru/read_satp_sel_lutinv }),
    .c({wb_ld_acc_fault,satp[5]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n5 [1],\cu_ru/medeleg [5]}),
    .mi({open_n19509,data_csr[5]}),
    .sr(rst_pad),
    .f({\cu_ru/medeleg_exc_ctrl/laf_target_s ,_al_u7879_o}),
    .q({open_n19513,\cu_ru/medeleg [5]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4113|_al_u4112  (
    .a({_al_u4107_o,open_n19514}),
    .b({\cu_ru/medeleg_exc_ctrl/n87_neg_lutinv ,\cu_ru/medeleg [5]}),
    .c({\cu_ru/medeleg_exc_ctrl/laf_target_s ,wb_ld_acc_fault}),
    .d({\cu_ru/medeleg_exc_ctrl/laf_target_m_lutinv ,priv[3]}),
    .f({_al_u4113_o,\cu_ru/medeleg_exc_ctrl/laf_target_m_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4114|cu_ru/medeleg_exc_ctrl/diam_reg  (
    .b({\cu_ru/medeleg [0],\cu_ru/mepc [0]}),
    .c({wb_ins_addr_mis,data_csr[0]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n5 [1],\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .mi({open_n19544,data_csr[0]}),
    .sr(rst_pad),
    .f({\cu_ru/medeleg_exc_ctrl/iam_target_s ,_al_u6696_o}),
    .q({open_n19559,\cu_ru/medeleg [0]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(D*~(C*~B*A))"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b1101111100000000),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b1101111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4117|exu/ill_ins_reg  (
    .a({\cu_ru/m_s_status/n5 [1],ex_ill_ins}),
    .b({priv[3],ex_ins_acc_fault}),
    .c({\cu_ru/medeleg [2],ex_ins_addr_mis}),
    .clk(clk_pad),
    .d({wb_ill_ins,ex_ins_page_fault}),
    .mi({open_n19564,ex_ill_ins}),
    .sr(\exu/n86 ),
    .f({_al_u4117_o,\exu/n17_lutinv }),
    .q({open_n19579,wb_ill_ins}));  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*B*~(~C*~A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000011001000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u4118|_al_u7211  (
    .a({open_n19580,_al_u7210_o}),
    .b({open_n19581,\cu_ru/medeleg_exc_ctrl/n80_neg_lutinv }),
    .c({_al_u4117_o,_al_u4126_o}),
    .d({\cu_ru/medeleg_exc_ctrl/n80_neg_lutinv ,_al_u4128_o}),
    .f({\cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o ,_al_u7211_o}));
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4119|cu_ru/medeleg_exc_ctrl/diaf_reg  (
    .b({open_n19604,\cu_ru/stval [1]}),
    .c({wb_ins_acc_fault,data_csr[1]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/medeleg [1],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n19608,data_csr[1]}),
    .sr(rst_pad),
    .f({_al_u4119_o,_al_u5347_o}),
    .q({open_n19623,\cu_ru/medeleg [1]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(~C*~(B*~D))"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b0000111100000011),
    .MODE("LOGIC"))
    \_al_u4121|_al_u4120  (
    .b({_al_u4119_o,\cu_ru/medeleg [1]}),
    .c({\cu_ru/medeleg_exc_ctrl/iaf_target_m_lutinv ,wb_ins_acc_fault}),
    .d({\cu_ru/m_s_status/n5 [1],priv[3]}),
    .f({_al_u4121_o,\cu_ru/medeleg_exc_ctrl/iaf_target_m_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4122|_al_u4127  (
    .c({_al_u4121_o,_al_u4126_o}),
    .d({\cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o ,\cu_ru/medeleg_exc_ctrl/n84_neg_lutinv }),
    .f({_al_u4122_o,_al_u4127_o}));
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4123|cu_ru/medeleg_exc_ctrl/dlam_reg  (
    .a({open_n19674,\cu_ru/read_sscratch_sel_lutinv }),
    .b({open_n19675,\cu_ru/read_medeleg_sel_lutinv }),
    .c({wb_ld_addr_mis,\cu_ru/sscratch [4]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/medeleg [4],\cu_ru/medeleg [4]}),
    .mi({open_n19679,data_csr[4]}),
    .sr(rst_pad),
    .f({_al_u4123_o,_al_u7551_o}),
    .q({open_n19694,\cu_ru/medeleg [4]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(~C*~(B*~D))"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b0000111100000011),
    .MODE("LOGIC"))
    \_al_u4125|_al_u4124  (
    .b({_al_u4123_o,\cu_ru/medeleg [4]}),
    .c({\cu_ru/medeleg_exc_ctrl/lam_target_m_lutinv ,wb_ld_addr_mis}),
    .d({\cu_ru/m_s_status/n5 [1],priv[3]}),
    .f({\cu_ru/medeleg_exc_ctrl/n84_neg_lutinv ,\cu_ru/medeleg_exc_ctrl/lam_target_m_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*~(C*~B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1101111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4126|cu_ru/medeleg_exc_ctrl/dsam_reg  (
    .a({\cu_ru/m_s_status/n5 [1],\cu_ru/read_sscratch_sel_lutinv }),
    .b({priv[3],\cu_ru/read_medeleg_sel_lutinv }),
    .c({\cu_ru/medeleg [6],\cu_ru/sscratch [6]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({wb_st_addr_mis,\cu_ru/medeleg [6]}),
    .mi({open_n19727,data_csr[6]}),
    .sr(rst_pad),
    .f({_al_u4126_o,_al_u7341_o}),
    .q({open_n19731,\cu_ru/medeleg [6]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~(~B*~D))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~(~B*~D))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000011000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4128|_al_u3246  (
    .b({priv[1],open_n19734}),
    .c({wb_ecall,priv[1]}),
    .d({priv[0],priv[0]}),
    .f({_al_u4128_o,\cu_ru/m_s_status/n5 [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*~(C*~B)))"),
    //.LUTF1("(~D*B*~(C*A))"),
    //.LUTG0("(A*~(~D*~(C*~B)))"),
    //.LUTG1("(~D*B*~(C*A))"),
    .INIT_LUTF0(16'b1010101000100000),
    .INIT_LUTF1(16'b0000000001001100),
    .INIT_LUTG0(16'b1010101000100000),
    .INIT_LUTG1(16'b0000000001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4129|_al_u6436  (
    .a({_al_u4113_o,_al_u4122_o}),
    .b({_al_u4122_o,_al_u4107_o}),
    .c({_al_u4127_o,_al_u4127_o}),
    .d({_al_u4128_o,_al_u4128_o}),
    .f({\cu_ru/medeleg_exc_ctrl/n98 [2],_al_u6436_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*B))"),
    //.LUT1("(~C*~(~B*D))"),
    .INIT_LUT0(16'b0001010101010101),
    .INIT_LUT1(16'b0000110000001111),
    .MODE("LOGIC"))
    \_al_u4132|_al_u4234  (
    .a({open_n19783,_al_u4138_o}),
    .b({_al_u4131_o,\cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o }),
    .c({_al_u3237_o,_al_u4131_o}),
    .d({\cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o ,_al_u4233_o}),
    .f({_al_u4132_o,_al_u4234_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~D*~C*~B*A)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4134|_al_u5161  (
    .a({_al_u4133_o,open_n19804}),
    .b({wb_st_acc_fault,open_n19805}),
    .c({wb_st_addr_mis,wb_ebreak}),
    .d({wb_st_page_fault,_al_u4133_o}),
    .f({_al_u4134_o,_al_u5161_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4136|_al_u5353  (
    .b({wb_ebreak,open_n19832}),
    .c({wb_ecall,wb_ebreak}),
    .d({_al_u4135_o,int_req}),
    .f({_al_u4136_o,_al_u5353_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4137|_al_u5098  (
    .c({_al_u4136_o,wb_int_acc}),
    .d({_al_u4134_o,_al_u4137_o}),
    .f({_al_u4137_o,_al_u5098_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4138|_al_u2844  (
    .c({wb_valid,wb_valid}),
    .d({_al_u4137_o,1'b0}),
    .f({_al_u4138_o,_al_u2844_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4139|cu_ru/m_s_ie/meie_reg  (
    .b({\cu_ru/m_sip [11],open_n19911}),
    .c({\cu_ru/mie ,_al_u3195_o}),
    .ce(\cu_ru/m_s_ie/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_sie [11],_al_u3191_o}),
    .mi({open_n19915,data_csr[11]}),
    .sr(rst_pad),
    .f({_al_u4139_o,\cu_ru/m_s_ie/n0 }),
    .q({open_n19930,\cu_ru/m_sie [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(D*~(C*~B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b1101111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4143|cu_ru/medeleg_exc_ctrl/dipf_reg  (
    .a({\cu_ru/m_s_status/n5 [1],open_n19931}),
    .b({priv[3],\cu_ru/stval [12]}),
    .c({\cu_ru/medeleg [12],data_csr[12]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({wb_ins_page_fault,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n19942,data_csr[12]}),
    .sr(rst_pad),
    .f({_al_u4143_o,_al_u5338_o}),
    .q({open_n19946,\cu_ru/medeleg [12]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUT1("~(~B*~(C*~(~D*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001111),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4144|cu_ru/m_s_cause/reg1_b2  (
    .a({\cu_ru/medeleg_exc_ctrl/n98 [2],open_n19947}),
    .b({_al_u4140_o,\cu_ru/trap_cause [2]}),
    .c({_al_u4142_o,\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u4143_o,_al_u6700_o}),
    .sr(rst_pad),
    .f({\cu_ru/trap_cause [2],open_n19961}),
    .q({open_n19965,\cu_ru/mcause [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4146|biu/cache_ctrl_logic/reg7_b15  (
    .b({uncache_data[15],open_n19968}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[15]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [15],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [15],uncache_data[15]}),
    .q({open_n19984,\biu/cache_ctrl_logic/pte_temp [15]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4148|biu/cache_ctrl_logic/reg7_b14  (
    .b({uncache_data[14],open_n19987}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[14]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [14],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [14],uncache_data[14]}),
    .q({open_n20007,\biu/cache_ctrl_logic/pte_temp [14]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4150|biu/cache_ctrl_logic/reg7_b13  (
    .b({uncache_data[13],open_n20010}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[13]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [13],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [13],uncache_data[13]}),
    .q({open_n20026,\biu/cache_ctrl_logic/pte_temp [13]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4152|biu/cache_ctrl_logic/reg7_b12  (
    .b({uncache_data[12],open_n20029}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[12]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [12],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [12],uncache_data[12]}),
    .q({open_n20045,\biu/cache_ctrl_logic/pte_temp [12]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4154|biu/cache_ctrl_logic/reg7_b11  (
    .b({uncache_data[11],open_n20048}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[11]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [11],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [11],uncache_data[11]}),
    .q({open_n20068,\biu/cache_ctrl_logic/pte_temp [11]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4156|biu/cache_ctrl_logic/reg7_b10  (
    .b({uncache_data[10],open_n20071}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[10]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [10],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [10],uncache_data[10]}),
    .q({open_n20091,\biu/cache_ctrl_logic/pte_temp [10]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u4158|_al_u7919  (
    .a({open_n20092,uncache_data[9]}),
    .b({uncache_data[9],uncache_data[25]}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,addr_ex[0]}),
    .d({\exu/lsu/n4 [9],addr_ex[1]}),
    .f({\biu/l1i_in [9],_al_u7919_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4160|biu/cache_ctrl_logic/reg7_b8  (
    .b({uncache_data[8],open_n20115}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[8]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [8],_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [8],uncache_data[8]}),
    .q({open_n20135,\biu/cache_ctrl_logic/pte_temp [8]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~B*~A)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~D*C*~B*~A)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000010000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000010000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4161|_al_u4162  (
    .a({open_n20136,_al_u4161_o}),
    .b({open_n20137,_al_u3216_o}),
    .c({\ins_dec/op_amo ,_al_u3217_o}),
    .d({\ins_dec/op_store ,_al_u3384_o}),
    .f({_al_u4161_o,_al_u4162_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4163|_al_u9115  (
    .b({_al_u3217_o,open_n20164}),
    .c({_al_u3384_o,rd_data_slt}),
    .d({\ins_dec/op_load ,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .f({\ins_dec/n48_lutinv ,\exu/alu_au/n39 [0]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4165|_al_u4178  (
    .c({_al_u3213_o,id_ins[16]}),
    .d({\ins_dec/mux24_b10_sel_is_0_o ,_al_u3214_o}),
    .f({_al_u4165_o,_al_u4178_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4166|ins_dec/reg8_b9  (
    .a({open_n20217,_al_u4166_o}),
    .b({open_n20218,_al_u4167_o}),
    .c({id_ins[29],_al_u4064_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4165_o,id_ins[28]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4166_o,open_n20235}),
    .q({open_n20239,as2[9]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4169|ins_dec/reg8_b8  (
    .a({open_n20240,_al_u4169_o}),
    .b({open_n20241,_al_u4170_o}),
    .c({id_ins[28],_al_u4064_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4165_o,id_ins[27]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4169_o,open_n20254}),
    .q({open_n20258,as2[8]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4170|_al_u4167  (
    .c({id_ins[19],id_ins[20]}),
    .d({_al_u3214_o,_al_u3214_o}),
    .f({_al_u4170_o,_al_u4167_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4172|ins_dec/reg8_b7  (
    .a({open_n20283,_al_u4172_o}),
    .b({open_n20284,_al_u4173_o}),
    .c({id_ins[27],_al_u4064_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4165_o,id_ins[26]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4172_o,open_n20301}),
    .q({open_n20305,as2[7]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C*~D))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0011001111110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4175|ins_dec/reg8_b6  (
    .a({_al_u3214_o,open_n20306}),
    .b({_al_u4064_o,_al_u4175_o}),
    .c({id_ins[25],id_ins[26]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[17],_al_u4165_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4175_o,open_n20323}),
    .q({open_n20327,as2[6]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4177|ins_dec/reg8_b5  (
    .a({open_n20328,_al_u4177_o}),
    .b({open_n20329,_al_u4178_o}),
    .c({id_ins[25],_al_u4064_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4165_o,id_ins[11]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4177_o,open_n20342}),
    .q({open_n20346,as2[5]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4182|ins_dec/reg8_b10  (
    .a({open_n20347,_al_u4182_o}),
    .b({open_n20348,_al_u4183_o}),
    .c({id_ins[30],_al_u4064_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4165_o,id_ins[29]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4182_o,open_n20361}),
    .q({open_n20365,as2[10]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4183|_al_u6207  (
    .b({open_n20368,_al_u3927_o}),
    .c({id_ins[21],id_ins[21]}),
    .d({_al_u3214_o,_al_u4086_o}),
    .f({_al_u4183_o,_al_u6207_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u4185|_al_u6112  (
    .b({\ins_dec/funct3_0_lutinv ,open_n20391}),
    .c({_al_u3927_o,_al_u3216_o}),
    .d({_al_u3926_o,\ins_dec/n239 }),
    .f({_al_u4185_o,_al_u6112_o}));
  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(D*C*A))"),
    //.LUT1("(C*~B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110110011001100),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4188|ins_dec/mem_csr_data_ds2_reg  (
    .a({open_n20412,_al_u3938_o}),
    .b({_al_u3217_o,\ins_dec/n141_lutinv }),
    .c({_al_u3384_o,_al_u3399_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_system,id_ins[27]}),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/n141_lutinv ,open_n20425}),
    .q({open_n20429,mem_csr_data_ds2}));  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4190|_al_u2893  (
    .b({open_n20432,\biu/bus_unit/addr_counter [7]}),
    .c({\biu/bus_unit/statu [0],\biu/bus_unit/last_addr [7]}),
    .d({_al_u3407_o,_al_u2890_o}),
    .f({\biu/bus_unit/n26 [0],_al_u2893_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C)*~(A)+~(D*~B)*C*~(A)+~(~(D*~B))*C*A+~(D*~B)*C*A)"),
    //.LUTF1("~(~D*~(B)*~((~C*A))+~D*B*~((~C*A))+~(~D)*B*(~C*A)+~D*B*(~C*A))"),
    //.LUTG0("(~(D*~B)*~(C)*~(A)+~(D*~B)*C*~(A)+~(~(D*~B))*C*A+~(D*~B)*C*A)"),
    //.LUTG1("~(~D*~(B)*~((~C*A))+~D*B*~((~C*A))+~(~D)*B*(~C*A)+~D*B*(~C*A))"),
    .INIT_LUTF0(16'b1110010011110101),
    .INIT_LUTF1(16'b1111011100000010),
    .INIT_LUTG0(16'b1110010011110101),
    .INIT_LUTG1(16'b1111011100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4191|_al_u4100  (
    .a({\biu/bus_unit/mux10_b3_sel_is_0_o ,_al_u2890_o}),
    .b({\biu/bus_unit/n26 [0],_al_u3407_o}),
    .c({_al_u2890_o,_al_u4099_o}),
    .d({_al_u4099_o,\biu/bus_unit/statu [3]}),
    .f({_al_u4191_o,_al_u4100_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~D*~(C*A)))"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(B*~(~D*~(C*A)))"),
    //.LUTG1("(~C*B*D)"),
    .INIT_LUTF0(16'b1100110010000000),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b1100110010000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4193|_al_u4192  (
    .a({open_n20481,\biu/bus_unit/n15_lutinv }),
    .b({_al_u2957_o,htrans_pad[0]}),
    .c({_al_u4192_o,hready_pad}),
    .d({_al_u4191_o,hresp_pad}),
    .f({_al_u4193_o,_al_u4192_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(~D*~C*~B*A)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"))
    \_al_u4194|_al_u2834  (
    .a({_al_u2833_o,open_n20506}),
    .b({\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ,open_n20507}),
    .c({\biu/cache_ctrl_logic/n75_lutinv ,rst_pad}),
    .d({_al_u2885_o,_al_u2833_o}),
    .f({_al_u4194_o,\biu/bus_unit/n37 }));
  // ../../RTL/CPU/BIU/bus_unit.v(163)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(~D*~A)))"),
    //.LUT1("(D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000000110001),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4197|biu/bus_unit/reg1_b0  (
    .a({open_n20528,_al_u4193_o}),
    .b({\biu/bus_unit/mmu/mux10_b0_sel_is_2_o ,_al_u4194_o}),
    .c({\biu/bus_unit/statu [0],_al_u4197_o}),
    .clk(clk_pad),
    .d({_al_u2704_o,_al_u2958_o}),
    .sr(rst_pad),
    .f({_al_u4197_o,open_n20542}),
    .q({open_n20546,\biu/bus_unit/statu [0]}));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4199|_al_u4202  (
    .a({open_n20547,\biu/cache_ctrl_logic/n149 }),
    .b({_al_u2905_o,_al_u4199_o}),
    .c({_al_u2907_o,_al_u4200_o}),
    .d({_al_u2903_o,_al_u4201_o}),
    .f({_al_u4199_o,\biu/cache_ctrl_logic/n140 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4200|_al_u2894  (
    .b({open_n20574,_al_u2893_o}),
    .c({_al_u2893_o,addr_ex[7]}),
    .d({_al_u2891_o,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .f({_al_u4200_o,\biu/l1d_addr [7]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4201|_al_u2902  (
    .a({_al_u2895_o,open_n20599}),
    .b({_al_u2897_o,_al_u2901_o}),
    .c({_al_u2899_o,addr_ex[3]}),
    .d({_al_u2901_o,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .f({_al_u4201_o,\biu/l1d_addr [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u4205|_al_u4204  (
    .b({\exu/alu_data_mem_csr [9],open_n20626}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[1]}),
    .d({_al_u4203_o,addr_ex[0]}),
    .f({_al_u4205_o,\exu/lsu/n2_lutinv }));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4206|biu/cache_ctrl_logic/reg7_b17  (
    .b({uncache_data[17],open_n20649}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[17]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4205_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [17],uncache_data[17]}),
    .q({open_n20669,\biu/cache_ctrl_logic/pte_temp [17]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b1111010100111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1111010100111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4208|_al_u4392  (
    .a({open_n20670,\exu/alu_data_mem_csr [8]}),
    .b({\exu/alu_data_mem_csr [8],\exu/alu_data_mem_csr [16]}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[0]}),
    .d({_al_u4207_o,addr_ex[1]}),
    .f({_al_u4208_o,_al_u4392_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4209|biu/cache_ctrl_logic/reg7_b16  (
    .b({uncache_data[16],open_n20697}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[16]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4208_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [16],uncache_data[16]}),
    .q({open_n20713,\biu/cache_ctrl_logic/pte_temp [16]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0000000010101100),
    .INIT_LUTF1(16'b1111010100111111),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b1111010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4210|_al_u4145  (
    .a({\exu/alu_data_mem_csr [7],\exu/alu_data_mem_csr [7]}),
    .b({\exu/alu_data_mem_csr [15],\exu/alu_data_mem_csr [15]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4210_o,\exu/lsu/n4 [15]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4212|biu/cache_ctrl_logic/reg7_b23  (
    .b({uncache_data[23],open_n20740}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[23]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4211_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [23],uncache_data[23]}),
    .q({open_n20756,\biu/cache_ctrl_logic/pte_temp [23]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0000000010101100),
    .INIT_LUTF1(16'b1111010100111111),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b1111010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4213|_al_u4147  (
    .a({\exu/alu_data_mem_csr [6],\exu/alu_data_mem_csr [6]}),
    .b({\exu/alu_data_mem_csr [14],\exu/alu_data_mem_csr [14]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4213_o,\exu/lsu/n4 [14]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1111001101011111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111001101011111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4214|_al_u4368  (
    .a({open_n20781,\exu/alu_data_mem_csr [22]}),
    .b({\exu/alu_data_mem_csr [22],\exu/alu_data_mem_csr [14]}),
    .c({\exu/lsu/n0_lutinv ,addr_ex[0]}),
    .d({_al_u4213_o,addr_ex[1]}),
    .f({_al_u4214_o,_al_u4368_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4215|biu/cache_ctrl_logic/reg7_b22  (
    .b({uncache_data[22],open_n20808}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[22]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4214_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [22],uncache_data[22]}),
    .q({open_n20828,\biu/cache_ctrl_logic/pte_temp [22]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b0000000010101100),
    .INIT_LUT1(16'b1111010100111111),
    .MODE("LOGIC"))
    \_al_u4216|_al_u4149  (
    .a({\exu/alu_data_mem_csr [5],\exu/alu_data_mem_csr [5]}),
    .b({\exu/alu_data_mem_csr [13],\exu/alu_data_mem_csr [13]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4216_o,\exu/lsu/n4 [13]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*~D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(B*~(~C*~D))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1100110011000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100110011000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4217|_al_u5128  (
    .b({\exu/alu_data_mem_csr [21],_al_u5127_o}),
    .c({\exu/lsu/n0_lutinv ,_al_u3222_o}),
    .d({_al_u4216_o,_al_u4217_o}),
    .f({_al_u4217_o,_al_u5128_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4218|biu/cache_ctrl_logic/reg7_b21  (
    .b({uncache_data[21],open_n20877}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[21]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4217_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [21],uncache_data[21]}),
    .q({open_n20897,\biu/cache_ctrl_logic/pte_temp [21]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b0000000010101100),
    .INIT_LUT1(16'b1111010100111111),
    .MODE("LOGIC"))
    \_al_u4219|_al_u4151  (
    .a({\exu/alu_data_mem_csr [4],\exu/alu_data_mem_csr [4]}),
    .b({\exu/alu_data_mem_csr [12],\exu/alu_data_mem_csr [12]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4219_o,\exu/lsu/n4 [12]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1111001101011111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111001101011111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4220|_al_u4376  (
    .a({open_n20918,\exu/alu_data_mem_csr [20]}),
    .b({\exu/alu_data_mem_csr [20],\exu/alu_data_mem_csr [12]}),
    .c({\exu/lsu/n0_lutinv ,addr_ex[0]}),
    .d({_al_u4219_o,addr_ex[1]}),
    .f({_al_u4220_o,_al_u4376_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4221|biu/cache_ctrl_logic/reg7_b20  (
    .b({uncache_data[20],open_n20945}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[20]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4220_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [20],uncache_data[20]}),
    .q({open_n20961,\biu/cache_ctrl_logic/pte_temp [20]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0000000010101100),
    .INIT_LUTF1(16'b1111010100111111),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b1111010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4222|_al_u4153  (
    .a({\exu/alu_data_mem_csr [3],\exu/alu_data_mem_csr [3]}),
    .b({\exu/alu_data_mem_csr [11],\exu/alu_data_mem_csr [11]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4222_o,\exu/lsu/n4 [11]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4224|biu/cache_ctrl_logic/reg7_b19  (
    .b({uncache_data[19],open_n20988}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[19]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4223_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [19],uncache_data[19]}),
    .q({open_n21004,\biu/cache_ctrl_logic/pte_temp [19]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0000000010101100),
    .INIT_LUTF1(16'b1111010100111111),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b1111010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4225|_al_u4155  (
    .a({\exu/alu_data_mem_csr [2],\exu/alu_data_mem_csr [2]}),
    .b({\exu/alu_data_mem_csr [10],\exu/alu_data_mem_csr [10]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4225_o,\exu/lsu/n4 [10]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*~D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(B*~(~C*~D))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1100110011000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100110011000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4226|_al_u5140  (
    .b({\exu/alu_data_mem_csr [18],_al_u5139_o}),
    .c({\exu/lsu/n0_lutinv ,_al_u3222_o}),
    .d({_al_u4225_o,_al_u4226_o}),
    .f({_al_u4226_o,_al_u5140_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4227|biu/cache_ctrl_logic/reg7_b18  (
    .b({uncache_data[18],open_n21057}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[18]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4226_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [18],uncache_data[18]}),
    .q({open_n21077,\biu/cache_ctrl_logic/pte_temp [18]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*~(~D*B*~A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*~(~D*B*~A))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111100001011),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4230|_al_u4229  (
    .a({_al_u4113_o,open_n21078}),
    .b({_al_u4127_o,open_n21079}),
    .c({_al_u4229_o,wb_ecall}),
    .d({_al_u4128_o,priv[1]}),
    .f({_al_u4230_o,_al_u4229_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"))
    \_al_u4231|_al_u4232  (
    .a({_al_u4230_o,open_n21104}),
    .b({\cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o ,_al_u4138_o}),
    .c({_al_u4143_o,_al_u4141_o}),
    .d({_al_u4121_o,\cu_ru/medeleg_exc_ctrl/n99 [0]}),
    .f({\cu_ru/medeleg_exc_ctrl/n99 [0],_al_u4232_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4233|_al_u4142  (
    .c({_al_u4139_o,_al_u4141_o}),
    .d({\cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ,_al_u4138_o}),
    .f({_al_u4233_o,_al_u4142_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("~(~C*~D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("~(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4235|cu_ru/m_s_cause/reg1_b63  (
    .b({open_n21155,\cu_ru/trap_target_m }),
    .c({_al_u4234_o,_al_u4234_o}),
    .clk(clk_pad),
    .d({_al_u4232_o,_al_u6698_o}),
    .sr(rst_pad),
    .f({\cu_ru/trap_cause [0],open_n21173}),
    .q({open_n21177,\cu_ru/mcause [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011111111110101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011111111110101),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4238|_al_u4237  (
    .a({open_n21178,\exu/alu_data_mem_csr [63]}),
    .b({open_n21179,\exu/alu_data_mem_csr [39]}),
    .c({_al_u4237_o,addr_ex[0]}),
    .d({_al_u4236_o,addr_ex[1]}),
    .f({_al_u4238_o,_al_u4237_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4239|biu/cache_ctrl_logic/reg7_b63  (
    .b({uncache_data[63],open_n21206}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[63]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4238_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [63],uncache_data[63]}),
    .q({open_n21226,\biu/cache_ctrl_logic/pte_temp [63]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0000110000001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4240|exu/reg2_b62  (
    .a({\exu/alu_data_mem_csr [62],open_n21227}),
    .b({\exu/alu_data_mem_csr [46],_al_u3468_o}),
    .c({addr_ex[0],\exu/alu_au/n55 [62]}),
    .clk(clk_pad),
    .d({addr_ex[1],\exu/alu_au/n53 [62]}),
    .sr(rst_pad),
    .f({_al_u4240_o,\exu/alu_data_mem_csr [62]}),
    .q({open_n21244,data_csr[62]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUTF0(16'b0000110000001010),
    .INIT_LUTF1(16'b1100000010100000),
    .INIT_LUTG0(16'b0000110000001010),
    .INIT_LUTG1(16'b1100000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4241|_al_u4272  (
    .a({\exu/alu_data_mem_csr [54],\exu/alu_data_mem_csr [54]}),
    .b({\exu/alu_data_mem_csr [38],\exu/alu_data_mem_csr [38]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4241_o,_al_u4272_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    .INIT_LUT0(16'b0000000000001111),
    .MODE("LOGIC"))
    _al_u4242 (
    .c({open_n21273,_al_u4241_o}),
    .d({open_n21276,_al_u4240_o}),
    .f({open_n21290,_al_u4242_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4243|biu/cache_ctrl_logic/reg7_b62  (
    .b({uncache_data[62],open_n21298}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[62]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4242_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [62],uncache_data[62]}),
    .q({open_n21314,\biu/cache_ctrl_logic/pte_temp [62]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0011111111110101),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0011111111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4245|exu/reg2_b61  (
    .a({\exu/alu_data_mem_csr [61],open_n21315}),
    .b({\exu/alu_data_mem_csr [37],_al_u3476_o}),
    .c({addr_ex[0],\exu/alu_au/n55 [61]}),
    .clk(clk_pad),
    .d({addr_ex[1],\exu/alu_au/n53 [61]}),
    .sr(rst_pad),
    .f({_al_u4245_o,\exu/alu_data_mem_csr [61]}),
    .q({open_n21336,data_csr[61]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111001101011111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111001101011111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4246|_al_u4244  (
    .a({open_n21337,\exu/alu_data_mem_csr [53]}),
    .b({open_n21338,\exu/alu_data_mem_csr [45]}),
    .c({_al_u4245_o,addr_ex[0]}),
    .d({_al_u4244_o,addr_ex[1]}),
    .f({_al_u4246_o,_al_u4244_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4247|biu/cache_ctrl_logic/reg7_b61  (
    .b({uncache_data[61],open_n21365}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[61]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4246_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [61],uncache_data[61]}),
    .q({open_n21381,\biu/cache_ctrl_logic/pte_temp [61]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0000110000001010),
    .INIT_LUTF1(16'b1111001101011111),
    .INIT_LUTG0(16'b0000110000001010),
    .INIT_LUTG1(16'b1111001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4248|_al_u4312  (
    .a({\exu/alu_data_mem_csr [52],\exu/alu_data_mem_csr [44]}),
    .b({\exu/alu_data_mem_csr [44],\exu/alu_data_mem_csr [28]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4248_o,_al_u4312_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0011111111110101),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0011111111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4249|exu/reg2_b60  (
    .a({\exu/alu_data_mem_csr [60],open_n21406}),
    .b({\exu/alu_data_mem_csr [36],_al_u3484_o}),
    .c({addr_ex[0],\exu/alu_au/n55 [60]}),
    .clk(clk_pad),
    .d({addr_ex[1],\exu/alu_au/n53 [60]}),
    .sr(rst_pad),
    .f({_al_u4249_o,\exu/alu_data_mem_csr [60]}),
    .q({open_n21427,data_csr[60]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4250|_al_u4254  (
    .c({_al_u4249_o,_al_u4253_o}),
    .d({_al_u4248_o,_al_u4252_o}),
    .f({_al_u4250_o,_al_u4254_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4251|biu/cache_ctrl_logic/reg7_b60  (
    .b({uncache_data[60],open_n21458}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[60]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4250_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [60],uncache_data[60]}),
    .q({open_n21478,\biu/cache_ctrl_logic/pte_temp [60]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0000110000001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4252|exu/reg2_b59  (
    .a({\exu/alu_data_mem_csr [59],open_n21479}),
    .b({\exu/alu_data_mem_csr [43],_al_u3499_o}),
    .c({addr_ex[0],\exu/alu_au/n55 [59]}),
    .clk(clk_pad),
    .d({addr_ex[1],\exu/alu_au/n53 [59]}),
    .sr(rst_pad),
    .f({_al_u4252_o,\exu/alu_data_mem_csr [59]}),
    .q({open_n21496,data_csr[59]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b1100000010100000),
    .MODE("LOGIC"))
    \_al_u4253|_al_u4284  (
    .a({\exu/alu_data_mem_csr [51],\exu/alu_data_mem_csr [51]}),
    .b({\exu/alu_data_mem_csr [35],\exu/alu_data_mem_csr [35]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4253_o,_al_u4284_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4255|biu/cache_ctrl_logic/reg7_b59  (
    .b({uncache_data[59],open_n21519}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[59]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4254_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [59],uncache_data[59]}),
    .q({open_n21539,\biu/cache_ctrl_logic/pte_temp [59]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*B*~D)"),
    //.LUT1("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110011),
    .INIT_LUT1(16'b0000110000001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4256|exu/reg2_b58  (
    .a({\exu/alu_data_mem_csr [58],open_n21540}),
    .b({\exu/alu_data_mem_csr [42],_al_u3507_o}),
    .c({addr_ex[0],\exu/alu_au/n55 [58]}),
    .clk(clk_pad),
    .d({addr_ex[1],\exu/alu_au/n53 [58]}),
    .sr(rst_pad),
    .f({_al_u4256_o,\exu/alu_data_mem_csr [58]}),
    .q({open_n21557,data_csr[58]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUTF0(16'b0000110000001010),
    .INIT_LUTF1(16'b1100000010100000),
    .INIT_LUTG0(16'b0000110000001010),
    .INIT_LUTG1(16'b1100000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4257|_al_u4288  (
    .a({\exu/alu_data_mem_csr [50],\exu/alu_data_mem_csr [50]}),
    .b({\exu/alu_data_mem_csr [34],\exu/alu_data_mem_csr [34]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4257_o,_al_u4288_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4258|_al_u6818  (
    .b({open_n21584,_al_u6816_o}),
    .c({_al_u4257_o,_al_u6817_o}),
    .d({_al_u4256_o,_al_u6815_o}),
    .f({_al_u4258_o,_al_u6818_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4259|biu/cache_ctrl_logic/reg7_b58  (
    .b({uncache_data[58],open_n21607}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[58]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4258_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [58],uncache_data[58]}),
    .q({open_n21627,\biu/cache_ctrl_logic/pte_temp [58]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0011111111110101),
    .INIT_LUTF1(16'b1111001101011111),
    .INIT_LUTG0(16'b0011111111110101),
    .INIT_LUTG1(16'b1111001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4260|_al_u4293  (
    .a({\exu/alu_data_mem_csr [49],\exu/alu_data_mem_csr [49]}),
    .b({\exu/alu_data_mem_csr [41],\exu/alu_data_mem_csr [25]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4260_o,_al_u4293_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0011111111110101),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0011111111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4261|exu/reg2_b57  (
    .a({\exu/alu_data_mem_csr [57],open_n21652}),
    .b({\exu/alu_data_mem_csr [33],_al_u3515_o}),
    .c({addr_ex[0],\exu/alu_au/n55 [57]}),
    .clk(clk_pad),
    .d({addr_ex[1],\exu/alu_au/n53 [57]}),
    .sr(rst_pad),
    .f({_al_u4261_o,\exu/alu_data_mem_csr [57]}),
    .q({open_n21673,data_csr[57]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4262|_al_u5702  (
    .b({open_n21676,_al_u5701_o}),
    .c({_al_u4261_o,_al_u3222_o}),
    .d({_al_u4260_o,_al_u4262_o}),
    .f({_al_u4262_o,_al_u5702_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4263|biu/cache_ctrl_logic/reg7_b57  (
    .b({uncache_data[57],open_n21699}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[57]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4262_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [57],uncache_data[57]}),
    .q({open_n21715,\biu/cache_ctrl_logic/pte_temp [57]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*~D)"),
    //.LUTF1("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("~(~C*B*~D)"),
    //.LUTG1("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110011),
    .INIT_LUTF1(16'b0000110000001010),
    .INIT_LUTG0(16'b1111111111110011),
    .INIT_LUTG1(16'b0000110000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4264|exu/reg2_b56  (
    .a({\exu/alu_data_mem_csr [56],open_n21716}),
    .b({\exu/alu_data_mem_csr [40],_al_u3523_o}),
    .c({addr_ex[0],\exu/alu_au/n55 [56]}),
    .clk(clk_pad),
    .d({addr_ex[1],\exu/alu_au/n53 [56]}),
    .sr(rst_pad),
    .f({_al_u4264_o,\exu/alu_data_mem_csr [56]}),
    .q({open_n21737,data_csr[56]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4266|_al_u4265  (
    .a({open_n21738,\exu/alu_data_mem_csr [48]}),
    .b({open_n21739,\exu/alu_data_mem_csr [32]}),
    .c({_al_u4265_o,addr_ex[0]}),
    .d({_al_u4264_o,addr_ex[1]}),
    .f({_al_u4266_o,_al_u4265_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4267|biu/cache_ctrl_logic/reg7_b56  (
    .b({uncache_data[56],open_n21762}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[56]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4266_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [56],uncache_data[56]}),
    .q({open_n21778,\biu/cache_ctrl_logic/pte_temp [56]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b0011111111110101),
    .MODE("LOGIC"))
    \_al_u4269|_al_u4364  (
    .a({\exu/alu_data_mem_csr [55],\exu/alu_data_mem_csr [31]}),
    .b({\exu/alu_data_mem_csr [31],\exu/alu_data_mem_csr [15]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4269_o,_al_u4364_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111001101011111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111001101011111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4270|_al_u4268  (
    .a({open_n21799,\exu/alu_data_mem_csr [47]}),
    .b({open_n21800,\exu/alu_data_mem_csr [39]}),
    .c({_al_u4269_o,addr_ex[0]}),
    .d({_al_u4268_o,addr_ex[1]}),
    .f({_al_u4270_o,_al_u4268_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4271|biu/cache_ctrl_logic/reg7_b55  (
    .b({uncache_data[55],open_n21827}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[55]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4270_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [55],uncache_data[55]}),
    .q({open_n21843,\biu/cache_ctrl_logic/pte_temp [55]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b1111001101011111),
    .INIT_LUT1(16'b1100000010100000),
    .MODE("LOGIC"))
    \_al_u4273|_al_u4336  (
    .a({\exu/alu_data_mem_csr [46],\exu/alu_data_mem_csr [30]}),
    .b({\exu/alu_data_mem_csr [30],\exu/alu_data_mem_csr [22]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4273_o,_al_u4336_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4274|_al_u4457  (
    .b({open_n21866,_al_u4455_o}),
    .c({_al_u4273_o,_al_u4456_o}),
    .d({_al_u4272_o,_al_u4454_o}),
    .f({_al_u4274_o,_al_u4457_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4275|biu/cache_ctrl_logic/reg7_b54  (
    .b({uncache_data[54],open_n21893}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[54]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4274_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [54],uncache_data[54]}),
    .q({open_n21913,\biu/cache_ctrl_logic/pte_temp [54]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b1100000010100000),
    .MODE("LOGIC"))
    \_al_u4277|_al_u4372  (
    .a({\exu/alu_data_mem_csr [45],\exu/alu_data_mem_csr [29]}),
    .b({\exu/alu_data_mem_csr [29],\exu/alu_data_mem_csr [13]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4277_o,_al_u4372_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000110000001010),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000110000001010),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4278|_al_u4276  (
    .a({open_n21934,\exu/alu_data_mem_csr [53]}),
    .b({open_n21935,\exu/alu_data_mem_csr [37]}),
    .c({_al_u4277_o,addr_ex[0]}),
    .d({_al_u4276_o,addr_ex[1]}),
    .f({_al_u4278_o,_al_u4276_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4279|biu/cache_ctrl_logic/reg7_b53  (
    .b({uncache_data[53],open_n21962}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[53]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4278_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [53],uncache_data[53]}),
    .q({open_n21982,\biu/cache_ctrl_logic/pte_temp [53]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b1111001101011111),
    .INIT_LUT1(16'b1100000010100000),
    .MODE("LOGIC"))
    \_al_u4281|_al_u4344  (
    .a({\exu/alu_data_mem_csr [44],\exu/alu_data_mem_csr [28]}),
    .b({\exu/alu_data_mem_csr [28],\exu/alu_data_mem_csr [20]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4281_o,_al_u4344_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4282|_al_u4280  (
    .a({open_n22003,\exu/alu_data_mem_csr [52]}),
    .b({open_n22004,\exu/alu_data_mem_csr [36]}),
    .c({_al_u4281_o,addr_ex[0]}),
    .d({_al_u4280_o,addr_ex[1]}),
    .f({_al_u4282_o,_al_u4280_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4283|biu/cache_ctrl_logic/reg7_b52  (
    .b({uncache_data[52],open_n22027}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[52]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4282_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [52],uncache_data[52]}),
    .q({open_n22047,\biu/cache_ctrl_logic/pte_temp [52]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b1100000010100000),
    .MODE("LOGIC"))
    \_al_u4285|_al_u4380  (
    .a({\exu/alu_data_mem_csr [43],\exu/alu_data_mem_csr [27]}),
    .b({\exu/alu_data_mem_csr [27],\exu/alu_data_mem_csr [11]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4285_o,_al_u4380_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4286|_al_u5727  (
    .b({open_n22070,_al_u2705_o}),
    .c({_al_u4285_o,\biu/bus_unit/mmu_hwdata [51]}),
    .d({_al_u4284_o,_al_u5726_o}),
    .f({_al_u4286_o,hwdata_pad[51]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4287|biu/cache_ctrl_logic/reg7_b51  (
    .b({uncache_data[51],open_n22097}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[51]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4286_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [51],uncache_data[51]}),
    .q({open_n22113,\biu/cache_ctrl_logic/pte_temp [51]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUT1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b0011111111110101),
    .INIT_LUT1(16'b1100000010100000),
    .MODE("LOGIC"))
    \_al_u4289|_al_u4321  (
    .a({\exu/alu_data_mem_csr [42],\exu/alu_data_mem_csr [42]}),
    .b({\exu/alu_data_mem_csr [26],\exu/alu_data_mem_csr [18]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4289_o,_al_u4321_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*~D))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(B*~(~C*~D))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1100110011000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1100110011000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4290|_al_u5730  (
    .b({open_n22136,_al_u5729_o}),
    .c({_al_u4289_o,_al_u3222_o}),
    .d({_al_u4288_o,_al_u4290_o}),
    .f({_al_u4290_o,_al_u5730_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4291|biu/cache_ctrl_logic/reg7_b50  (
    .b({uncache_data[50],open_n22163}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[50]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4290_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [50],uncache_data[50]}),
    .q({open_n22179,\biu/cache_ctrl_logic/pte_temp [50]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111001101011111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4294|_al_u4292  (
    .a({open_n22180,\exu/alu_data_mem_csr [41]}),
    .b({open_n22181,\exu/alu_data_mem_csr [33]}),
    .c({_al_u4293_o,addr_ex[0]}),
    .d({_al_u4292_o,addr_ex[1]}),
    .f({_al_u4294_o,_al_u4292_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4295|biu/cache_ctrl_logic/reg7_b49  (
    .b({uncache_data[49],open_n22204}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[49]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4294_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [49],uncache_data[49]}),
    .q({open_n22224,\biu/cache_ctrl_logic/pte_temp [49]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b1111001101011111),
    .MODE("LOGIC"))
    \_al_u4296|_al_u4328  (
    .a({\exu/alu_data_mem_csr [40],\exu/alu_data_mem_csr [40]}),
    .b({\exu/alu_data_mem_csr [32],\exu/alu_data_mem_csr [24]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4296_o,_al_u4328_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT_LUTF0(16'b1111001101011111),
    .INIT_LUTF1(16'b0011111111110101),
    .INIT_LUTG0(16'b1111001101011111),
    .INIT_LUTG1(16'b0011111111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4297|_al_u4360  (
    .a({\exu/alu_data_mem_csr [48],\exu/alu_data_mem_csr [24]}),
    .b({\exu/alu_data_mem_csr [24],\exu/alu_data_mem_csr [16]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4297_o,_al_u4360_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4298|_al_u7169  (
    .b({open_n22271,_al_u7167_o}),
    .c({_al_u4297_o,_al_u7168_o}),
    .d({_al_u4296_o,_al_u7166_o}),
    .f({_al_u4298_o,_al_u7169_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4299|biu/cache_ctrl_logic/reg7_b48  (
    .b({uncache_data[48],open_n22298}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[48]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4298_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [48],uncache_data[48]}),
    .q({open_n22318,\biu/cache_ctrl_logic/pte_temp [48]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUTF0(16'b1111001101011111),
    .INIT_LUTF1(16'b0000110000001010),
    .INIT_LUTG0(16'b1111001101011111),
    .INIT_LUTG1(16'b0000110000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4300|_al_u4332  (
    .a({\exu/alu_data_mem_csr [47],\exu/alu_data_mem_csr [31]}),
    .b({\exu/alu_data_mem_csr [31],\exu/alu_data_mem_csr [23]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4300_o,_al_u4332_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4302|_al_u4301  (
    .a({open_n22343,\exu/alu_data_mem_csr [39]}),
    .b({open_n22344,\exu/alu_data_mem_csr [23]}),
    .c({_al_u4301_o,addr_ex[0]}),
    .d({_al_u4300_o,addr_ex[1]}),
    .f({_al_u4302_o,_al_u4301_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4303|biu/cache_ctrl_logic/reg7_b47  (
    .b({uncache_data[47],open_n22371}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[47]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4302_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [47],uncache_data[47]}),
    .q({open_n22387,\biu/cache_ctrl_logic/pte_temp [47]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111001101011111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4306|_al_u4304  (
    .a({open_n22388,\exu/alu_data_mem_csr [38]}),
    .b({open_n22389,\exu/alu_data_mem_csr [30]}),
    .c({_al_u4305_o,addr_ex[0]}),
    .d({_al_u4304_o,addr_ex[1]}),
    .f({_al_u4306_o,_al_u4304_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4307|biu/cache_ctrl_logic/reg7_b46  (
    .b({uncache_data[46],open_n22412}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[46]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4306_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [46],uncache_data[46]}),
    .q({open_n22428,\biu/cache_ctrl_logic/pte_temp [46]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUTF0(16'b1111001101011111),
    .INIT_LUTF1(16'b0000110000001010),
    .INIT_LUTG0(16'b1111001101011111),
    .INIT_LUTG1(16'b0000110000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4308|_al_u4340  (
    .a({\exu/alu_data_mem_csr [45],\exu/alu_data_mem_csr [29]}),
    .b({\exu/alu_data_mem_csr [29],\exu/alu_data_mem_csr [21]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4308_o,_al_u4340_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4310|_al_u4309  (
    .a({open_n22453,\exu/alu_data_mem_csr [37]}),
    .b({open_n22454,\exu/alu_data_mem_csr [21]}),
    .c({_al_u4309_o,addr_ex[0]}),
    .d({_al_u4308_o,addr_ex[1]}),
    .f({_al_u4310_o,_al_u4309_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4311|biu/cache_ctrl_logic/reg7_b45  (
    .b({uncache_data[45],open_n22477}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[45]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4310_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [45],uncache_data[45]}),
    .q({open_n22497,\biu/cache_ctrl_logic/pte_temp [45]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4314|_al_u4313  (
    .a({open_n22498,\exu/alu_data_mem_csr [36]}),
    .b({open_n22499,\exu/alu_data_mem_csr [20]}),
    .c({_al_u4313_o,addr_ex[0]}),
    .d({_al_u4312_o,addr_ex[1]}),
    .f({_al_u4314_o,_al_u4313_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4315|biu/cache_ctrl_logic/reg7_b44  (
    .b({uncache_data[44],open_n22526}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[44]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4314_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [44],uncache_data[44]}),
    .q({open_n22546,\biu/cache_ctrl_logic/pte_temp [44]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b1111001101011111),
    .INIT_LUTF1(16'b1111001101011111),
    .INIT_LUTG0(16'b1111001101011111),
    .INIT_LUTG1(16'b1111001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4316|_al_u4348  (
    .a({\exu/alu_data_mem_csr [35],\exu/alu_data_mem_csr [27]}),
    .b({\exu/alu_data_mem_csr [27],\exu/alu_data_mem_csr [19]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4316_o,_al_u4348_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011111111110101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011111111110101),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4318|_al_u4317  (
    .a({open_n22571,\exu/alu_data_mem_csr [43]}),
    .b({open_n22572,\exu/alu_data_mem_csr [19]}),
    .c({_al_u4317_o,addr_ex[0]}),
    .d({_al_u4316_o,addr_ex[1]}),
    .f({_al_u4318_o,_al_u4317_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4319|biu/cache_ctrl_logic/reg7_b43  (
    .b({uncache_data[43],open_n22599}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[43]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4318_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [43],uncache_data[43]}),
    .q({open_n22619,\biu/cache_ctrl_logic/pte_temp [43]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111001101011111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111001101011111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4322|_al_u4320  (
    .a({open_n22620,\exu/alu_data_mem_csr [34]}),
    .b({open_n22621,\exu/alu_data_mem_csr [26]}),
    .c({_al_u4321_o,addr_ex[0]}),
    .d({_al_u4320_o,addr_ex[1]}),
    .f({_al_u4322_o,_al_u4320_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4323|biu/cache_ctrl_logic/reg7_b42  (
    .b({uncache_data[42],open_n22648}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[42]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4322_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [42],uncache_data[42]}),
    .q({open_n22664,\biu/cache_ctrl_logic/pte_temp [42]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b0011111111110101),
    .MODE("LOGIC"))
    \_al_u4325|_al_u4203  (
    .a({\exu/alu_data_mem_csr [41],\exu/alu_data_mem_csr [17]}),
    .b({\exu/alu_data_mem_csr [17],\exu/alu_data_mem_csr [1]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4325_o,_al_u4203_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111001101011111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4326|_al_u4324  (
    .a({open_n22685,\exu/alu_data_mem_csr [33]}),
    .b({open_n22686,\exu/alu_data_mem_csr [25]}),
    .c({_al_u4325_o,addr_ex[0]}),
    .d({_al_u4324_o,addr_ex[1]}),
    .f({_al_u4326_o,_al_u4324_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4327|biu/cache_ctrl_logic/reg7_b41  (
    .b({uncache_data[41],open_n22709}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[41]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4326_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [41],uncache_data[41]}),
    .q({open_n22725,\biu/cache_ctrl_logic/pte_temp [41]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4330|_al_u4329  (
    .a({open_n22726,\exu/alu_data_mem_csr [32]}),
    .b({open_n22727,\exu/alu_data_mem_csr [16]}),
    .c({_al_u4329_o,addr_ex[0]}),
    .d({_al_u4328_o,addr_ex[1]}),
    .f({_al_u4330_o,_al_u4329_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4331|biu/cache_ctrl_logic/reg7_b40  (
    .b({uncache_data[40],open_n22750}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[40]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4330_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [40],uncache_data[40]}),
    .q({open_n22770,\biu/cache_ctrl_logic/pte_temp [40]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011111111110101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011111111110101),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4334|_al_u4333  (
    .a({open_n22771,\exu/alu_data_mem_csr [39]}),
    .b({open_n22772,\exu/alu_data_mem_csr [15]}),
    .c({_al_u4333_o,addr_ex[0]}),
    .d({_al_u4332_o,addr_ex[1]}),
    .f({_al_u4334_o,_al_u4333_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4335|biu/cache_ctrl_logic/reg7_b39  (
    .b({uncache_data[39],open_n22799}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[39]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4334_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [39],uncache_data[39]}),
    .q({open_n22819,\biu/cache_ctrl_logic/pte_temp [39]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011111111110101),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4338|_al_u4337  (
    .a({open_n22820,\exu/alu_data_mem_csr [38]}),
    .b({open_n22821,\exu/alu_data_mem_csr [14]}),
    .c({_al_u4337_o,addr_ex[0]}),
    .d({_al_u4336_o,addr_ex[1]}),
    .f({_al_u4338_o,_al_u4337_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4339|biu/cache_ctrl_logic/reg7_b38  (
    .b({uncache_data[38],open_n22844}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[38]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4338_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [38],uncache_data[38]}),
    .q({open_n22864,\biu/cache_ctrl_logic/pte_temp [38]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011111111110101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011111111110101),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4342|_al_u4341  (
    .a({open_n22865,\exu/alu_data_mem_csr [37]}),
    .b({open_n22866,\exu/alu_data_mem_csr [13]}),
    .c({_al_u4341_o,addr_ex[0]}),
    .d({_al_u4340_o,addr_ex[1]}),
    .f({_al_u4342_o,_al_u4341_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4343|biu/cache_ctrl_logic/reg7_b37  (
    .b({uncache_data[37],open_n22893}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[37]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4342_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [37],uncache_data[37]}),
    .q({open_n22909,\biu/cache_ctrl_logic/pte_temp [37]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011111111110101),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u4346|_al_u4345  (
    .a({open_n22910,\exu/alu_data_mem_csr [36]}),
    .b({open_n22911,\exu/alu_data_mem_csr [12]}),
    .c({_al_u4345_o,addr_ex[0]}),
    .d({_al_u4344_o,addr_ex[1]}),
    .f({_al_u4346_o,_al_u4345_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4347|biu/cache_ctrl_logic/reg7_b36  (
    .b({uncache_data[36],open_n22934}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[36]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4346_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [36],uncache_data[36]}),
    .q({open_n22950,\biu/cache_ctrl_logic/pte_temp [36]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011111111110101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011111111110101),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4350|_al_u4349  (
    .a({open_n22951,\exu/alu_data_mem_csr [35]}),
    .b({open_n22952,\exu/alu_data_mem_csr [11]}),
    .c({_al_u4349_o,addr_ex[0]}),
    .d({_al_u4348_o,addr_ex[1]}),
    .f({_al_u4350_o,_al_u4349_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4351|biu/cache_ctrl_logic/reg7_b35  (
    .b({uncache_data[35],open_n22979}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[35]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4350_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [35],uncache_data[35]}),
    .q({open_n22995,\biu/cache_ctrl_logic/pte_temp [35]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUTF0(16'b0000110000001010),
    .INIT_LUTF1(16'b1100000010100000),
    .INIT_LUTG0(16'b0000110000001010),
    .INIT_LUTG1(16'b1100000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4353|_al_u4384  (
    .a({\exu/alu_data_mem_csr [26],\exu/alu_data_mem_csr [26]}),
    .b({\exu/alu_data_mem_csr [10],\exu/alu_data_mem_csr [10]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4353_o,_al_u4384_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4354|_al_u4352  (
    .a({open_n23020,\exu/alu_data_mem_csr [34]}),
    .b({open_n23021,\exu/alu_data_mem_csr [18]}),
    .c({_al_u4353_o,addr_ex[0]}),
    .d({_al_u4352_o,addr_ex[1]}),
    .f({_al_u4354_o,_al_u4352_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4355|biu/cache_ctrl_logic/reg7_b34  (
    .b({uncache_data[34],open_n23044}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[34]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4354_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [34],uncache_data[34]}),
    .q({open_n23064,\biu/cache_ctrl_logic/pte_temp [34]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b1010000011000000),
    .MODE("LOGIC"))
    \_al_u4357|_al_u4388  (
    .a({\exu/alu_data_mem_csr [9],\exu/alu_data_mem_csr [9]}),
    .b({\exu/alu_data_mem_csr [25],\exu/alu_data_mem_csr [25]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u4357_o,_al_u4388_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4358|_al_u4356  (
    .a({open_n23085,\exu/alu_data_mem_csr [33]}),
    .b({open_n23086,\exu/alu_data_mem_csr [17]}),
    .c({_al_u4357_o,addr_ex[0]}),
    .d({_al_u4356_o,addr_ex[1]}),
    .f({_al_u4358_o,_al_u4356_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4359|biu/cache_ctrl_logic/reg7_b33  (
    .b({uncache_data[33],open_n23109}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[33]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4358_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [33],uncache_data[33]}),
    .q({open_n23129,\biu/cache_ctrl_logic/pte_temp [33]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4362|_al_u4361  (
    .a({open_n23130,\exu/alu_data_mem_csr [8]}),
    .b({open_n23131,\exu/alu_data_mem_csr [32]}),
    .c({_al_u4361_o,addr_ex[0]}),
    .d({_al_u4360_o,addr_ex[1]}),
    .f({_al_u4362_o,_al_u4361_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4363|biu/cache_ctrl_logic/reg7_b32  (
    .b({uncache_data[32],open_n23158}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[32]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4362_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [32],uncache_data[32]}),
    .q({open_n23174,\biu/cache_ctrl_logic/pte_temp [32]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4366|_al_u4365  (
    .a({open_n23175,\exu/alu_data_mem_csr [7]}),
    .b({open_n23176,\exu/alu_data_mem_csr [23]}),
    .c({_al_u4365_o,addr_ex[0]}),
    .d({_al_u4364_o,addr_ex[1]}),
    .f({_al_u4366_o,_al_u4365_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4367|biu/cache_ctrl_logic/reg7_b31  (
    .b({uncache_data[31],open_n23199}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[31]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4366_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [31],uncache_data[31]}),
    .q({open_n23215,\biu/cache_ctrl_logic/pte_temp [31]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4370|_al_u4369  (
    .a({open_n23216,\exu/alu_data_mem_csr [6]}),
    .b({open_n23217,\exu/alu_data_mem_csr [30]}),
    .c({_al_u4369_o,addr_ex[0]}),
    .d({_al_u4368_o,addr_ex[1]}),
    .f({_al_u4370_o,_al_u4369_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4371|biu/cache_ctrl_logic/reg7_b30  (
    .b({uncache_data[30],open_n23244}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[30]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4370_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [30],uncache_data[30]}),
    .q({open_n23260,\biu/cache_ctrl_logic/pte_temp [30]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4374|_al_u4373  (
    .a({open_n23261,\exu/alu_data_mem_csr [5]}),
    .b({open_n23262,\exu/alu_data_mem_csr [21]}),
    .c({_al_u4373_o,addr_ex[0]}),
    .d({_al_u4372_o,addr_ex[1]}),
    .f({_al_u4374_o,_al_u4373_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4375|biu/cache_ctrl_logic/reg7_b29  (
    .b({uncache_data[29],open_n23285}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[29]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4374_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [29],uncache_data[29]}),
    .q({open_n23305,\biu/cache_ctrl_logic/pte_temp [29]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4378|_al_u4377  (
    .a({open_n23306,\exu/alu_data_mem_csr [4]}),
    .b({open_n23307,\exu/alu_data_mem_csr [28]}),
    .c({_al_u4377_o,addr_ex[0]}),
    .d({_al_u4376_o,addr_ex[1]}),
    .f({_al_u4378_o,_al_u4377_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4379|biu/cache_ctrl_logic/reg7_b28  (
    .b({uncache_data[28],open_n23334}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[28]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4378_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [28],uncache_data[28]}),
    .q({open_n23354,\biu/cache_ctrl_logic/pte_temp [28]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4382|_al_u4381  (
    .a({open_n23355,\exu/alu_data_mem_csr [3]}),
    .b({open_n23356,\exu/alu_data_mem_csr [19]}),
    .c({_al_u4381_o,addr_ex[0]}),
    .d({_al_u4380_o,addr_ex[1]}),
    .f({_al_u4382_o,_al_u4381_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4383|biu/cache_ctrl_logic/reg7_b27  (
    .b({uncache_data[27],open_n23379}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[27]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4382_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [27],uncache_data[27]}),
    .q({open_n23395,\biu/cache_ctrl_logic/pte_temp [27]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4386|_al_u4385  (
    .a({open_n23396,\exu/alu_data_mem_csr [2]}),
    .b({open_n23397,\exu/alu_data_mem_csr [18]}),
    .c({_al_u4385_o,addr_ex[0]}),
    .d({_al_u4384_o,addr_ex[1]}),
    .f({_al_u4386_o,_al_u4385_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000110011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4387|biu/cache_ctrl_logic/reg7_b26  (
    .b({uncache_data[26],open_n23424}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[26]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4386_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [26],uncache_data[26]}),
    .q({open_n23440,\biu/cache_ctrl_logic/pte_temp [26]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u4390|_al_u4389  (
    .a({open_n23441,\exu/alu_data_mem_csr [17]}),
    .b({open_n23442,\exu/alu_data_mem_csr [1]}),
    .c({_al_u4389_o,addr_ex[0]}),
    .d({_al_u4388_o,addr_ex[1]}),
    .f({_al_u4390_o,_al_u4389_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4391|biu/cache_ctrl_logic/reg7_b25  (
    .b({uncache_data[25],open_n23465}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[25]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4390_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [25],uncache_data[25]}),
    .q({open_n23485,\biu/cache_ctrl_logic/pte_temp [25]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011111111110101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011111111110101),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4394|_al_u4393  (
    .a({open_n23486,\exu/alu_data_mem_csr [24]}),
    .b({open_n23487,\exu/alu_data_mem_csr [0]}),
    .c({_al_u4393_o,addr_ex[0]}),
    .d({_al_u4392_o,addr_ex[1]}),
    .f({_al_u4394_o,_al_u4393_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4395|biu/cache_ctrl_logic/reg7_b24  (
    .b({uncache_data[24],open_n23514}),
    .c({\biu/bus_unit/mux1_b1_sel_is_0_o ,hrdata_pad[24]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4394_o,_al_u2705_o}),
    .sr(rst_pad),
    .f({\biu/l1i_in [24],uncache_data[24]}),
    .q({open_n23534,\biu/cache_ctrl_logic/pte_temp [24]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4397|biu/cache_ctrl_logic/reg1_b73  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n212 [9],\biu/cache_ctrl_logic/pa_temp [73]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [73],addr_ex[9]}),
    .mi({open_n23545,\biu/cache_ctrl_logic/pa_temp [73]}),
    .sr(rst_pad),
    .f({_al_u4397_o,_al_u4401_o}),
    .q({open_n23549,\biu/cache_ctrl_logic/l1i_pa [73]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4398|ins_fetch/reg0_b9  (
    .a({open_n23550,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[9],\ins_fetch/n1 [7]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4397_o,addr_if[9]}),
    .mi({open_n23554,addr_if[9]}),
    .sr(rst_pad),
    .f({_al_u4398_o,_al_u9301_o}),
    .q({open_n23569,id_ins_pc[9]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~D*C*B*A)"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4399|_al_u2912  (
    .a({_al_u2847_o,_al_u2847_o}),
    .b({\biu/cache_ctrl_logic/statu [2],\biu/cache_ctrl_logic/statu [2]}),
    .c({\biu/cache_ctrl_logic/statu [3],\biu/cache_ctrl_logic/statu [3]}),
    .d({\biu/cache_ctrl_logic/statu [4],\biu/cache_ctrl_logic/statu [4]}),
    .f({_al_u4399_o,\biu/cache_ctrl_logic/n75_lutinv }));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4402|biu/cache_ctrl_logic/reg4_b73  (
    .a({open_n23594,_al_u3947_o}),
    .b({_al_u4400_o,_al_u4399_o}),
    .c({_al_u4401_o,\biu/cache_ctrl_logic/n209 [9]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4398_o,\biu/cache_ctrl_logic/l1d_pa [73]}),
    .mi({open_n23598,\biu/cache_ctrl_logic/pa_temp [73]}),
    .sr(rst_pad),
    .f({_al_u4402_o,_al_u4400_o}),
    .q({open_n23613,\biu/cache_ctrl_logic/l1d_pa [73]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4404|_al_u4752  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [9],\biu/cache_ctrl_logic/n207 [12]}),
    .d({_al_u4402_o,_al_u4751_o}),
    .f({\biu/maddress [9],\biu/maddress [12]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4406|biu/cache_ctrl_logic/reg1_b72  (
    .a({open_n23636,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[8],\biu/cache_ctrl_logic/l1d_pa [72]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4405_o,\biu/cache_ctrl_logic/pa_temp [72]}),
    .mi({open_n23647,\biu/cache_ctrl_logic/pa_temp [72]}),
    .sr(rst_pad),
    .f({_al_u4406_o,_al_u4405_o}),
    .q({open_n23651,\biu/cache_ctrl_logic/l1i_pa [72]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4407|_al_u4549  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [72],\biu/cache_ctrl_logic/l1i_pa [107]}),
    .d({addr_ex[8],addr_ex[43]}),
    .f({_al_u4407_o,_al_u4549_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4408|_al_u4713  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [8],\biu/cache_ctrl_logic/n209 [18]}),
    .d({\biu/cache_ctrl_logic/n212 [8],\biu/cache_ctrl_logic/n212 [18]}),
    .f({_al_u4408_o,_al_u4713_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u4409|_al_u4833  (
    .b({_al_u4407_o,open_n23694}),
    .c({_al_u4408_o,_al_u2952_o}),
    .d({_al_u4406_o,_al_u4832_o}),
    .f({_al_u4409_o,_al_u4833_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4410|_al_u4746  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [8],\biu/cache_ctrl_logic/n207 [13]}),
    .d({_al_u4409_o,_al_u4745_o}),
    .f({\biu/maddress [8],\biu/maddress [13]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4411|_al_u4543  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [71],\biu/cache_ctrl_logic/l1i_pa [108]}),
    .d({addr_ex[7],addr_ex[44]}),
    .f({_al_u4411_o,_al_u4543_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4412|ins_fetch/reg0_b7  (
    .a({open_n23757,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[7],\ins_fetch/n1 [5]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4411_o,addr_if[7]}),
    .mi({open_n23768,addr_if[7]}),
    .sr(rst_pad),
    .f({_al_u4412_o,_al_u9320_o}),
    .q({open_n23772,id_ins_pc[7]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4413|_al_u4683  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [7],\biu/cache_ctrl_logic/n209 [23]}),
    .d({\biu/cache_ctrl_logic/n212 [7],\biu/cache_ctrl_logic/n212 [23]}),
    .f({_al_u4413_o,_al_u4683_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4415|biu/cache_ctrl_logic/reg1_b71  (
    .a({open_n23797,_al_u3945_o}),
    .b({_al_u4413_o,_al_u3947_o}),
    .c({_al_u4414_o,\biu/cache_ctrl_logic/l1d_pa [71]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4412_o,\biu/cache_ctrl_logic/pa_temp [71]}),
    .mi({open_n23808,\biu/cache_ctrl_logic/pa_temp [71]}),
    .sr(rst_pad),
    .f({_al_u4415_o,_al_u4414_o}),
    .q({open_n23812,\biu/cache_ctrl_logic/l1i_pa [71]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4416|_al_u4740  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [7],\biu/cache_ctrl_logic/n207 [14]}),
    .d({_al_u4415_o,_al_u4739_o}),
    .f({\biu/maddress [7],\biu/maddress [14]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4418|biu/cache_ctrl_logic/reg1_b127  (
    .a({open_n23839,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[63],\biu/cache_ctrl_logic/l1d_pa [127]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4417_o,\biu/cache_ctrl_logic/pa_temp [127]}),
    .mi({open_n23850,\biu/cache_ctrl_logic/pa_temp [127]}),
    .sr(rst_pad),
    .f({_al_u4418_o,_al_u4417_o}),
    .q({open_n23854,\biu/cache_ctrl_logic/l1i_pa [127]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4420|_al_u4672  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [63],\biu/cache_ctrl_logic/n209 [25]}),
    .d({\biu/cache_ctrl_logic/n212 [63],\biu/cache_ctrl_logic/n212 [25]}),
    .f({_al_u4420_o,_al_u4672_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4421|_al_u4419  (
    .a({open_n23879,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4419_o,_al_u3950_o}),
    .c({_al_u4420_o,\biu/cache_ctrl_logic/l1i_pa [127]}),
    .d({_al_u4418_o,addr_ex[63]}),
    .f({_al_u4421_o,_al_u4419_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4422|_al_u4734  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [63],\biu/cache_ctrl_logic/n207 [15]}),
    .d({_al_u4421_o,_al_u4733_o}),
    .f({\biu/maddress [63],\biu/maddress [15]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4425|_al_u4687  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/n212 [62],\biu/cache_ctrl_logic/n212 [22]}),
    .d({\biu/cache_ctrl_logic/l1i_pa [126],\biu/cache_ctrl_logic/l1i_pa [86]}),
    .f({_al_u4425_o,_al_u4687_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4427|biu/cache_ctrl_logic/reg1_b126  (
    .a({open_n23954,_al_u3945_o}),
    .b({_al_u4425_o,_al_u3947_o}),
    .c({_al_u4426_o,\biu/cache_ctrl_logic/l1d_pa [126]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4424_o,\biu/cache_ctrl_logic/pa_temp [126]}),
    .mi({open_n23958,\biu/cache_ctrl_logic/pa_temp [126]}),
    .sr(rst_pad),
    .f({_al_u4427_o,_al_u4426_o}),
    .q({open_n23973,\biu/cache_ctrl_logic/l1i_pa [126]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4428|_al_u4728  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [62],\biu/cache_ctrl_logic/n207 [16]}),
    .d({_al_u4427_o,_al_u4727_o}),
    .f({\biu/maddress [62],\biu/maddress [16]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u4429|_al_u4659  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/n212 [61],\biu/cache_ctrl_logic/n212 [27]}),
    .d({\biu/cache_ctrl_logic/l1i_pa [125],\biu/cache_ctrl_logic/l1i_pa [91]}),
    .f({_al_u4429_o,_al_u4659_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4430|biu/cache_ctrl_logic/reg0_b61  (
    .a({open_n24016,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[61],\ins_fetch/n1 [59]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4429_o,addr_if[61]}),
    .mi({open_n24027,addr_if[61]}),
    .sr(rst_pad),
    .f({_al_u4430_o,_al_u9325_o}),
    .q({open_n24031,\biu/cache_ctrl_logic/l1i_va [61]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4433|biu/cache_ctrl_logic/reg1_b125  (
    .a({open_n24032,_al_u3945_o}),
    .b({_al_u4431_o,_al_u3947_o}),
    .c({_al_u4432_o,\biu/cache_ctrl_logic/l1d_pa [125]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4430_o,\biu/cache_ctrl_logic/pa_temp [125]}),
    .mi({open_n24036,\biu/cache_ctrl_logic/pa_temp [125]}),
    .sr(rst_pad),
    .f({_al_u4433_o,_al_u4432_o}),
    .q({open_n24051,\biu/cache_ctrl_logic/l1i_pa [125]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4434|_al_u4722  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [61],\biu/cache_ctrl_logic/n207 [17]}),
    .d({_al_u4433_o,_al_u4721_o}),
    .f({\biu/maddress [61],\biu/maddress [17]}));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4435|ins_fetch/reg0_b60  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,open_n24074}),
    .b({_al_u4399_o,\biu/bus_unit/mmu/n19_lutinv }),
    .c({\biu/cache_ctrl_logic/n209 [60],addr_if[60]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/n212 [60],_al_u4435_o}),
    .mi({open_n24078,addr_if[60]}),
    .sr(rst_pad),
    .f({_al_u4435_o,_al_u4436_o}),
    .q({open_n24093,id_ins_pc[60]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4439|biu/cache_ctrl_logic/reg4_b124  (
    .a({open_n24094,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4437_o,_al_u3947_o}),
    .c({_al_u4438_o,\biu/cache_ctrl_logic/l1d_pa [124]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4436_o,addr_ex[60]}),
    .mi({open_n24105,\biu/cache_ctrl_logic/pa_temp [124]}),
    .sr(rst_pad),
    .f({_al_u4439_o,_al_u4437_o}),
    .q({open_n24109,\biu/cache_ctrl_logic/l1d_pa [124]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4440|_al_u4716  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [60],\biu/cache_ctrl_logic/n207 [18]}),
    .d({_al_u4439_o,_al_u4715_o}),
    .f({\biu/maddress [60],\biu/maddress [18]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4441|_al_u4822  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [6],\biu/cache_ctrl_logic/n209 [0]}),
    .d({addr_ex[6],addr_ex[0]}),
    .f({_al_u4441_o,_al_u4822_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4442|ins_fetch/reg0_b6  (
    .a({open_n24160,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[6],\ins_fetch/n1 [4]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4441_o,addr_if[6]}),
    .mi({open_n24164,addr_if[6]}),
    .sr(rst_pad),
    .f({_al_u4442_o,_al_u9385_o}),
    .q({open_n24179,id_ins_pc[6]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4445|biu/cache_ctrl_logic/reg4_b70  (
    .a({open_n24180,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4443_o,_al_u3947_o}),
    .c({_al_u4444_o,\biu/cache_ctrl_logic/n212 [6]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4442_o,\biu/cache_ctrl_logic/l1d_pa [70]}),
    .mi({open_n24191,\biu/cache_ctrl_logic/pa_temp [70]}),
    .sr(rst_pad),
    .f({_al_u4445_o,_al_u4443_o}),
    .q({open_n24195,\biu/cache_ctrl_logic/l1d_pa [70]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4446|_al_u4710  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [6],\biu/cache_ctrl_logic/n207 [19]}),
    .d({_al_u4445_o,_al_u4709_o}),
    .f({\biu/maddress [6],\biu/maddress [19]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u4447|_al_u4605  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/n212 [59],\biu/cache_ctrl_logic/n212 [35]}),
    .d({\biu/cache_ctrl_logic/l1i_pa [123],\biu/cache_ctrl_logic/l1i_pa [99]}),
    .f({_al_u4447_o,_al_u4605_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4448|biu/cache_ctrl_logic/reg0_b59  (
    .a({open_n24242,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[59],\ins_fetch/n1 [57]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4447_o,addr_if[59]}),
    .mi({open_n24246,addr_if[59]}),
    .sr(rst_pad),
    .f({_al_u4448_o,_al_u9335_o}),
    .q({open_n24261,\biu/cache_ctrl_logic/l1i_va [59]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4451|biu/cache_ctrl_logic/reg1_b123  (
    .a({open_n24262,_al_u3945_o}),
    .b({_al_u4449_o,_al_u3947_o}),
    .c({_al_u4450_o,\biu/cache_ctrl_logic/l1d_pa [123]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4448_o,\biu/cache_ctrl_logic/pa_temp [123]}),
    .mi({open_n24273,\biu/cache_ctrl_logic/pa_temp [123]}),
    .sr(rst_pad),
    .f({_al_u4451_o,_al_u4450_o}),
    .q({open_n24277,\biu/cache_ctrl_logic/l1i_pa [123]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4452|_al_u4704  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [59],\biu/cache_ctrl_logic/n207 [20]}),
    .d({_al_u4451_o,_al_u4703_o}),
    .f({\biu/maddress [59],\biu/maddress [20]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4454|biu/cache_ctrl_logic/reg1_b122  (
    .a({open_n24300,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[58],\biu/cache_ctrl_logic/l1d_pa [122]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4453_o,\biu/cache_ctrl_logic/pa_temp [122]}),
    .mi({open_n24311,\biu/cache_ctrl_logic/pa_temp [122]}),
    .sr(rst_pad),
    .f({_al_u4454_o,_al_u4453_o}),
    .q({open_n24315,\biu/cache_ctrl_logic/l1i_pa [122]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4455|_al_u4581  (
    .a({_al_u3950_o,_al_u3950_o}),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [58],\biu/cache_ctrl_logic/n209 [39]}),
    .d({\biu/cache_ctrl_logic/l1i_pa [122],\biu/cache_ctrl_logic/l1i_pa [103]}),
    .f({_al_u4455_o,_al_u4581_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4456|_al_u4732  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .c({\biu/cache_ctrl_logic/n212 [58],\biu/cache_ctrl_logic/n212 [15]}),
    .d({addr_ex[58],addr_ex[15]}),
    .f({_al_u4456_o,_al_u4732_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4458|_al_u4698  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [58],\biu/cache_ctrl_logic/n207 [21]}),
    .d({_al_u4457_o,_al_u4697_o}),
    .f({\biu/maddress [58],\biu/maddress [21]}));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4459|ins_fetch/reg0_b57  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,open_n24382}),
    .b({_al_u3950_o,\biu/bus_unit/mmu/n19_lutinv }),
    .c({\biu/cache_ctrl_logic/n212 [57],addr_if[57]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [121],_al_u4459_o}),
    .mi({open_n24393,addr_if[57]}),
    .sr(rst_pad),
    .f({_al_u4459_o,_al_u4460_o}),
    .q({open_n24397,id_ins_pc[57]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4463|biu/cache_ctrl_logic/reg1_b121  (
    .a({open_n24398,_al_u3945_o}),
    .b({_al_u4461_o,_al_u3947_o}),
    .c({_al_u4462_o,\biu/cache_ctrl_logic/l1d_pa [121]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4460_o,\biu/cache_ctrl_logic/pa_temp [121]}),
    .mi({open_n24402,\biu/cache_ctrl_logic/pa_temp [121]}),
    .sr(rst_pad),
    .f({_al_u4463_o,_al_u4462_o}),
    .q({open_n24417,\biu/cache_ctrl_logic/l1i_pa [121]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4464|_al_u4692  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [57],\biu/cache_ctrl_logic/n207 [22]}),
    .d({_al_u4463_o,_al_u4691_o}),
    .f({\biu/maddress [57],\biu/maddress [22]}));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4465|ins_fetch/reg0_b56  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,open_n24444}),
    .b({_al_u4399_o,\biu/bus_unit/mmu/n19_lutinv }),
    .c({\biu/cache_ctrl_logic/n209 [56],addr_if[56]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_ex[56],_al_u4465_o}),
    .mi({open_n24455,addr_if[56]}),
    .sr(rst_pad),
    .f({_al_u4465_o,_al_u4466_o}),
    .q({open_n24459,id_ins_pc[56]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4467|_al_u4591  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/n212 [56],\biu/cache_ctrl_logic/n212 [37]}),
    .d({\biu/cache_ctrl_logic/l1i_pa [120],\biu/cache_ctrl_logic/l1i_pa [101]}),
    .f({_al_u4467_o,_al_u4591_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4469|biu/cache_ctrl_logic/reg1_b120  (
    .a({open_n24484,_al_u3945_o}),
    .b({_al_u4467_o,_al_u3947_o}),
    .c({_al_u4468_o,\biu/cache_ctrl_logic/l1d_pa [120]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4466_o,\biu/cache_ctrl_logic/pa_temp [120]}),
    .mi({open_n24488,\biu/cache_ctrl_logic/pa_temp [120]}),
    .sr(rst_pad),
    .f({_al_u4469_o,_al_u4468_o}),
    .q({open_n24503,\biu/cache_ctrl_logic/l1i_pa [120]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4470|_al_u4686  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [56],\biu/cache_ctrl_logic/n207 [23]}),
    .d({_al_u4469_o,_al_u4685_o}),
    .f({\biu/maddress [56],\biu/maddress [23]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4473|biu/cache_ctrl_logic/reg1_b119  (
    .a({_al_u3950_o,_al_u3945_o}),
    .b({_al_u4399_o,_al_u3947_o}),
    .c({\biu/cache_ctrl_logic/n209 [55],\biu/cache_ctrl_logic/l1d_pa [119]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [119],\biu/cache_ctrl_logic/pa_temp [119]}),
    .mi({open_n24540,\biu/cache_ctrl_logic/pa_temp [119]}),
    .sr(rst_pad),
    .f({_al_u4473_o,_al_u4471_o}),
    .q({open_n24544,\biu/cache_ctrl_logic/l1i_pa [119]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4475|ins_fetch/reg0_b55  (
    .b({_al_u4473_o,\biu/bus_unit/mmu/n19_lutinv }),
    .c({_al_u4474_o,addr_if[55]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4472_o,_al_u4471_o}),
    .mi({open_n24550,addr_if[55]}),
    .sr(rst_pad),
    .f({_al_u4475_o,_al_u4472_o}),
    .q({open_n24565,id_ins_pc[55]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4476|_al_u4680  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [55],\biu/cache_ctrl_logic/n207 [24]}),
    .d({_al_u4475_o,_al_u4679_o}),
    .f({\biu/maddress [55],\biu/maddress [24]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4478|biu/cache_ctrl_logic/reg1_b118  (
    .a({open_n24588,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[54],\biu/cache_ctrl_logic/l1d_pa [118]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4477_o,\biu/cache_ctrl_logic/pa_temp [118]}),
    .mi({open_n24599,\biu/cache_ctrl_logic/pa_temp [118]}),
    .sr(rst_pad),
    .f({_al_u4478_o,_al_u4477_o}),
    .q({open_n24603,\biu/cache_ctrl_logic/l1i_pa [118]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4480|_al_u4651  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [54],\biu/cache_ctrl_logic/n209 [28]}),
    .d({\biu/cache_ctrl_logic/n212 [54],\biu/cache_ctrl_logic/n212 [28]}),
    .f({_al_u4480_o,_al_u4651_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4481|_al_u4479  (
    .a({open_n24624,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4479_o,_al_u3950_o}),
    .c({_al_u4480_o,\biu/cache_ctrl_logic/l1i_pa [118]}),
    .d({_al_u4478_o,addr_ex[54]}),
    .f({_al_u4481_o,_al_u4479_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4482|_al_u4674  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [54],\biu/cache_ctrl_logic/n207 [25]}),
    .d({_al_u4481_o,_al_u4673_o}),
    .f({\biu/maddress [54],\biu/maddress [25]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4483|_al_u4639  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [53],\biu/cache_ctrl_logic/n209 [3]}),
    .d({\biu/cache_ctrl_logic/n212 [53],\biu/cache_ctrl_logic/n212 [3]}),
    .f({_al_u4483_o,_al_u4639_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4484|biu/cache_ctrl_logic/reg0_b53  (
    .a({open_n24695,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[53],\ins_fetch/n1 [51]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4483_o,addr_if[53]}),
    .mi({open_n24699,addr_if[53]}),
    .sr(rst_pad),
    .f({_al_u4484_o,_al_u9371_o}),
    .q({open_n24714,\biu/cache_ctrl_logic/l1i_va [53]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4487|biu/cache_ctrl_logic/reg4_b117  (
    .a({open_n24715,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4485_o,_al_u3947_o}),
    .c({_al_u4486_o,\biu/cache_ctrl_logic/l1d_pa [117]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4484_o,addr_ex[53]}),
    .mi({open_n24726,\biu/cache_ctrl_logic/pa_temp [117]}),
    .sr(rst_pad),
    .f({_al_u4487_o,_al_u4485_o}),
    .q({open_n24730,\biu/cache_ctrl_logic/l1d_pa [117]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4488|_al_u4668  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [53],\biu/cache_ctrl_logic/n207 [26]}),
    .d({_al_u4487_o,_al_u4667_o}),
    .f({\biu/maddress [53],\biu/maddress [26]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4489|_al_u4701  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [52],\biu/cache_ctrl_logic/n209 [20]}),
    .d({addr_ex[52],addr_ex[20]}),
    .f({_al_u4489_o,_al_u4701_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4490|biu/cache_ctrl_logic/reg0_b52  (
    .a({open_n24777,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[52],\ins_fetch/n1 [50]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4489_o,addr_if[52]}),
    .mi({open_n24788,addr_if[52]}),
    .sr(rst_pad),
    .f({_al_u4490_o,_al_u9378_o}),
    .q({open_n24792,\biu/cache_ctrl_logic/l1i_va [52]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4493|biu/cache_ctrl_logic/reg4_b116  (
    .a({open_n24793,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4491_o,_al_u3947_o}),
    .c({_al_u4492_o,\biu/cache_ctrl_logic/n212 [52]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4490_o,\biu/cache_ctrl_logic/l1d_pa [116]}),
    .mi({open_n24797,\biu/cache_ctrl_logic/pa_temp [116]}),
    .sr(rst_pad),
    .f({_al_u4493_o,_al_u4491_o}),
    .q({open_n24812,\biu/cache_ctrl_logic/l1d_pa [116]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4494|_al_u4662  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [52],\biu/cache_ctrl_logic/n207 [27]}),
    .d({_al_u4493_o,_al_u4661_o}),
    .f({\biu/maddress [52],\biu/maddress [27]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4496|biu/cache_ctrl_logic/reg1_b115  (
    .a({open_n24839,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[51],\biu/cache_ctrl_logic/l1d_pa [115]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4495_o,\biu/cache_ctrl_logic/pa_temp [115]}),
    .mi({open_n24843,\biu/cache_ctrl_logic/pa_temp [115]}),
    .sr(rst_pad),
    .f({_al_u4496_o,_al_u4495_o}),
    .q({open_n24858,\biu/cache_ctrl_logic/l1i_pa [115]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4497|_al_u4531  (
    .a({_al_u3950_o,_al_u3950_o}),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [51],\biu/cache_ctrl_logic/n209 [46]}),
    .d({\biu/cache_ctrl_logic/l1i_pa [115],\biu/cache_ctrl_logic/l1i_pa [110]}),
    .f({_al_u4497_o,_al_u4531_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C@B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100001100000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4498|biu/cache_ctrl_logic/reg3_b51  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,open_n24879}),
    .b({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/l1i_va [51]}),
    .c({\biu/cache_ctrl_logic/n212 [51],addr_ex[51]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[51],_al_u6401_o}),
    .mi({open_n24890,addr_ex[51]}),
    .sr(rst_pad),
    .f({_al_u4498_o,_al_u6402_o}),
    .q({open_n24894,\biu/cache_ctrl_logic/l1d_va [51]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u4499|_al_u6315  (
    .b({_al_u4497_o,open_n24897}),
    .c({_al_u4498_o,\biu/cache_ctrl_logic/l1d_pte [4]}),
    .d({_al_u4496_o,\biu/bus_unit/mmu/n7_lutinv }),
    .f({_al_u4499_o,\biu/cache_ctrl_logic/n30 }));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4500|_al_u4656  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [51],\biu/cache_ctrl_logic/n207 [28]}),
    .d({_al_u4499_o,_al_u4655_o}),
    .f({\biu/maddress [51],\biu/maddress [28]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4501|biu/cache_ctrl_logic/reg1_b114  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n212 [50],\biu/cache_ctrl_logic/pa_temp [114]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [114],addr_ex[50]}),
    .mi({open_n24950,\biu/cache_ctrl_logic/pa_temp [114]}),
    .sr(rst_pad),
    .f({_al_u4501_o,_al_u4504_o}),
    .q({open_n24954,\biu/cache_ctrl_logic/l1i_pa [114]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4505|biu/cache_ctrl_logic/reg4_b114  (
    .a({open_n24955,_al_u3947_o}),
    .b({_al_u4503_o,_al_u4399_o}),
    .c({_al_u4504_o,\biu/cache_ctrl_logic/n209 [50]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4502_o,\biu/cache_ctrl_logic/l1d_pa [114]}),
    .mi({open_n24959,\biu/cache_ctrl_logic/pa_temp [114]}),
    .sr(rst_pad),
    .f({_al_u4505_o,_al_u4503_o}),
    .q({open_n24974,\biu/cache_ctrl_logic/l1d_pa [114]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4506|_al_u4650  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [50],\biu/cache_ctrl_logic/n207 [29]}),
    .d({_al_u4505_o,_al_u4649_o}),
    .f({\biu/maddress [50],\biu/maddress [29]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4507|_al_u4612  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [5],\biu/cache_ctrl_logic/n209 [34]}),
    .d({\biu/cache_ctrl_logic/n212 [5],\biu/cache_ctrl_logic/n212 [34]}),
    .f({_al_u4507_o,_al_u4612_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4508|ins_fetch/reg0_b5  (
    .a({open_n25017,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[5],\ins_fetch/n1 [3]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4507_o,addr_if[5]}),
    .mi({open_n25021,addr_if[5]}),
    .sr(rst_pad),
    .f({_al_u4508_o,_al_u9456_o}),
    .q({open_n25036,id_ins_pc[5]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4509|_al_u4617  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [69],\biu/cache_ctrl_logic/l1i_pa [97]}),
    .d({addr_ex[5],addr_ex[33]}),
    .f({_al_u4509_o,_al_u4617_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4511|biu/cache_ctrl_logic/reg1_b69  (
    .a({open_n25057,_al_u3945_o}),
    .b({_al_u4509_o,_al_u3947_o}),
    .c({_al_u4510_o,\biu/cache_ctrl_logic/l1d_pa [69]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4508_o,\biu/cache_ctrl_logic/pa_temp [69]}),
    .mi({open_n25061,\biu/cache_ctrl_logic/pa_temp [69]}),
    .sr(rst_pad),
    .f({_al_u4511_o,_al_u4510_o}),
    .q({open_n25076,\biu/cache_ctrl_logic/l1i_pa [69]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4512|_al_u4584  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [5],\biu/cache_ctrl_logic/n207 [39]}),
    .d({_al_u4511_o,_al_u4583_o}),
    .f({\biu/maddress [5],\biu/maddress [39]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4514|biu/cache_ctrl_logic/reg1_b113  (
    .a({open_n25103,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[49],\biu/cache_ctrl_logic/l1d_pa [113]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4513_o,\biu/cache_ctrl_logic/pa_temp [113]}),
    .mi({open_n25107,\biu/cache_ctrl_logic/pa_temp [113]}),
    .sr(rst_pad),
    .f({_al_u4514_o,_al_u4513_o}),
    .q({open_n25122,\biu/cache_ctrl_logic/l1i_pa [113]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4516|exu/reg5_b49  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,open_n25123}),
    .b({\biu/cache_ctrl_logic/n97_lutinv ,open_n25124}),
    .c({\biu/cache_ctrl_logic/n212 [49],addr_ex[49]}),
    .clk(clk_pad),
    .d({addr_ex[49],ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({_al_u4516_o,open_n25138}),
    .q({open_n25142,wb_exc_code[49]}));  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4517|_al_u4515  (
    .a({open_n25143,_al_u3950_o}),
    .b({_al_u4515_o,_al_u4399_o}),
    .c({_al_u4516_o,\biu/cache_ctrl_logic/n209 [49]}),
    .d({_al_u4514_o,\biu/cache_ctrl_logic/l1i_pa [113]}),
    .f({_al_u4517_o,_al_u4515_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4518|_al_u4572  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [49],\biu/cache_ctrl_logic/n207 [40]}),
    .d({_al_u4517_o,_al_u4571_o}),
    .f({\biu/maddress [49],\biu/maddress [40]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4520|biu/cache_ctrl_logic/reg1_b112  (
    .a({open_n25190,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[48],\biu/cache_ctrl_logic/l1d_pa [112]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4519_o,\biu/cache_ctrl_logic/pa_temp [112]}),
    .mi({open_n25201,\biu/cache_ctrl_logic/pa_temp [112]}),
    .sr(rst_pad),
    .f({_al_u4520_o,_al_u4519_o}),
    .q({open_n25205,\biu/cache_ctrl_logic/l1i_pa [112]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("~(C@D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4521|biu/cache_ctrl_logic/reg3_b48  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,open_n25206}),
    .b({_al_u3950_o,open_n25207}),
    .c({\biu/cache_ctrl_logic/l1i_pa [112],addr_ex[48]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[48],\biu/cache_ctrl_logic/l1i_va [48]}),
    .mi({open_n25218,addr_ex[48]}),
    .sr(rst_pad),
    .f({_al_u4521_o,_al_u6365_o}),
    .q({open_n25222,\biu/cache_ctrl_logic/l1d_va [48]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4522|_al_u4555  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [48],\biu/cache_ctrl_logic/n209 [42]}),
    .d({\biu/cache_ctrl_logic/n212 [48],\biu/cache_ctrl_logic/n212 [42]}),
    .f({_al_u4522_o,_al_u4555_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4523|_al_u6291  (
    .a({open_n25243,_al_u6276_o}),
    .b({_al_u4521_o,_al_u6280_o}),
    .c({_al_u4522_o,_al_u6285_o}),
    .d({_al_u4520_o,_al_u6290_o}),
    .f({_al_u4523_o,_al_u6291_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4524|_al_u4566  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [48],\biu/cache_ctrl_logic/n207 [41]}),
    .d({_al_u4523_o,_al_u4565_o}),
    .f({\biu/maddress [48],\biu/maddress [41]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4527|biu/cache_ctrl_logic/reg1_b111  (
    .a({_al_u3950_o,_al_u3945_o}),
    .b({_al_u4399_o,_al_u3947_o}),
    .c({\biu/cache_ctrl_logic/n209 [47],\biu/cache_ctrl_logic/l1d_pa [111]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [111],\biu/cache_ctrl_logic/pa_temp [111]}),
    .mi({open_n25300,\biu/cache_ctrl_logic/pa_temp [111]}),
    .sr(rst_pad),
    .f({_al_u4527_o,_al_u4525_o}),
    .q({open_n25304,\biu/cache_ctrl_logic/l1i_pa [111]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4529|ins_fetch/reg0_b47  (
    .b({_al_u4527_o,\biu/bus_unit/mmu/n19_lutinv }),
    .c({_al_u4528_o,addr_if[47]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4526_o,_al_u4525_o}),
    .mi({open_n25310,addr_if[47]}),
    .sr(rst_pad),
    .f({_al_u4529_o,_al_u4526_o}),
    .q({open_n25325,id_ins_pc[47]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4530|_al_u4560  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [47],\biu/cache_ctrl_logic/n207 [42]}),
    .d({_al_u4529_o,_al_u4559_o}),
    .f({\biu/maddress [47],\biu/maddress [42]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4532|biu/cache_ctrl_logic/reg0_b46  (
    .a({open_n25352,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[46],\ins_fetch/n1 [44]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4531_o,addr_if[46]}),
    .mi({open_n25363,addr_if[46]}),
    .sr(rst_pad),
    .f({_al_u4532_o,_al_u9425_o}),
    .q({open_n25367,\biu/cache_ctrl_logic/l1i_va [46]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4533|_al_u4666  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .c({\biu/cache_ctrl_logic/n212 [46],\biu/cache_ctrl_logic/n212 [26]}),
    .d({addr_ex[46],addr_ex[26]}),
    .f({_al_u4533_o,_al_u4666_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4535|biu/cache_ctrl_logic/reg1_b110  (
    .a({open_n25388,_al_u3945_o}),
    .b({_al_u4533_o,_al_u3947_o}),
    .c({_al_u4534_o,\biu/cache_ctrl_logic/l1d_pa [110]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4532_o,\biu/cache_ctrl_logic/pa_temp [110]}),
    .mi({open_n25392,\biu/cache_ctrl_logic/pa_temp [110]}),
    .sr(rst_pad),
    .f({_al_u4535_o,_al_u4534_o}),
    .q({open_n25407,\biu/cache_ctrl_logic/l1i_pa [110]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4536|_al_u4554  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [46],\biu/cache_ctrl_logic/n207 [43]}),
    .d({_al_u4535_o,_al_u4553_o}),
    .f({\biu/maddress [46],\biu/maddress [43]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4537|biu/cache_ctrl_logic/reg1_b109  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n212 [45],\biu/cache_ctrl_logic/pa_temp [109]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [109],addr_ex[45]}),
    .mi({open_n25437,\biu/cache_ctrl_logic/pa_temp [109]}),
    .sr(rst_pad),
    .f({_al_u4537_o,_al_u4540_o}),
    .q({open_n25452,\biu/cache_ctrl_logic/l1i_pa [109]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4541|biu/cache_ctrl_logic/reg4_b109  (
    .a({open_n25453,_al_u3947_o}),
    .b({_al_u4539_o,_al_u4399_o}),
    .c({_al_u4540_o,\biu/cache_ctrl_logic/n209 [45]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4538_o,\biu/cache_ctrl_logic/l1d_pa [109]}),
    .mi({open_n25464,\biu/cache_ctrl_logic/pa_temp [109]}),
    .sr(rst_pad),
    .f({_al_u4541_o,_al_u4539_o}),
    .q({open_n25468,\biu/cache_ctrl_logic/l1d_pa [109]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4542|_al_u4548  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c(\biu/cache_ctrl_logic/n207 [45:44]),
    .d({_al_u4541_o,_al_u4547_o}),
    .f(\biu/maddress [45:44]));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100110001),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4544|ins_fetch/reg0_b44  (
    .a({open_n25491,\biu/cache_ctrl_logic/l1i_va [44]}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,\biu/cache_ctrl_logic/l1i_va [54]}),
    .c({addr_if[44],addr_if[44]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4543_o,addr_if[54]}),
    .mi({open_n25502,addr_if[44]}),
    .sr(rst_pad),
    .f({_al_u4544_o,_al_u9254_o}),
    .q({open_n25506,id_ins_pc[44]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4545|_al_u4551  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c(\biu/cache_ctrl_logic/n209 [44:43]),
    .d(\biu/cache_ctrl_logic/n212 [44:43]),
    .f({_al_u4545_o,_al_u4551_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4547|biu/cache_ctrl_logic/reg1_b108  (
    .a({open_n25531,_al_u3945_o}),
    .b({_al_u4545_o,_al_u3947_o}),
    .c({_al_u4546_o,\biu/cache_ctrl_logic/l1d_pa [108]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4544_o,\biu/cache_ctrl_logic/pa_temp [108]}),
    .mi({open_n25535,\biu/cache_ctrl_logic/pa_temp [108]}),
    .sr(rst_pad),
    .f({_al_u4547_o,_al_u4546_o}),
    .q({open_n25550,\biu/cache_ctrl_logic/l1i_pa [108]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4550|biu/cache_ctrl_logic/reg0_b43  (
    .a({open_n25551,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[43],\ins_fetch/n1 [41]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4549_o,addr_if[43]}),
    .mi({open_n25555,addr_if[43]}),
    .sr(rst_pad),
    .f({_al_u4550_o,_al_u9444_o}),
    .q({open_n25570,\biu/cache_ctrl_logic/l1i_va [43]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4553|biu/cache_ctrl_logic/reg1_b107  (
    .a({open_n25571,_al_u3945_o}),
    .b({_al_u4551_o,_al_u3947_o}),
    .c({_al_u4552_o,\biu/cache_ctrl_logic/l1d_pa [107]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4550_o,\biu/cache_ctrl_logic/pa_temp [107]}),
    .mi({open_n25582,\biu/cache_ctrl_logic/pa_temp [107]}),
    .sr(rst_pad),
    .f({_al_u4553_o,_al_u4552_o}),
    .q({open_n25586,\biu/cache_ctrl_logic/l1i_pa [107]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4556|_al_u2914  (
    .b({\biu/bus_unit/mmu/n19_lutinv ,open_n25589}),
    .c({addr_if[42],\biu/bus_unit/mmu/n19_lutinv }),
    .d({_al_u4555_o,\biu/cache_ctrl_logic/n75_lutinv }),
    .f({_al_u4556_o,_al_u2914_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4559|biu/cache_ctrl_logic/reg4_b106  (
    .a({open_n25610,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4557_o,_al_u3947_o}),
    .c({_al_u4558_o,\biu/cache_ctrl_logic/l1d_pa [106]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4556_o,addr_ex[42]}),
    .mi({open_n25621,\biu/cache_ctrl_logic/pa_temp [106]}),
    .sr(rst_pad),
    .f({_al_u4559_o,_al_u4557_o}),
    .q({open_n25625,\biu/cache_ctrl_logic/l1d_pa [106]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4561|biu/cache_ctrl_logic/reg1_b105  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n212 [41],\biu/cache_ctrl_logic/pa_temp [105]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [105],addr_ex[41]}),
    .mi({open_n25629,\biu/cache_ctrl_logic/pa_temp [105]}),
    .sr(rst_pad),
    .f({_al_u4561_o,_al_u4564_o}),
    .q({open_n25644,\biu/cache_ctrl_logic/l1i_pa [105]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4562|_al_u4742  (
    .b({\biu/bus_unit/mmu/n19_lutinv ,\biu/bus_unit/mmu/n19_lutinv }),
    .c({addr_if[41],addr_if[13]}),
    .d({_al_u4561_o,_al_u4741_o}),
    .f({_al_u4562_o,_al_u4742_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4565|biu/cache_ctrl_logic/reg4_b105  (
    .a({open_n25671,_al_u3947_o}),
    .b({_al_u4563_o,_al_u4399_o}),
    .c({_al_u4564_o,\biu/cache_ctrl_logic/n209 [41]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4562_o,\biu/cache_ctrl_logic/l1d_pa [105]}),
    .mi({open_n25682,\biu/cache_ctrl_logic/pa_temp [105]}),
    .sr(rst_pad),
    .f({_al_u4565_o,_al_u4563_o}),
    .q({open_n25686,\biu/cache_ctrl_logic/l1d_pa [105]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4567|biu/cache_ctrl_logic/reg1_b104  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n212 [40],\biu/cache_ctrl_logic/pa_temp [104]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [104],addr_ex[40]}),
    .mi({open_n25697,\biu/cache_ctrl_logic/pa_temp [104]}),
    .sr(rst_pad),
    .f({_al_u4567_o,_al_u4570_o}),
    .q({open_n25701,\biu/cache_ctrl_logic/l1i_pa [104]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4568|biu/cache_ctrl_logic/reg0_b40  (
    .a({open_n25702,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[40],\ins_fetch/n1 [38]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4567_o,addr_if[40]}),
    .mi({open_n25713,addr_if[40]}),
    .sr(rst_pad),
    .f({_al_u4568_o,_al_u9468_o}),
    .q({open_n25717,\biu/cache_ctrl_logic/l1i_va [40]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4571|biu/cache_ctrl_logic/reg4_b104  (
    .a({open_n25718,_al_u3947_o}),
    .b({_al_u4569_o,_al_u4399_o}),
    .c({_al_u4570_o,\biu/cache_ctrl_logic/n209 [40]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4568_o,\biu/cache_ctrl_logic/l1d_pa [104]}),
    .mi({open_n25722,\biu/cache_ctrl_logic/pa_temp [104]}),
    .sr(rst_pad),
    .f({_al_u4571_o,_al_u4569_o}),
    .q({open_n25737,\biu/cache_ctrl_logic/l1d_pa [104]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4573|_al_u4621  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [4],\biu/cache_ctrl_logic/n209 [32]}),
    .d({addr_ex[4],addr_ex[32]}),
    .f({_al_u4573_o,_al_u4621_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4574|ins_fetch/reg0_b4  (
    .a({open_n25762,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[4],\ins_fetch/n1 [2]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4573_o,addr_if[4]}),
    .mi({open_n25773,addr_if[4]}),
    .sr(rst_pad),
    .f({_al_u4574_o,_al_u9525_o}),
    .q({open_n25777,id_ins_pc[4]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4577|biu/cache_ctrl_logic/reg4_b68  (
    .a({open_n25778,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4575_o,_al_u3947_o}),
    .c({_al_u4576_o,\biu/cache_ctrl_logic/n212 [4]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4574_o,\biu/cache_ctrl_logic/l1d_pa [68]}),
    .mi({open_n25789,\biu/cache_ctrl_logic/pa_temp [68]}),
    .sr(rst_pad),
    .f({_al_u4577_o,_al_u4575_o}),
    .q({open_n25793,\biu/cache_ctrl_logic/l1d_pa [68]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C*~B))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0011000011111111),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4578|_al_u4764  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [4],\biu/cache_ctrl_logic/n207 [10]}),
    .d({_al_u4577_o,_al_u4763_o}),
    .f({\biu/maddress [4],\biu/maddress [10]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4580|biu/cache_ctrl_logic/reg1_b103  (
    .a({open_n25816,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[39],\biu/cache_ctrl_logic/l1d_pa [103]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4579_o,\biu/cache_ctrl_logic/pa_temp [103]}),
    .mi({open_n25827,\biu/cache_ctrl_logic/pa_temp [103]}),
    .sr(rst_pad),
    .f({_al_u4580_o,_al_u4579_o}),
    .q({open_n25831,\biu/cache_ctrl_logic/l1i_pa [103]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4583|exu/reg3_b39  (
    .a({open_n25832,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4581_o,\biu/cache_ctrl_logic/n97_lutinv }),
    .c({_al_u4582_o,\biu/cache_ctrl_logic/n212 [39]}),
    .clk(clk_pad),
    .d({_al_u4580_o,addr_ex[39]}),
    .mi({open_n25844,addr_ex[39]}),
    .sr(rst_pad),
    .f({_al_u4583_o,_al_u4582_o}),
    .q({open_n25848,new_pc[39]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4586|biu/cache_ctrl_logic/reg1_b102  (
    .a({open_n25849,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[38],\biu/cache_ctrl_logic/l1d_pa [102]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4585_o,\biu/cache_ctrl_logic/pa_temp [102]}),
    .mi({open_n25853,\biu/cache_ctrl_logic/pa_temp [102]}),
    .sr(rst_pad),
    .f({_al_u4586_o,_al_u4585_o}),
    .q({open_n25868,\biu/cache_ctrl_logic/l1i_pa [102]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4588|biu/cache_ctrl_logic/reg3_b29  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/l1i_va [29]}),
    .b({_al_u4399_o,\biu/cache_ctrl_logic/l1i_va [38]}),
    .c({\biu/cache_ctrl_logic/n209 [38],addr_ex[29]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[38],addr_ex[38]}),
    .mi({open_n25872,addr_ex[29]}),
    .sr(rst_pad),
    .f({_al_u4588_o,_al_u6416_o}),
    .q({open_n25887,\biu/cache_ctrl_logic/l1d_va [29]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4589|_al_u4587  (
    .a({open_n25888,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4587_o,_al_u3950_o}),
    .c({_al_u4588_o,\biu/cache_ctrl_logic/n212 [38]}),
    .d({_al_u4586_o,\biu/cache_ctrl_logic/l1i_pa [102]}),
    .f({_al_u4589_o,_al_u4587_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0000000011001010),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4590|_al_u6216  (
    .a({open_n25913,\biu/maddress [38]}),
    .b({_al_u4403_o,\biu/maddress [29]}),
    .c({\biu/cache_ctrl_logic/n207 [38],\biu/bus_unit/mmu/i [0]}),
    .d({_al_u4589_o,\biu/bus_unit/mmu/i [1]}),
    .f({\biu/maddress [38],_al_u6216_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4592|biu/cache_ctrl_logic/reg0_b37  (
    .a({open_n25934,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[37],\ins_fetch/n1 [35]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4591_o,addr_if[37]}),
    .mi({open_n25938,addr_if[37]}),
    .sr(rst_pad),
    .f({_al_u4592_o,_al_u9487_o}),
    .q({open_n25953,\biu/cache_ctrl_logic/l1i_va [37]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4595|biu/cache_ctrl_logic/reg4_b101  (
    .a({open_n25954,_al_u3947_o}),
    .b({_al_u4593_o,_al_u4399_o}),
    .c({_al_u4594_o,\biu/cache_ctrl_logic/n209 [37]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4592_o,\biu/cache_ctrl_logic/l1d_pa [101]}),
    .mi({open_n25958,\biu/cache_ctrl_logic/pa_temp [101]}),
    .sr(rst_pad),
    .f({_al_u4595_o,_al_u4593_o}),
    .q({open_n25973,\biu/cache_ctrl_logic/l1d_pa [101]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0000000011001010),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0000000011001010),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4596|_al_u6219  (
    .a({open_n25974,\biu/maddress [37]}),
    .b({_al_u4403_o,\biu/maddress [28]}),
    .c({\biu/cache_ctrl_logic/n207 [37],\biu/bus_unit/mmu/i [0]}),
    .d({_al_u4595_o,\biu/bus_unit/mmu/i [1]}),
    .f({\biu/maddress [37],_al_u6219_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4598|biu/cache_ctrl_logic/reg0_b36  (
    .a({open_n25999,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[36],\ins_fetch/n1 [34]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4597_o,addr_if[36]}),
    .mi({open_n26003,addr_if[36]}),
    .sr(rst_pad),
    .f({_al_u4598_o,_al_u9494_o}),
    .q({open_n26018,\biu/cache_ctrl_logic/l1i_va [36]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4601|biu/cache_ctrl_logic/reg4_b100  (
    .a({open_n26019,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4599_o,_al_u3947_o}),
    .c({_al_u4600_o,\biu/cache_ctrl_logic/n212 [36]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4598_o,\biu/cache_ctrl_logic/l1d_pa [100]}),
    .mi({open_n26030,\biu/cache_ctrl_logic/pa_temp [100]}),
    .sr(rst_pad),
    .f({_al_u4601_o,_al_u4599_o}),
    .q({open_n26034,\biu/cache_ctrl_logic/l1d_pa [100]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0000000011001010),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0000000011001010),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4602|_al_u6222  (
    .a({open_n26035,\biu/maddress [36]}),
    .b({_al_u4403_o,\biu/maddress [27]}),
    .c({\biu/cache_ctrl_logic/n207 [36],\biu/bus_unit/mmu/i [0]}),
    .d({_al_u4601_o,\biu/bus_unit/mmu/i [1]}),
    .f({\biu/maddress [36],_al_u6222_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4604|exu/reg3_b35  (
    .a({open_n26060,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u4399_o}),
    .c({addr_if[35],\biu/cache_ctrl_logic/n209 [35]}),
    .clk(clk_pad),
    .d({_al_u4603_o,addr_ex[35]}),
    .mi({open_n26065,addr_ex[35]}),
    .sr(rst_pad),
    .f({_al_u4604_o,_al_u4603_o}),
    .q({open_n26080,new_pc[35]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4607|biu/cache_ctrl_logic/reg1_b99  (
    .a({open_n26081,_al_u3945_o}),
    .b({_al_u4605_o,_al_u3947_o}),
    .c({_al_u4606_o,\biu/cache_ctrl_logic/l1d_pa [99]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4604_o,\biu/cache_ctrl_logic/pa_temp [99]}),
    .mi({open_n26092,\biu/cache_ctrl_logic/pa_temp [99]}),
    .sr(rst_pad),
    .f({_al_u4607_o,_al_u4606_o}),
    .q({open_n26096,\biu/cache_ctrl_logic/l1i_pa [99]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0000000011001010),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4608|_al_u6225  (
    .a({open_n26097,\biu/maddress [35]}),
    .b({_al_u4403_o,\biu/maddress [26]}),
    .c({\biu/cache_ctrl_logic/n207 [35],\biu/bus_unit/mmu/i [0]}),
    .d({_al_u4607_o,\biu/bus_unit/mmu/i [1]}),
    .f({\biu/maddress [35],_al_u6225_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4610|biu/cache_ctrl_logic/reg1_b98  (
    .a({open_n26118,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[34],\biu/cache_ctrl_logic/l1d_pa [98]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4609_o,\biu/cache_ctrl_logic/pa_temp [98]}),
    .mi({open_n26122,\biu/cache_ctrl_logic/pa_temp [98]}),
    .sr(rst_pad),
    .f({_al_u4610_o,_al_u4609_o}),
    .q({open_n26137,\biu/cache_ctrl_logic/l1i_pa [98]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4613|_al_u4611  (
    .a({open_n26138,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4611_o,_al_u3950_o}),
    .c({_al_u4612_o,\biu/cache_ctrl_logic/l1i_pa [98]}),
    .d({_al_u4610_o,addr_ex[34]}),
    .f({_al_u4613_o,_al_u4611_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0000000011001010),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4614|_al_u6228  (
    .a({open_n26163,\biu/maddress [34]}),
    .b({_al_u4403_o,\biu/maddress [25]}),
    .c({\biu/cache_ctrl_logic/n207 [34],\biu/bus_unit/mmu/i [0]}),
    .d({_al_u4613_o,\biu/bus_unit/mmu/i [1]}),
    .f({\biu/maddress [34],_al_u6228_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4616|_al_u4615  (
    .a({open_n26184,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u4399_o}),
    .c({addr_if[33],\biu/cache_ctrl_logic/n209 [33]}),
    .d({_al_u4615_o,\biu/cache_ctrl_logic/n212 [33]}),
    .f({_al_u4616_o,_al_u4615_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4619|biu/cache_ctrl_logic/reg1_b97  (
    .a({open_n26209,_al_u3945_o}),
    .b({_al_u4617_o,_al_u3947_o}),
    .c({_al_u4618_o,\biu/cache_ctrl_logic/l1d_pa [97]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4616_o,\biu/cache_ctrl_logic/pa_temp [97]}),
    .mi({open_n26213,\biu/cache_ctrl_logic/pa_temp [97]}),
    .sr(rst_pad),
    .f({_al_u4619_o,_al_u4618_o}),
    .q({open_n26228,\biu/cache_ctrl_logic/l1i_pa [97]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0000000011001010),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0000000011001010),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4620|_al_u6231  (
    .a({open_n26229,\biu/maddress [33]}),
    .b({_al_u4403_o,\biu/maddress [24]}),
    .c({\biu/cache_ctrl_logic/n207 [33],\biu/bus_unit/mmu/i [0]}),
    .d({_al_u4619_o,\biu/bus_unit/mmu/i [1]}),
    .f({\biu/maddress [33],_al_u6231_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4622|biu/cache_ctrl_logic/reg0_b32  (
    .a({open_n26254,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[32],\ins_fetch/n1 [30]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4621_o,addr_if[32]}),
    .mi({open_n26265,addr_if[32]}),
    .sr(rst_pad),
    .f({_al_u4622_o,_al_u9518_o}),
    .q({open_n26269,\biu/cache_ctrl_logic/l1i_va [32]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4625|biu/cache_ctrl_logic/reg4_b96  (
    .a({open_n26270,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4623_o,_al_u3947_o}),
    .c({_al_u4624_o,\biu/cache_ctrl_logic/n212 [32]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4622_o,\biu/cache_ctrl_logic/l1d_pa [96]}),
    .mi({open_n26274,\biu/cache_ctrl_logic/pa_temp [96]}),
    .sr(rst_pad),
    .f({_al_u4625_o,_al_u4623_o}),
    .q({open_n26289,\biu/cache_ctrl_logic/l1d_pa [96]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0000000011001010),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0000000011001010),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4626|_al_u6234  (
    .a({open_n26290,\biu/maddress [32]}),
    .b({_al_u4403_o,\biu/maddress [23]}),
    .c({\biu/cache_ctrl_logic/n207 [32],\biu/bus_unit/mmu/i [0]}),
    .d({_al_u4625_o,\biu/bus_unit/mmu/i [1]}),
    .f({\biu/maddress [32],_al_u6234_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4629|biu/cache_ctrl_logic/reg1_b95  (
    .a({_al_u3950_o,_al_u3945_o}),
    .b({_al_u4399_o,_al_u3947_o}),
    .c({\biu/cache_ctrl_logic/n209 [31],\biu/cache_ctrl_logic/l1d_pa [95]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [95],\biu/cache_ctrl_logic/pa_temp [95]}),
    .mi({open_n26325,\biu/cache_ctrl_logic/pa_temp [95]}),
    .sr(rst_pad),
    .f({_al_u4629_o,_al_u4627_o}),
    .q({open_n26329,\biu/cache_ctrl_logic/l1i_pa [95]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4631|ins_fetch/reg0_b31  (
    .b({_al_u4629_o,\biu/bus_unit/mmu/n19_lutinv }),
    .c({_al_u4630_o,addr_if[31]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4628_o,_al_u4627_o}),
    .mi({open_n26342,addr_if[31]}),
    .sr(rst_pad),
    .f({_al_u4631_o,_al_u4628_o}),
    .q({open_n26346,id_ins_pc[31]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0000000011001010),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4632|_al_u6237  (
    .a({open_n26347,\biu/maddress [31]}),
    .b({_al_u4403_o,\biu/maddress [22]}),
    .c({\biu/cache_ctrl_logic/n207 [31],\biu/bus_unit/mmu/i [0]}),
    .d({_al_u4631_o,\biu/bus_unit/mmu/i [1]}),
    .f({\biu/maddress [31],_al_u6237_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4634|_al_u4633  (
    .a({open_n26368,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u4399_o}),
    .c({addr_if[30],\biu/cache_ctrl_logic/n209 [30]}),
    .d({_al_u4633_o,addr_ex[30]}),
    .f({_al_u4634_o,_al_u4633_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4637|biu/cache_ctrl_logic/reg4_b94  (
    .a({open_n26393,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4635_o,_al_u3947_o}),
    .c({_al_u4636_o,\biu/cache_ctrl_logic/n212 [30]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4634_o,\biu/cache_ctrl_logic/l1d_pa [94]}),
    .mi({open_n26404,\biu/cache_ctrl_logic/pa_temp [94]}),
    .sr(rst_pad),
    .f({_al_u4637_o,_al_u4635_o}),
    .q({open_n26408,\biu/cache_ctrl_logic/l1d_pa [94]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("~(D*~(C*~B))"),
    .INIT_LUT0(16'b0000000011001010),
    .INIT_LUT1(16'b0011000011111111),
    .MODE("LOGIC"))
    \_al_u4638|_al_u6240  (
    .a({open_n26409,\biu/maddress [30]}),
    .b({_al_u4403_o,\biu/maddress [21]}),
    .c({\biu/cache_ctrl_logic/n207 [30],\biu/bus_unit/mmu/i [0]}),
    .d({_al_u4637_o,\biu/bus_unit/mmu/i [1]}),
    .f({\biu/maddress [30],_al_u6240_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4640|ins_fetch/reg0_b3  (
    .a({open_n26430,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[3],\ins_fetch/n1 [1]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4639_o,addr_if[3]}),
    .mi({open_n26441,addr_if[3]}),
    .sr(rst_pad),
    .f({_al_u4640_o,_al_u9598_o}),
    .q({open_n26445,id_ins_pc[3]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4643|biu/cache_ctrl_logic/reg4_b67  (
    .a({open_n26446,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4641_o,_al_u3947_o}),
    .c({_al_u4642_o,\biu/cache_ctrl_logic/l1d_pa [67]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4640_o,addr_ex[3]}),
    .mi({open_n26457,\biu/cache_ctrl_logic/pa_temp [67]}),
    .sr(rst_pad),
    .f({_al_u4643_o,_al_u4641_o}),
    .q({open_n26461,\biu/cache_ctrl_logic/l1d_pa [67]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C*~B))"),
    //.LUTF1("~(D*~(C*~B))"),
    //.LUTG0("~(D*~(C*~B))"),
    //.LUTG1("~(D*~(C*~B))"),
    .INIT_LUTF0(16'b0011000011111111),
    .INIT_LUTF1(16'b0011000011111111),
    .INIT_LUTG0(16'b0011000011111111),
    .INIT_LUTG1(16'b0011000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4644|_al_u4758  (
    .b({_al_u4403_o,_al_u4403_o}),
    .c({\biu/cache_ctrl_logic/n207 [3],\biu/cache_ctrl_logic/n207 [11]}),
    .d({_al_u4643_o,_al_u4757_o}),
    .f({\biu/maddress [3],\biu/maddress [11]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4646|_al_u4645  (
    .a({open_n26488,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u4399_o}),
    .c({addr_if[29],\biu/cache_ctrl_logic/n209 [29]}),
    .d({_al_u4645_o,\biu/cache_ctrl_logic/n212 [29]}),
    .f({_al_u4646_o,_al_u4645_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4649|biu/cache_ctrl_logic/reg4_b93  (
    .a({open_n26509,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4647_o,_al_u3947_o}),
    .c({_al_u4648_o,\biu/cache_ctrl_logic/l1d_pa [93]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4646_o,addr_ex[29]}),
    .mi({open_n26513,\biu/cache_ctrl_logic/pa_temp [93]}),
    .sr(rst_pad),
    .f({_al_u4649_o,_al_u4647_o}),
    .q({open_n26528,\biu/cache_ctrl_logic/l1d_pa [93]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4652|biu/cache_ctrl_logic/reg0_b28  (
    .a({open_n26529,\ins_fetch/n27 }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,pip_flush}),
    .c({addr_if[28],\ins_fetch/n1 [26]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4651_o,addr_if[28]}),
    .mi({open_n26533,addr_if[28]}),
    .sr(rst_pad),
    .f({_al_u4652_o,_al_u9551_o}),
    .q({open_n26548,\biu/cache_ctrl_logic/l1i_va [28]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4653|biu/cache_ctrl_logic/reg3_b28  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,open_n26549}),
    .b({_al_u3950_o,\biu/cache_ctrl_logic/l1i_va [28]}),
    .c({\biu/cache_ctrl_logic/l1i_pa [92],addr_ex[28]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[28],_al_u6410_o}),
    .mi({open_n26553,addr_ex[28]}),
    .sr(rst_pad),
    .f({_al_u4653_o,_al_u6411_o}),
    .q({open_n26568,\biu/cache_ctrl_logic/l1d_va [28]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4655|biu/cache_ctrl_logic/reg1_b92  (
    .a({open_n26569,_al_u3945_o}),
    .b({_al_u4653_o,_al_u3947_o}),
    .c({_al_u4654_o,\biu/cache_ctrl_logic/l1d_pa [92]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4652_o,\biu/cache_ctrl_logic/pa_temp [92]}),
    .mi({open_n26580,\biu/cache_ctrl_logic/pa_temp [92]}),
    .sr(rst_pad),
    .f({_al_u4655_o,_al_u4654_o}),
    .q({open_n26584,\biu/cache_ctrl_logic/l1i_pa [92]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u4657|_al_u4597  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4399_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/n209 [27],\biu/cache_ctrl_logic/n209 [36]}),
    .d({addr_ex[27],addr_ex[36]}),
    .f({_al_u4657_o,_al_u4597_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4658|_al_u4718  (
    .b({\biu/bus_unit/mmu/n19_lutinv ,\biu/bus_unit/mmu/n19_lutinv }),
    .c({addr_if[27],addr_if[17]}),
    .d({_al_u4657_o,_al_u4717_o}),
    .f({_al_u4658_o,_al_u4718_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4661|biu/cache_ctrl_logic/reg1_b91  (
    .a({open_n26631,_al_u3945_o}),
    .b({_al_u4659_o,_al_u3947_o}),
    .c({_al_u4660_o,\biu/cache_ctrl_logic/l1d_pa [91]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4658_o,\biu/cache_ctrl_logic/pa_temp [91]}),
    .mi({open_n26635,\biu/cache_ctrl_logic/pa_temp [91]}),
    .sr(rst_pad),
    .f({_al_u4661_o,_al_u4660_o}),
    .q({open_n26650,\biu/cache_ctrl_logic/l1i_pa [91]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4664|biu/cache_ctrl_logic/reg1_b90  (
    .a({open_n26651,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[26],\biu/cache_ctrl_logic/l1d_pa [90]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4663_o,\biu/cache_ctrl_logic/pa_temp [90]}),
    .mi({open_n26655,\biu/cache_ctrl_logic/pa_temp [90]}),
    .sr(rst_pad),
    .f({_al_u4664_o,_al_u4663_o}),
    .q({open_n26670,\biu/cache_ctrl_logic/l1i_pa [90]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4667|_al_u4665  (
    .a({open_n26671,_al_u3950_o}),
    .b({_al_u4665_o,_al_u4399_o}),
    .c({_al_u4666_o,\biu/cache_ctrl_logic/n209 [26]}),
    .d({_al_u4664_o,\biu/cache_ctrl_logic/l1i_pa [90]}),
    .f({_al_u4667_o,_al_u4665_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4670|biu/cache_ctrl_logic/reg1_b89  (
    .a({open_n26696,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[25],\biu/cache_ctrl_logic/l1d_pa [89]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4669_o,\biu/cache_ctrl_logic/pa_temp [89]}),
    .mi({open_n26707,\biu/cache_ctrl_logic/pa_temp [89]}),
    .sr(rst_pad),
    .f({_al_u4670_o,_al_u4669_o}),
    .q({open_n26711,\biu/cache_ctrl_logic/l1i_pa [89]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4673|_al_u4671  (
    .a({open_n26712,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4671_o,_al_u3950_o}),
    .c({_al_u4672_o,\biu/cache_ctrl_logic/l1i_pa [89]}),
    .d({_al_u4670_o,addr_ex[25]}),
    .f({_al_u4673_o,_al_u4671_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4675|biu/cache_ctrl_logic/reg1_b88  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n212 [24],\biu/cache_ctrl_logic/pa_temp [88]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [88],addr_ex[24]}),
    .mi({open_n26740,\biu/cache_ctrl_logic/pa_temp [88]}),
    .sr(rst_pad),
    .f({_al_u4675_o,_al_u4678_o}),
    .q({open_n26755,\biu/cache_ctrl_logic/l1i_pa [88]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4676|ins_fetch/reg0_b24  (
    .a({open_n26756,\biu/cache_ctrl_logic/l1i_va [24]}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,\biu/cache_ctrl_logic/l1i_va [58]}),
    .c({addr_if[24],addr_if[24]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4675_o,addr_if[58]}),
    .mi({open_n26767,addr_if[24]}),
    .sr(rst_pad),
    .f({_al_u4676_o,_al_u9208_o}),
    .q({open_n26771,id_ins_pc[24]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4679|biu/cache_ctrl_logic/reg4_b88  (
    .a({open_n26772,_al_u3947_o}),
    .b({_al_u4677_o,_al_u4399_o}),
    .c({_al_u4678_o,\biu/cache_ctrl_logic/n209 [24]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4676_o,\biu/cache_ctrl_logic/l1d_pa [88]}),
    .mi({open_n26783,\biu/cache_ctrl_logic/pa_temp [88]}),
    .sr(rst_pad),
    .f({_al_u4679_o,_al_u4677_o}),
    .q({open_n26787,\biu/cache_ctrl_logic/l1d_pa [88]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4682|exu/reg3_b23  (
    .a({open_n26788,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3950_o}),
    .c({addr_if[23],\biu/cache_ctrl_logic/l1i_pa [87]}),
    .clk(clk_pad),
    .d({_al_u4681_o,addr_ex[23]}),
    .mi({open_n26793,addr_ex[23]}),
    .sr(rst_pad),
    .f({_al_u4682_o,_al_u4681_o}),
    .q({open_n26808,new_pc[23]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4685|biu/cache_ctrl_logic/reg1_b87  (
    .a({open_n26809,_al_u3945_o}),
    .b({_al_u4683_o,_al_u3947_o}),
    .c({_al_u4684_o,\biu/cache_ctrl_logic/l1d_pa [87]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4682_o,\biu/cache_ctrl_logic/pa_temp [87]}),
    .mi({open_n26820,\biu/cache_ctrl_logic/pa_temp [87]}),
    .sr(rst_pad),
    .f({_al_u4685_o,_al_u4684_o}),
    .q({open_n26824,\biu/cache_ctrl_logic/l1i_pa [87]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4688|ins_fetch/reg0_b22  (
    .a({open_n26825,\biu/cache_ctrl_logic/l1i_va [22]}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,\biu/cache_ctrl_logic/l1i_va [48]}),
    .c({addr_if[22],addr_if[22]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4687_o,addr_if[48]}),
    .mi({open_n26836,addr_if[22]}),
    .sr(rst_pad),
    .f({_al_u4688_o,_al_u9225_o}),
    .q({open_n26840,id_ins_pc[22]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4691|biu/cache_ctrl_logic/reg1_b86  (
    .a({open_n26841,_al_u3945_o}),
    .b({_al_u4689_o,_al_u3947_o}),
    .c({_al_u4690_o,\biu/cache_ctrl_logic/l1d_pa [86]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4688_o,\biu/cache_ctrl_logic/pa_temp [86]}),
    .mi({open_n26845,\biu/cache_ctrl_logic/pa_temp [86]}),
    .sr(rst_pad),
    .f({_al_u4691_o,_al_u4690_o}),
    .q({open_n26860,\biu/cache_ctrl_logic/l1i_pa [86]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4693|biu/cache_ctrl_logic/reg1_b85  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n212 [21],\biu/cache_ctrl_logic/pa_temp [85]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [85],addr_ex[21]}),
    .mi({open_n26871,\biu/cache_ctrl_logic/pa_temp [85]}),
    .sr(rst_pad),
    .f({_al_u4693_o,_al_u4696_o}),
    .q({open_n26875,\biu/cache_ctrl_logic/l1i_pa [85]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4697|biu/cache_ctrl_logic/reg4_b85  (
    .a({open_n26876,_al_u3947_o}),
    .b({_al_u4695_o,_al_u4399_o}),
    .c({_al_u4696_o,\biu/cache_ctrl_logic/n209 [21]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4694_o,\biu/cache_ctrl_logic/l1d_pa [85]}),
    .mi({open_n26880,\biu/cache_ctrl_logic/pa_temp [85]}),
    .sr(rst_pad),
    .f({_al_u4697_o,_al_u4695_o}),
    .q({open_n26895,\biu/cache_ctrl_logic/l1d_pa [85]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4700|_al_u4699  (
    .a({open_n26896,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3950_o}),
    .c({addr_if[20],\biu/cache_ctrl_logic/n212 [20]}),
    .d({_al_u4699_o,\biu/cache_ctrl_logic/l1i_pa [84]}),
    .f({_al_u4700_o,_al_u4699_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4703|biu/cache_ctrl_logic/reg1_b84  (
    .a({open_n26917,_al_u3945_o}),
    .b({_al_u4701_o,_al_u3947_o}),
    .c({_al_u4702_o,\biu/cache_ctrl_logic/l1d_pa [84]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4700_o,\biu/cache_ctrl_logic/pa_temp [84]}),
    .mi({open_n26921,\biu/cache_ctrl_logic/pa_temp [84]}),
    .sr(rst_pad),
    .f({_al_u4703_o,_al_u4702_o}),
    .q({open_n26936,\biu/cache_ctrl_logic/l1i_pa [84]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4706|_al_u4705  (
    .a({open_n26937,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u4399_o}),
    .c({addr_if[19],\biu/cache_ctrl_logic/n209 [19]}),
    .d({_al_u4705_o,addr_ex[19]}),
    .f({_al_u4706_o,_al_u4705_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4709|biu/cache_ctrl_logic/reg4_b83  (
    .a({open_n26962,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4707_o,_al_u3947_o}),
    .c({_al_u4708_o,\biu/cache_ctrl_logic/n212 [19]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4706_o,\biu/cache_ctrl_logic/l1d_pa [83]}),
    .mi({open_n26966,\biu/cache_ctrl_logic/pa_temp [83]}),
    .sr(rst_pad),
    .f({_al_u4709_o,_al_u4707_o}),
    .q({open_n26981,\biu/cache_ctrl_logic/l1d_pa [83]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4712|_al_u4711  (
    .a({open_n26982,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3950_o}),
    .c({addr_if[18],\biu/cache_ctrl_logic/l1i_pa [82]}),
    .d({_al_u4711_o,addr_ex[18]}),
    .f({_al_u4712_o,_al_u4711_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4715|biu/cache_ctrl_logic/reg1_b82  (
    .a({open_n27003,_al_u3945_o}),
    .b({_al_u4713_o,_al_u3947_o}),
    .c({_al_u4714_o,\biu/cache_ctrl_logic/l1d_pa [82]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4712_o,\biu/cache_ctrl_logic/pa_temp [82]}),
    .mi({open_n27014,\biu/cache_ctrl_logic/pa_temp [82]}),
    .sr(rst_pad),
    .f({_al_u4715_o,_al_u4714_o}),
    .q({open_n27018,\biu/cache_ctrl_logic/l1i_pa [82]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4717|biu/cache_ctrl_logic/reg1_b81  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n212 [17],\biu/cache_ctrl_logic/pa_temp [81]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [81],addr_ex[17]}),
    .mi({open_n27029,\biu/cache_ctrl_logic/pa_temp [81]}),
    .sr(rst_pad),
    .f({_al_u4717_o,_al_u4720_o}),
    .q({open_n27033,\biu/cache_ctrl_logic/l1i_pa [81]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4721|biu/cache_ctrl_logic/reg4_b81  (
    .a({open_n27034,_al_u3947_o}),
    .b({_al_u4719_o,_al_u4399_o}),
    .c({_al_u4720_o,\biu/cache_ctrl_logic/n209 [17]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4718_o,\biu/cache_ctrl_logic/l1d_pa [81]}),
    .mi({open_n27045,\biu/cache_ctrl_logic/pa_temp [81]}),
    .sr(rst_pad),
    .f({_al_u4721_o,_al_u4719_o}),
    .q({open_n27049,\biu/cache_ctrl_logic/l1d_pa [81]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4723|biu/cache_ctrl_logic/reg1_b80  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n212 [16],\biu/cache_ctrl_logic/pa_temp [80]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [80],addr_ex[16]}),
    .mi({open_n27053,\biu/cache_ctrl_logic/pa_temp [80]}),
    .sr(rst_pad),
    .f({_al_u4723_o,_al_u4726_o}),
    .q({open_n27068,\biu/cache_ctrl_logic/l1i_pa [80]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D@C))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000001000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4724|biu/cache_ctrl_logic/reg3_b16  (
    .a({open_n27069,_al_u6389_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u6390_o}),
    .c({addr_if[16],\biu/cache_ctrl_logic/l1i_va [16]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4723_o,addr_ex[16]}),
    .mi({open_n27080,addr_ex[16]}),
    .sr(rst_pad),
    .f({_al_u4724_o,_al_u6391_o}),
    .q({open_n27084,\biu/cache_ctrl_logic/l1d_va [16]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4727|biu/cache_ctrl_logic/reg4_b80  (
    .a({open_n27085,_al_u3947_o}),
    .b({_al_u4725_o,_al_u4399_o}),
    .c({_al_u4726_o,\biu/cache_ctrl_logic/n209 [16]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4724_o,\biu/cache_ctrl_logic/l1d_pa [80]}),
    .mi({open_n27096,\biu/cache_ctrl_logic/pa_temp [80]}),
    .sr(rst_pad),
    .f({_al_u4727_o,_al_u4725_o}),
    .q({open_n27100,\biu/cache_ctrl_logic/l1d_pa [80]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4730|biu/cache_ctrl_logic/reg1_b79  (
    .a({open_n27101,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[15],\biu/cache_ctrl_logic/l1d_pa [79]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4729_o,\biu/cache_ctrl_logic/pa_temp [79]}),
    .mi({open_n27112,\biu/cache_ctrl_logic/pa_temp [79]}),
    .sr(rst_pad),
    .f({_al_u4730_o,_al_u4729_o}),
    .q({open_n27116,\biu/cache_ctrl_logic/l1i_pa [79]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u4733|_al_u4731  (
    .a({open_n27117,_al_u3950_o}),
    .b({_al_u4731_o,_al_u4399_o}),
    .c({_al_u4732_o,\biu/cache_ctrl_logic/n209 [15]}),
    .d({_al_u4730_o,\biu/cache_ctrl_logic/l1i_pa [79]}),
    .f({_al_u4733_o,_al_u4731_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4736|biu/cache_ctrl_logic/reg1_b78  (
    .a({open_n27138,_al_u3945_o}),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .c({addr_if[14],\biu/cache_ctrl_logic/l1d_pa [78]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4735_o,\biu/cache_ctrl_logic/pa_temp [78]}),
    .mi({open_n27142,\biu/cache_ctrl_logic/pa_temp [78]}),
    .sr(rst_pad),
    .f({_al_u4736_o,_al_u4735_o}),
    .q({open_n27157,\biu/cache_ctrl_logic/l1i_pa [78]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4738|biu/cache_ctrl_logic/reg3_b14  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/l1i_va [14]}),
    .b({_al_u4399_o,\biu/cache_ctrl_logic/l1i_va [22]}),
    .c({\biu/cache_ctrl_logic/n209 [14],addr_ex[14]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[14],addr_ex[22]}),
    .mi({open_n27161,addr_ex[14]}),
    .sr(rst_pad),
    .f({_al_u4738_o,_al_u6392_o}),
    .q({open_n27176,\biu/cache_ctrl_logic/l1d_va [14]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4739|_al_u4737  (
    .a({open_n27177,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4737_o,_al_u3950_o}),
    .c({_al_u4738_o,\biu/cache_ctrl_logic/n212 [14]}),
    .d({_al_u4736_o,\biu/cache_ctrl_logic/l1i_pa [78]}),
    .f({_al_u4739_o,_al_u4737_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4741|biu/cache_ctrl_logic/reg1_b77  (
    .a({_al_u3950_o,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4399_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n209 [13],\biu/cache_ctrl_logic/n212 [13]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [77],\biu/cache_ctrl_logic/pa_temp [77]}),
    .mi({open_n27205,\biu/cache_ctrl_logic/pa_temp [77]}),
    .sr(rst_pad),
    .f({_al_u4741_o,_al_u4744_o}),
    .q({open_n27220,\biu/cache_ctrl_logic/l1i_pa [77]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4745|biu/cache_ctrl_logic/reg4_b77  (
    .a({open_n27221,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4743_o,_al_u3947_o}),
    .c({_al_u4744_o,\biu/cache_ctrl_logic/l1d_pa [77]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4742_o,addr_ex[13]}),
    .mi({open_n27225,\biu/cache_ctrl_logic/pa_temp [77]}),
    .sr(rst_pad),
    .f({_al_u4745_o,_al_u4743_o}),
    .q({open_n27240,\biu/cache_ctrl_logic/l1d_pa [77]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4748|_al_u4747  (
    .a({open_n27241,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({\biu/bus_unit/mmu/n19_lutinv ,_al_u4399_o}),
    .c({addr_if[12],\biu/cache_ctrl_logic/n209 [12]}),
    .d({_al_u4747_o,\biu/cache_ctrl_logic/n212 [12]}),
    .f({_al_u4748_o,_al_u4747_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4751|biu/cache_ctrl_logic/reg4_b76  (
    .a({open_n27262,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u4749_o,_al_u3947_o}),
    .c({_al_u4750_o,\biu/cache_ctrl_logic/l1d_pa [76]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4748_o,addr_ex[12]}),
    .mi({open_n27273,\biu/cache_ctrl_logic/pa_temp [76]}),
    .sr(rst_pad),
    .f({_al_u4751_o,_al_u4749_o}),
    .q({open_n27277,\biu/cache_ctrl_logic/l1d_pa [76]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4753|biu/cache_ctrl_logic/reg1_b75  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/n212 [11],\biu/cache_ctrl_logic/pa_temp [75]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pa [75],addr_ex[11]}),
    .mi({open_n27281,\biu/cache_ctrl_logic/pa_temp [75]}),
    .sr(rst_pad),
    .f({_al_u4753_o,_al_u4756_o}),
    .q({open_n27296,\biu/cache_ctrl_logic/l1i_pa [75]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4754|_al_u4694  (
    .b({\biu/bus_unit/mmu/n19_lutinv ,\biu/bus_unit/mmu/n19_lutinv }),
    .c({addr_if[11],addr_if[21]}),
    .d({_al_u4753_o,_al_u4693_o}),
    .f({_al_u4754_o,_al_u4694_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4757|biu/cache_ctrl_logic/reg4_b75  (
    .a({open_n27319,_al_u3947_o}),
    .b({_al_u4755_o,_al_u4399_o}),
    .c({_al_u4756_o,\biu/cache_ctrl_logic/n209 [11]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4754_o,\biu/cache_ctrl_logic/l1d_pa [75]}),
    .mi({open_n27323,\biu/cache_ctrl_logic/pa_temp [75]}),
    .sr(rst_pad),
    .f({_al_u4757_o,_al_u4755_o}),
    .q({open_n27338,\biu/cache_ctrl_logic/l1d_pa [75]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4760|ins_fetch/reg0_b10  (
    .b({\biu/bus_unit/mmu/n19_lutinv ,open_n27341}),
    .c({addr_if[10],1'b0}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u4759_o,if_hold}),
    .mi({open_n27345,addr_if[10]}),
    .sr(rst_pad),
    .f({_al_u4760_o,\ins_fetch/n9 }),
    .q({open_n27360,id_ins_pc[10]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4761|biu/cache_ctrl_logic/reg1_b74  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3947_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [74],\biu/cache_ctrl_logic/l1d_pa [74]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({addr_ex[10],\biu/cache_ctrl_logic/pa_temp [74]}),
    .mi({open_n27364,\biu/cache_ctrl_logic/pa_temp [74]}),
    .sr(rst_pad),
    .f({_al_u4761_o,_al_u4759_o}),
    .q({open_n27379,\biu/cache_ctrl_logic/l1i_pa [74]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4763|_al_u4762  (
    .a({open_n27380,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u4761_o,_al_u4399_o}),
    .c({_al_u4762_o,\biu/cache_ctrl_logic/n209 [10]}),
    .d({_al_u4760_o,\biu/cache_ctrl_logic/n212 [10]}),
    .f({_al_u4763_o,_al_u4762_o}));
  // ../../RTL/CPU/BIU/bus_unit.v(163)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~D)"),
    //.LUTF1("(~(D*~B)*~(C)*~(A)+~(D*~B)*C*~(A)+~(~(D*~B))*C*A+~(D*~B)*C*A)"),
    //.LUTG0("~(C*~D)"),
    //.LUTG1("(~(D*~B)*~(C)*~(A)+~(D*~B)*C*~(A)+~(~(D*~B))*C*A+~(D*~B)*C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100001111),
    .INIT_LUTF1(16'b1110010011110101),
    .INIT_LUTG0(16'b1111111100001111),
    .INIT_LUTG1(16'b1110010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4766|biu/bus_unit/reg1_b2  (
    .a({_al_u3404_o,open_n27405}),
    .b({_al_u3407_o,open_n27406}),
    .c({_al_u4099_o,_al_u4766_o}),
    .clk(clk_pad),
    .d({\biu/bus_unit/statu [2],_al_u4765_o}),
    .sr(rst_pad),
    .f({_al_u4766_o,open_n27424}),
    .q({open_n27428,\biu/bus_unit/statu [2]}));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*~B)*~(D)*~(A)+~(~C*~B)*D*~(A)+~(~(~C*~B))*D*A+~(~C*~B)*D*A)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(~C*~B)*~(D)*~(A)+~(~C*~B)*D*~(A)+~(~(~C*~B))*D*A+~(~C*~B)*D*A)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111001010100),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111111001010100),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4768|biu/cache_ctrl_logic/reg5_b7  (
    .a({_al_u3945_o,\biu/cache_ctrl_logic/n149 }),
    .b({_al_u3947_o,_al_u3947_o}),
    .c({\biu/cache_ctrl_logic/l1d_pte [7],\biu/cache_ctrl_logic/l1d_pte [7]}),
    .clk(clk_pad),
    .d(2'b00),
    .sr(rst_pad),
    .f({_al_u4768_o,open_n27446}),
    .q({open_n27450,\biu/cache_ctrl_logic/l1d_pte [7]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*~B)*~(D)*~(A)+~(~C*~B)*D*~(A)+~(~(~C*~B))*D*A+~(~C*~B)*D*A)"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(~(~C*~B)*~(D)*~(A)+~(~C*~B)*D*~(A)+~(~(~C*~B))*D*A+~(~C*~B)*D*A)"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111001010100),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b1111111001010100),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4769|biu/cache_ctrl_logic/reg2_b7  (
    .a({_al_u2705_o,\biu/cache_ctrl_logic/n135 }),
    .b({_al_u4768_o,_al_u3950_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1i_pte [7]}),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [7],1'b0}),
    .sr(rst_pad),
    .f({_al_u4769_o,open_n27468}),
    .q({open_n27472,\biu/cache_ctrl_logic/l1i_pte [7]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(~C*D))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4770|_al_u5747  (
    .b({_al_u4769_o,_al_u2705_o}),
    .c({_al_u3222_o,\biu/bus_unit/mmu_hwdata [46]}),
    .d({\exu/lsu/n1 [7],_al_u5746_o}),
    .f({_al_u4770_o,hwdata_pad[46]}));
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4771|biu/bus_unit/mmu/reg3_b7  (
    .a({open_n27499,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [7],\biu/bus_unit/mmu_hwdata [7]}),
    .clk(clk_pad),
    .d({_al_u4770_o,hrdata_pad[7]}),
    .sr(rst_pad),
    .f({hwdata_pad[7],open_n27517}),
    .q({open_n27521,\biu/bus_unit/mmu_hwdata [7]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4774|biu/cache_ctrl_logic/reg2_b6  (
    .a({open_n27522,_al_u2705_o}),
    .b({_al_u4773_o,_al_u4772_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\exu/lsu/n1 [6],\biu/cache_ctrl_logic/pte_temp [6]}),
    .mi({open_n27533,\biu/cache_ctrl_logic/pte_temp [6]}),
    .sr(rst_pad),
    .f({_al_u4774_o,_al_u4773_o}),
    .q({open_n27537,\biu/cache_ctrl_logic/l1i_pte [6]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4778|biu/cache_ctrl_logic/reg2_b5  (
    .a({open_n27538,_al_u2705_o}),
    .b({_al_u4777_o,_al_u4776_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\exu/lsu/n1 [5],\biu/cache_ctrl_logic/pte_temp [5]}),
    .mi({open_n27549,\biu/cache_ctrl_logic/pte_temp [5]}),
    .sr(rst_pad),
    .f({_al_u4778_o,_al_u4777_o}),
    .q({open_n27553,\biu/cache_ctrl_logic/l1i_pte [5]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4779|biu/bus_unit/mmu/reg3_b5  (
    .a({open_n27554,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [5],\biu/bus_unit/mmu_hwdata [5]}),
    .clk(clk_pad),
    .d({_al_u4778_o,hrdata_pad[5]}),
    .sr(rst_pad),
    .f({hwdata_pad[5],open_n27568}),
    .q({open_n27572,\biu/bus_unit/mmu_hwdata [5]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4780|biu/cache_ctrl_logic/reg2_b4  (
    .a({_al_u3947_o,_al_u2705_o}),
    .b({_al_u3950_o,_al_u4780_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [4],_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [4],\biu/cache_ctrl_logic/pte_temp [4]}),
    .mi({open_n27583,\biu/cache_ctrl_logic/pte_temp [4]}),
    .sr(rst_pad),
    .f({_al_u4780_o,_al_u4781_o}),
    .q({open_n27587,\biu/cache_ctrl_logic/l1i_pte [4]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u4782|_al_u5735  (
    .b({_al_u4781_o,_al_u2705_o}),
    .c({_al_u3222_o,\biu/bus_unit/mmu_hwdata [49]}),
    .d({\exu/lsu/n1 [4],_al_u5734_o}),
    .f({_al_u4782_o,hwdata_pad[49]}));
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4783|biu/bus_unit/mmu/reg3_b4  (
    .a({open_n27610,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [4],\biu/bus_unit/mmu_hwdata [4]}),
    .clk(clk_pad),
    .d({_al_u4782_o,hrdata_pad[4]}),
    .sr(rst_pad),
    .f({hwdata_pad[4],open_n27624}),
    .q({open_n27628,\biu/bus_unit/mmu_hwdata [4]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4784|biu/cache_ctrl_logic/reg2_b3  (
    .a({_al_u3947_o,_al_u2705_o}),
    .b({_al_u3950_o,_al_u4784_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [3],_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [3],\biu/cache_ctrl_logic/pte_temp [3]}),
    .mi({open_n27632,\biu/cache_ctrl_logic/pte_temp [3]}),
    .sr(rst_pad),
    .f({_al_u4784_o,_al_u4785_o}),
    .q({open_n27647,\biu/cache_ctrl_logic/l1i_pte [3]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(~C*D))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4786|_al_u4787  (
    .b({_al_u4785_o,_al_u2705_o}),
    .c({_al_u3222_o,\biu/bus_unit/mmu_hwdata [3]}),
    .d({\exu/lsu/n1 [3],_al_u4786_o}),
    .f({_al_u4786_o,hwdata_pad[3]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4788|biu/cache_ctrl_logic/reg2_b2  (
    .a({_al_u3947_o,_al_u2705_o}),
    .b({_al_u3950_o,_al_u4788_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [2],_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [2],\biu/cache_ctrl_logic/pte_temp [2]}),
    .mi({open_n27684,\biu/cache_ctrl_logic/pte_temp [2]}),
    .sr(rst_pad),
    .f({_al_u4788_o,_al_u4789_o}),
    .q({open_n27688,\biu/cache_ctrl_logic/l1i_pte [2]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u4790|_al_u4791  (
    .b({_al_u4789_o,_al_u2705_o}),
    .c({_al_u3222_o,\biu/bus_unit/mmu_hwdata [2]}),
    .d({\exu/lsu/n1 [2],_al_u4790_o}),
    .f({_al_u4790_o,hwdata_pad[2]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4792|biu/cache_ctrl_logic/reg2_b1  (
    .a({_al_u3947_o,_al_u2705_o}),
    .b({_al_u3950_o,_al_u4792_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [1],_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [1],\biu/cache_ctrl_logic/pte_temp [1]}),
    .mi({open_n27714,\biu/cache_ctrl_logic/pte_temp [1]}),
    .sr(rst_pad),
    .f({_al_u4792_o,_al_u4793_o}),
    .q({open_n27729,\biu/cache_ctrl_logic/l1i_pte [1]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(~C*D))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4794|_al_u5723  (
    .b({_al_u4793_o,_al_u2705_o}),
    .c({_al_u3222_o,\biu/bus_unit/mmu_hwdata [52]}),
    .d({\exu/lsu/n1 [1],_al_u5722_o}),
    .f({_al_u4794_o,hwdata_pad[52]}));
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4795|biu/bus_unit/mmu/reg3_b1  (
    .a({open_n27756,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [1],\biu/bus_unit/mmu_hwdata [1]}),
    .clk(clk_pad),
    .d({_al_u4794_o,hrdata_pad[1]}),
    .sr(rst_pad),
    .f({hwdata_pad[1],open_n27770}),
    .q({open_n27774,\biu/bus_unit/mmu_hwdata [1]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(B*~(~C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4798|biu/cache_ctrl_logic/reg5_b0  (
    .b({_al_u4797_o,_al_u3947_o}),
    .c({_al_u3222_o,\biu/cache_ctrl_logic/l1d_pte [0]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\exu/lsu/n1 [0],_al_u4796_o}),
    .mi({open_n27780,\biu/cache_ctrl_logic/pte_temp [0]}),
    .sr(rst_pad),
    .f({_al_u4798_o,_al_u4797_o}),
    .q({open_n27795,\biu/cache_ctrl_logic/l1d_pte [0]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(C)*~(B)+~D*C*~(B)+~(~D)*C*B+~D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b1100000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b1100000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4799|biu/bus_unit/mmu/reg3_b0  (
    .a({open_n27796,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [0],\biu/bus_unit/mmu_hwdata [0]}),
    .clk(clk_pad),
    .d({_al_u4798_o,hrdata_pad[0]}),
    .sr(rst_pad),
    .f({hwdata_pad[0],open_n27814}),
    .q({open_n27818,\biu/bus_unit/mmu_hwdata [0]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~A*~(D*~(~C*~B)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000101010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4802|ins_dec/rd_data_sub_reg  (
    .a({\ins_dec/ins_srli ,open_n27819}),
    .b({\ins_dec/funct7_0_lutinv ,\ins_dec/funct7_32_lutinv }),
    .c({\ins_dec/funct7_32_lutinv ,_al_u3925_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4801_o,\ins_dec/funct3_0_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u4802_o,open_n27832}),
    .q({open_n27836,rd_data_sub}));  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*~C*B*~A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*~C*B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000010000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000010000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4804|ins_dec/reg10_b26  (
    .a({id_ins[26],open_n27837}),
    .b({_al_u3216_o,open_n27838}),
    .c({_al_u3217_o,id_ins[26]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3384_o,id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u4804_o,open_n27855}),
    .q({open_n27859,ex_exc_code[26]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u4806|_al_u4803  (
    .a({open_n27860,\ins_dec/op_32_imm_lutinv }),
    .b({\ins_dec/ins_srai ,_al_u3216_o}),
    .c({\ins_dec/funct7_32_lutinv ,_al_u3217_o}),
    .d({\ins_dec/n38 ,_al_u3384_o}),
    .f({_al_u4806_o,\ins_dec/n38 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4809|_al_u4808  (
    .a({open_n27881,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u3950_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [66],\biu/cache_ctrl_logic/n209 [2]}),
    .d({_al_u4808_o,\biu/cache_ctrl_logic/n212 [2]}),
    .f({_al_u4809_o,_al_u4808_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4811|biu/cache_ctrl_logic/reg1_b66  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u4810_o,_al_u3947_o}),
    .c({\biu/cache_ctrl_logic/n75_lutinv ,\biu/cache_ctrl_logic/l1d_pa [66]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({addr_ex[2],\biu/cache_ctrl_logic/pa_temp [66]}),
    .mi({open_n27909,\biu/cache_ctrl_logic/pa_temp [66]}),
    .sr(rst_pad),
    .f({_al_u4811_o,_al_u4810_o}),
    .q({open_n27924,\biu/cache_ctrl_logic/l1i_pa [66]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4813|biu/cache_ctrl_logic/reg6_b66  (
    .b({_al_u4403_o,_al_u2705_o}),
    .c({\biu/cache_ctrl_logic/n207 [2],\biu/paddress [66]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4812_o,_al_u4813_o}),
    .mi({open_n27937,\biu/paddress [66]}),
    .sr(rst_pad),
    .f({_al_u4813_o,haddr_pad[2]}),
    .q({open_n27941,\biu/cache_ctrl_logic/pa_temp [66]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u4816|_al_u4815  (
    .a({open_n27942,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({_al_u3950_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [65],\biu/cache_ctrl_logic/n209 [1]}),
    .d({_al_u4815_o,addr_ex[1]}),
    .f({_al_u4816_o,_al_u4815_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4818|biu/cache_ctrl_logic/reg1_b65  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u4817_o,_al_u3947_o}),
    .c({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/l1d_pa [65]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/n212 [1],\biu/cache_ctrl_logic/pa_temp [65]}),
    .mi({open_n27973,\biu/cache_ctrl_logic/pa_temp [65]}),
    .sr(rst_pad),
    .f({_al_u4818_o,_al_u4817_o}),
    .q({open_n27977,\biu/cache_ctrl_logic/l1i_pa [65]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000100000001),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4819|ins_fetch/reg2_b1  (
    .a({_al_u4816_o,_al_u6733_o}),
    .b({_al_u4818_o,_al_u6734_o}),
    .c({\biu/bus_unit/mmu/n19_lutinv ,\cu_ru/m_s_status/n2 }),
    .ce(pip_flush),
    .clk(clk_pad),
    .d({addr_if[1],\cu_ru/mepc [1]}),
    .sr(rst_pad),
    .f({_al_u4819_o,open_n27990}),
    .q({open_n27994,addr_if[1]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4820|biu/cache_ctrl_logic/reg6_b65  (
    .b({_al_u4403_o,_al_u2705_o}),
    .c({\biu/cache_ctrl_logic/n207 [1],\biu/paddress [65]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4819_o,_al_u4820_o}),
    .mi({open_n28000,\biu/paddress [65]}),
    .sr(rst_pad),
    .f({_al_u4820_o,haddr_pad[1]}),
    .q({open_n28015,\biu/cache_ctrl_logic/pa_temp [65]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4823|biu/cache_ctrl_logic/reg1_b64  (
    .a({open_n28016,\biu/cache_ctrl_logic/n97_lutinv }),
    .b({_al_u3950_o,_al_u3945_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [64],\biu/cache_ctrl_logic/n212 [0]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({_al_u4822_o,\biu/cache_ctrl_logic/pa_temp [64]}),
    .mi({open_n28020,\biu/cache_ctrl_logic/pa_temp [64]}),
    .sr(rst_pad),
    .f({_al_u4823_o,_al_u4824_o}),
    .q({open_n28035,\biu/cache_ctrl_logic/l1i_pa [64]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4826|biu/cache_ctrl_logic/reg4_b64  (
    .a({_al_u4823_o,_al_u2705_o}),
    .b({_al_u4825_o,_al_u4824_o}),
    .c({\biu/bus_unit/mmu/n19_lutinv ,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_if[0],\biu/cache_ctrl_logic/l1d_pa [64]}),
    .mi({open_n28039,\biu/cache_ctrl_logic/pa_temp [64]}),
    .sr(rst_pad),
    .f({_al_u4826_o,_al_u4825_o}),
    .q({open_n28054,\biu/cache_ctrl_logic/l1d_pa [64]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4827|biu/cache_ctrl_logic/reg6_b64  (
    .b({_al_u4403_o,_al_u2705_o}),
    .c({\biu/cache_ctrl_logic/n207 [0],\biu/paddress [64]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u4826_o,_al_u4827_o}),
    .mi({open_n28060,\biu/paddress [64]}),
    .sr(rst_pad),
    .f({_al_u4827_o,haddr_pad[0]}),
    .q({open_n28075,\biu/cache_ctrl_logic/pa_temp [64]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~C*~B))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(A*~(D*~C*~B))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b1010100010101010),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b1010100010101010),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4829|_al_u4830  (
    .a({open_n28076,_al_u4829_o}),
    .b({_al_u3404_o,_al_u2890_o}),
    .c({_al_u4099_o,_al_u3407_o}),
    .d({_al_u2890_o,\biu/bus_unit/statu [1]}),
    .f({_al_u4829_o,_al_u4830_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A*~(~D*C))"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b0001000100000001),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u4832|_al_u4831  (
    .a({open_n28101,_al_u4830_o}),
    .b({_al_u3403_o,_al_u3403_o}),
    .c({_al_u4099_o,_al_u3404_o}),
    .d({_al_u4831_o,hresp_pad}),
    .f({_al_u4832_o,_al_u4831_o}));
  // ../../RTL/CPU/BIU/bus_unit.v(163)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(~C*B))"),
    //.LUT1("(~D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011111111),
    .INIT_LUT1(16'b0000000011001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4835|biu/bus_unit/reg1_b1  (
    .b({_al_u2847_o,_al_u4194_o}),
    .c({_al_u3944_o,_al_u4835_o}),
    .clk(clk_pad),
    .d({_al_u4834_o,_al_u4833_o}),
    .sr(rst_pad),
    .f({_al_u4835_o,open_n28137}),
    .q({open_n28141,\biu/bus_unit/statu [1]}));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(D*~(C*B*A))"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0111111100000000),
    .MODE("LOGIC"))
    \_al_u4839|_al_u4838  (
    .a({_al_u4134_o,open_n28142}),
    .b({_al_u4136_o,1'b0}),
    .c({_al_u4838_o,1'b0}),
    .d({wb_valid,_al_u4837_o}),
    .f({ex_nop,_al_u4838_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4842|biu/cache_ctrl_logic/reg2_b15  (
    .a({open_n28163,_al_u2705_o}),
    .b({_al_u4841_o,_al_u4840_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [15],\biu/cache_ctrl_logic/pte_temp [15]}),
    .mi({open_n28174,\biu/cache_ctrl_logic/pte_temp [15]}),
    .sr(rst_pad),
    .f({_al_u4842_o,_al_u4841_o}),
    .q({open_n28178,\biu/cache_ctrl_logic/l1i_pte [15]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4843|biu/bus_unit/mmu/reg3_b15  (
    .a({open_n28179,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [15],\biu/bus_unit/mmu_hwdata [15]}),
    .clk(clk_pad),
    .d({_al_u4842_o,hrdata_pad[15]}),
    .sr(rst_pad),
    .f({hwdata_pad[15],open_n28197}),
    .q({open_n28201,\biu/bus_unit/mmu_hwdata [15]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4845|biu/cache_ctrl_logic/reg2_b14  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u4844_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [14]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [14],\biu/cache_ctrl_logic/pte_temp [14]}),
    .mi({open_n28205,\biu/cache_ctrl_logic/pte_temp [14]}),
    .sr(rst_pad),
    .f({_al_u4845_o,_al_u4844_o}),
    .q({open_n28220,\biu/cache_ctrl_logic/l1i_pte [14]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u4846|_al_u5806  (
    .b({_al_u4845_o,_al_u5805_o}),
    .c({_al_u3222_o,_al_u3222_o}),
    .d({\exu/lsu/n4 [14],_al_u4366_o}),
    .f({_al_u4846_o,_al_u5806_o}));
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4847|biu/bus_unit/mmu/reg3_b14  (
    .a({open_n28243,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [14],\biu/bus_unit/mmu_hwdata [14]}),
    .clk(clk_pad),
    .d({_al_u4846_o,hrdata_pad[14]}),
    .sr(rst_pad),
    .f({hwdata_pad[14],open_n28261}),
    .q({open_n28265,\biu/bus_unit/mmu_hwdata [14]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4850|biu/cache_ctrl_logic/reg2_b13  (
    .a({open_n28266,_al_u2705_o}),
    .b({_al_u4849_o,_al_u4848_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [13],\biu/cache_ctrl_logic/pte_temp [13]}),
    .mi({open_n28270,\biu/cache_ctrl_logic/pte_temp [13]}),
    .sr(rst_pad),
    .f({_al_u4850_o,_al_u4849_o}),
    .q({open_n28285,\biu/cache_ctrl_logic/l1i_pte [13]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4851|biu/bus_unit/mmu/reg3_b13  (
    .a({open_n28286,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [13],\biu/bus_unit/mmu_hwdata [13]}),
    .clk(clk_pad),
    .d({_al_u4850_o,hrdata_pad[13]}),
    .sr(rst_pad),
    .f({hwdata_pad[13],open_n28300}),
    .q({open_n28304,\biu/bus_unit/mmu_hwdata [13]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4854|biu/cache_ctrl_logic/reg2_b12  (
    .a({open_n28305,_al_u2705_o}),
    .b({_al_u4853_o,_al_u4852_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [12],\biu/cache_ctrl_logic/pte_temp [12]}),
    .mi({open_n28309,\biu/cache_ctrl_logic/pte_temp [12]}),
    .sr(rst_pad),
    .f({_al_u4854_o,_al_u4853_o}),
    .q({open_n28324,\biu/cache_ctrl_logic/l1i_pte [12]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4855|biu/bus_unit/mmu/reg3_b12  (
    .a({open_n28325,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [12],\biu/bus_unit/mmu_hwdata [12]}),
    .clk(clk_pad),
    .d({_al_u4854_o,hrdata_pad[12]}),
    .sr(rst_pad),
    .f({hwdata_pad[12],open_n28339}),
    .q({open_n28343,\biu/bus_unit/mmu_hwdata [12]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4857|biu/cache_ctrl_logic/reg2_b11  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u4856_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [11]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [11],\biu/cache_ctrl_logic/pte_temp [11]}),
    .mi({open_n28347,\biu/cache_ctrl_logic/pte_temp [11]}),
    .sr(rst_pad),
    .f({_al_u4857_o,_al_u4856_o}),
    .q({open_n28362,\biu/cache_ctrl_logic/l1i_pte [11]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*~D))"),
    //.LUTF1("(B*~(~C*D))"),
    //.LUTG0("(B*~(~C*~D))"),
    //.LUTG1("(B*~(~C*D))"),
    .INIT_LUTF0(16'b1100110011000000),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b1100110011000000),
    .INIT_LUTG1(16'b1100000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4858|_al_u5710  (
    .b({_al_u4857_o,_al_u5709_o}),
    .c({_al_u3222_o,_al_u3222_o}),
    .d({\exu/lsu/n4 [11],_al_u4270_o}),
    .f({_al_u4858_o,_al_u5710_o}));
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4859|biu/bus_unit/mmu/reg3_b11  (
    .a({open_n28389,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [11],\biu/bus_unit/mmu_hwdata [11]}),
    .clk(clk_pad),
    .d({_al_u4858_o,hrdata_pad[11]}),
    .sr(rst_pad),
    .f({hwdata_pad[11],open_n28407}),
    .q({open_n28411,\biu/bus_unit/mmu_hwdata [11]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4862|biu/cache_ctrl_logic/reg2_b10  (
    .a({open_n28412,_al_u2705_o}),
    .b({_al_u4861_o,_al_u4860_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\exu/lsu/n4 [10],\biu/cache_ctrl_logic/pte_temp [10]}),
    .mi({open_n28423,\biu/cache_ctrl_logic/pte_temp [10]}),
    .sr(rst_pad),
    .f({_al_u4862_o,_al_u4861_o}),
    .q({open_n28427,\biu/cache_ctrl_logic/l1i_pte [10]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4863|biu/bus_unit/mmu/reg3_b10  (
    .a({open_n28428,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [10],\biu/bus_unit/mmu_hwdata [10]}),
    .clk(clk_pad),
    .d({_al_u4862_o,hrdata_pad[10]}),
    .sr(rst_pad),
    .f({hwdata_pad[10],open_n28446}),
    .q({open_n28450,\biu/bus_unit/mmu_hwdata [10]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4865|biu/cache_ctrl_logic/reg2_b9  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u4864_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [9]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [9],\biu/cache_ctrl_logic/pte_temp [9]}),
    .mi({open_n28454,\biu/cache_ctrl_logic/pte_temp [9]}),
    .sr(rst_pad),
    .f({_al_u4865_o,_al_u4864_o}),
    .q({open_n28469,\biu/cache_ctrl_logic/l1i_pte [9]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b0000000011001010),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u4866|_al_u4157  (
    .a({open_n28470,\exu/alu_data_mem_csr [9]}),
    .b({_al_u4865_o,\exu/alu_data_mem_csr [1]}),
    .c({_al_u3222_o,addr_ex[0]}),
    .d({\exu/lsu/n4 [9],addr_ex[1]}),
    .f({_al_u4866_o,\exu/lsu/n4 [9]}));
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~D)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(C*~D)"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100001111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111100001111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4867|biu/bus_unit/mmu/reg3_b9  (
    .b({_al_u2705_o,open_n28493}),
    .c({\biu/bus_unit/mmu_hwdata [9],_al_u2966_o}),
    .clk(clk_pad),
    .d({_al_u4866_o,_al_u2963_o}),
    .sr(rst_pad),
    .f({hwdata_pad[9],open_n28511}),
    .q({open_n28515,\biu/bus_unit/mmu_hwdata [9]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4869|biu/cache_ctrl_logic/reg2_b8  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u4868_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [8]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [8],\biu/cache_ctrl_logic/pte_temp [8]}),
    .mi({open_n28519,\biu/cache_ctrl_logic/pte_temp [8]}),
    .sr(rst_pad),
    .f({_al_u4869_o,_al_u4868_o}),
    .q({open_n28534,\biu/cache_ctrl_logic/l1i_pte [8]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("(B*~(~C*D))"),
    .INIT_LUT0(16'b0000000011001010),
    .INIT_LUT1(16'b1100000011001100),
    .MODE("LOGIC"))
    \_al_u4870|_al_u4159  (
    .a({open_n28535,\exu/alu_data_mem_csr [8]}),
    .b({_al_u4869_o,\exu/alu_data_mem_csr [0]}),
    .c({_al_u3222_o,addr_ex[0]}),
    .d({\exu/lsu/n4 [8],addr_ex[1]}),
    .f({_al_u4870_o,\exu/lsu/n4 [8]}));
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4871|biu/bus_unit/mmu/reg3_b8  (
    .a({open_n28556,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [8],\biu/bus_unit/mmu_hwdata [8]}),
    .clk(clk_pad),
    .d({_al_u4870_o,hrdata_pad[8]}),
    .sr(rst_pad),
    .f({hwdata_pad[8],open_n28570}),
    .q({open_n28574,\biu/bus_unit/mmu_hwdata [8]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~B)*~(~D*A))"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(~(C*~B)*~(~D*A))"),
    //.LUTG1("(~C*~B*~D)"),
    .INIT_LUTF0(16'b1100111101000101),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1100111101000101),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4872|_al_u9170  (
    .a({open_n28575,id_rs1_index[3]}),
    .b(id_rs1_index[1:0]),
    .c({id_rs1_index[0],wb_rd_index[0]}),
    .d({id_rs1_index[2],wb_rd_index[3]}),
    .f({_al_u4872_o,_al_u9170_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4874|ins_dec/reg7_b9  (
    .a({\cu_ru/n45_lutinv ,open_n28600}),
    .b({\cu_ru/al_ram_gpr_do_i0_009 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_009 ,id_ins_pc[9]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[9]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[9],open_n28613}),
    .q({open_n28617,as1[9]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4877|ins_dec/reg7_b8  (
    .a({\cu_ru/n45_lutinv ,open_n28618}),
    .b({\cu_ru/al_ram_gpr_do_i0_008 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_008 ,id_ins_pc[8]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[8]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[8],open_n28635}),
    .q({open_n28639,as1[8]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4879|ins_dec/reg7_b7  (
    .a({\cu_ru/n45_lutinv ,open_n28640}),
    .b({\cu_ru/al_ram_gpr_do_i0_007 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_007 ,id_ins_pc[7]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[7]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[7],open_n28657}),
    .q({open_n28661,as1[7]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4881|_al_u5001  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_063 ,\cu_ru/al_ram_gpr_do_i0_000 }),
    .c({\cu_ru/al_ram_gpr_do_i1_063 ,\cu_ru/al_ram_gpr_do_i1_000 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[63],rs1_data[0]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4883|_al_u4993  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_062 ,\cu_ru/al_ram_gpr_do_i0_012 }),
    .c({\cu_ru/al_ram_gpr_do_i1_062 ,\cu_ru/al_ram_gpr_do_i1_012 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[62],rs1_data[12]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"))
    \_al_u4885|_al_u4991  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_061 ,\cu_ru/al_ram_gpr_do_i0_013 }),
    .c({\cu_ru/al_ram_gpr_do_i1_061 ,\cu_ru/al_ram_gpr_do_i1_013 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[61],rs1_data[13]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"))
    \_al_u4887|_al_u4989  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_060 ,\cu_ru/al_ram_gpr_do_i0_014 }),
    .c({\cu_ru/al_ram_gpr_do_i1_060 ,\cu_ru/al_ram_gpr_do_i1_014 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[60],rs1_data[14]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4889|ins_dec/reg7_b6  (
    .a({\cu_ru/n45_lutinv ,open_n28750}),
    .b({\cu_ru/al_ram_gpr_do_i0_006 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_006 ,id_ins_pc[6]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[6]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[6],open_n28763}),
    .q({open_n28767,as1[6]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4891|_al_u4985  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_059 ,\cu_ru/al_ram_gpr_do_i0_016 }),
    .c({\cu_ru/al_ram_gpr_do_i1_059 ,\cu_ru/al_ram_gpr_do_i1_016 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[59],rs1_data[16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4893|_al_u4983  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_058 ,\cu_ru/al_ram_gpr_do_i0_017 }),
    .c({\cu_ru/al_ram_gpr_do_i1_058 ,\cu_ru/al_ram_gpr_do_i1_017 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[58],rs1_data[17]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"))
    \_al_u4895|_al_u4981  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_057 ,\cu_ru/al_ram_gpr_do_i0_018 }),
    .c({\cu_ru/al_ram_gpr_do_i1_057 ,\cu_ru/al_ram_gpr_do_i1_018 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[57],rs1_data[18]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"))
    \_al_u4897|_al_u4979  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_056 ,\cu_ru/al_ram_gpr_do_i0_019 }),
    .c({\cu_ru/al_ram_gpr_do_i1_056 ,\cu_ru/al_ram_gpr_do_i1_019 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[56],rs1_data[19]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4899|_al_u4975  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_055 ,\cu_ru/al_ram_gpr_do_i0_020 }),
    .c({\cu_ru/al_ram_gpr_do_i1_055 ,\cu_ru/al_ram_gpr_do_i1_020 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[55],rs1_data[20]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4901|_al_u4973  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_054 ,\cu_ru/al_ram_gpr_do_i0_021 }),
    .c({\cu_ru/al_ram_gpr_do_i1_054 ,\cu_ru/al_ram_gpr_do_i1_021 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[54],rs1_data[21]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"))
    \_al_u4903|_al_u4971  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_053 ,\cu_ru/al_ram_gpr_do_i0_022 }),
    .c({\cu_ru/al_ram_gpr_do_i1_053 ,\cu_ru/al_ram_gpr_do_i1_022 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[53],rs1_data[22]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"))
    \_al_u4905|_al_u4969  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_052 ,\cu_ru/al_ram_gpr_do_i0_023 }),
    .c({\cu_ru/al_ram_gpr_do_i1_052 ,\cu_ru/al_ram_gpr_do_i1_023 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[52],rs1_data[23]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4907|_al_u4967  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_051 ,\cu_ru/al_ram_gpr_do_i0_024 }),
    .c({\cu_ru/al_ram_gpr_do_i1_051 ,\cu_ru/al_ram_gpr_do_i1_024 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[51],rs1_data[24]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4909|_al_u4965  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_050 ,\cu_ru/al_ram_gpr_do_i0_025 }),
    .c({\cu_ru/al_ram_gpr_do_i1_050 ,\cu_ru/al_ram_gpr_do_i1_025 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[50],rs1_data[25]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4911|ins_dec/reg7_b5  (
    .a({\cu_ru/n45_lutinv ,open_n28992}),
    .b({\cu_ru/al_ram_gpr_do_i0_005 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_005 ,id_ins_pc[5]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[5]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[5],open_n29009}),
    .q({open_n29013,as1[5]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"))
    \_al_u4913|_al_u4963  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_049 ,\cu_ru/al_ram_gpr_do_i0_026 }),
    .c({\cu_ru/al_ram_gpr_do_i1_049 ,\cu_ru/al_ram_gpr_do_i1_026 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[49],rs1_data[26]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"))
    \_al_u4915|_al_u4961  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_048 ,\cu_ru/al_ram_gpr_do_i0_027 }),
    .c({\cu_ru/al_ram_gpr_do_i1_048 ,\cu_ru/al_ram_gpr_do_i1_027 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[48],rs1_data[27]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4917|_al_u4959  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_047 ,\cu_ru/al_ram_gpr_do_i0_028 }),
    .c({\cu_ru/al_ram_gpr_do_i1_047 ,\cu_ru/al_ram_gpr_do_i1_028 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[47],rs1_data[28]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4919|_al_u4957  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_046 ,\cu_ru/al_ram_gpr_do_i0_029 }),
    .c({\cu_ru/al_ram_gpr_do_i1_046 ,\cu_ru/al_ram_gpr_do_i1_029 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[46],rs1_data[29]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"))
    \_al_u4921|_al_u4953  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_045 ,\cu_ru/al_ram_gpr_do_i0_030 }),
    .c({\cu_ru/al_ram_gpr_do_i1_045 ,\cu_ru/al_ram_gpr_do_i1_030 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[45],rs1_data[30]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4923|_al_u4949  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_044 ,\cu_ru/al_ram_gpr_do_i0_032 }),
    .c({\cu_ru/al_ram_gpr_do_i1_044 ,\cu_ru/al_ram_gpr_do_i1_032 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[44],rs1_data[32]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4925|_al_u4947  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_043 ,\cu_ru/al_ram_gpr_do_i0_033 }),
    .c({\cu_ru/al_ram_gpr_do_i1_043 ,\cu_ru/al_ram_gpr_do_i1_033 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[43],rs1_data[33]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"))
    \_al_u4927|_al_u4943  (
    .a({\cu_ru/n45_lutinv ,\cu_ru/n45_lutinv }),
    .b({\cu_ru/al_ram_gpr_do_i0_042 ,\cu_ru/al_ram_gpr_do_i0_035 }),
    .c({\cu_ru/al_ram_gpr_do_i1_042 ,\cu_ru/al_ram_gpr_do_i1_035 }),
    .d({\cu_ru/n46 [4],\cu_ru/n46 [4]}),
    .f({rs1_data[42],rs1_data[35]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4933|ins_dec/reg7_b4  (
    .a({\cu_ru/n45_lutinv ,open_n29190}),
    .b({\cu_ru/al_ram_gpr_do_i0_004 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_004 ,id_ins_pc[4]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[4]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[4],open_n29207}),
    .q({open_n29211,as1[4]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4955|ins_dec/reg7_b3  (
    .a({\cu_ru/n45_lutinv ,open_n29212}),
    .b({\cu_ru/al_ram_gpr_do_i0_003 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_003 ,id_ins_pc[3]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[3]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[3],open_n29225}),
    .q({open_n29229,as1[3]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4977|ins_dec/reg7_b2  (
    .a({\cu_ru/n45_lutinv ,open_n29230}),
    .b({\cu_ru/al_ram_gpr_do_i0_002 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_002 ,id_ins_pc[2]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[2]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[2],open_n29243}),
    .q({open_n29247,as1[2]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u4987|_al_u3965  (
    .a({\cu_ru/n45_lutinv ,open_n29248}),
    .b({\cu_ru/al_ram_gpr_do_i0_015 ,1'b0}),
    .c({\cu_ru/al_ram_gpr_do_i1_015 ,\ins_fetch/ins_hold [15]}),
    .d({\cu_ru/n46 [4],\ins_fetch/ins_shift [15]}),
    .f({rs1_data[15],id_ins[15]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4995|ins_dec/reg7_b11  (
    .a({\cu_ru/n45_lutinv ,open_n29273}),
    .b({\cu_ru/al_ram_gpr_do_i0_011 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_011 ,id_ins_pc[11]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[11]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[11],open_n29290}),
    .q({open_n29294,as1[11]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4997|ins_dec/reg7_b10  (
    .a({\cu_ru/n45_lutinv ,open_n29295}),
    .b({\cu_ru/al_ram_gpr_do_i0_010 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_010 ,id_ins_pc[10]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[10]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[10],open_n29308}),
    .q({open_n29312,as1[10]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u4999|ins_dec/reg7_b1  (
    .a({\cu_ru/n45_lutinv ,open_n29313}),
    .b({\cu_ru/al_ram_gpr_do_i0_001 ,_al_u4875_o}),
    .c({\cu_ru/al_ram_gpr_do_i1_001 ,id_ins_pc[1]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n46 [4],rs1_data[1]}),
    .sr(\ins_dec/n107 ),
    .f({rs1_data[1],open_n29326}),
    .q({open_n29330,as1[1]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*~A))"),
    //.LUT1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100100011001100),
    .INIT_LUT1(16'b1100111101000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5003|biu/bus_unit/mmu/reg1_b63  (
    .a({_al_u2914_o,\biu/maddress [63]}),
    .b({_al_u2698_o,_al_u5003_o}),
    .c({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,_al_u2914_o}),
    .clk(clk_pad),
    .d({\biu/paddress [63],_al_u2698_o}),
    .sr(rst_pad),
    .f({_al_u5003_o,open_n29344}),
    .q({open_n29348,\biu/paddress [63]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*~A))"),
    //.LUT1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100100011001100),
    .INIT_LUT1(16'b1100111101000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5005|biu/bus_unit/mmu/reg1_b62  (
    .a({_al_u2914_o,\biu/maddress [62]}),
    .b({_al_u2698_o,_al_u5005_o}),
    .c({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,_al_u2914_o}),
    .clk(clk_pad),
    .d({\biu/paddress [62],_al_u2698_o}),
    .sr(rst_pad),
    .f({_al_u5005_o,open_n29362}),
    .q({open_n29366,\biu/paddress [62]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*~A))"),
    //.LUTF1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(B*~(D*~C*~A))"),
    //.LUTG1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100100011001100),
    .INIT_LUTF1(16'b1100111101000100),
    .INIT_LUTG0(16'b1100100011001100),
    .INIT_LUTG1(16'b1100111101000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5007|biu/bus_unit/mmu/reg1_b61  (
    .a({_al_u2914_o,\biu/maddress [61]}),
    .b({_al_u2698_o,_al_u5007_o}),
    .c({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,_al_u2914_o}),
    .clk(clk_pad),
    .d({\biu/paddress [61],_al_u2698_o}),
    .sr(rst_pad),
    .f({_al_u5007_o,open_n29384}),
    .q({open_n29388,\biu/paddress [61]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*~A))"),
    //.LUTF1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(B*~(D*~C*~A))"),
    //.LUTG1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100100011001100),
    .INIT_LUTF1(16'b1100111101000100),
    .INIT_LUTG0(16'b1100100011001100),
    .INIT_LUTG1(16'b1100111101000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5009|biu/bus_unit/mmu/reg1_b60  (
    .a({_al_u2914_o,\biu/maddress [60]}),
    .b({_al_u2698_o,_al_u5009_o}),
    .c({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,_al_u2914_o}),
    .clk(clk_pad),
    .d({\biu/paddress [60],_al_u2698_o}),
    .sr(rst_pad),
    .f({_al_u5009_o,open_n29406}),
    .q({open_n29410,\biu/paddress [60]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*~A))"),
    //.LUT1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100100011001100),
    .INIT_LUT1(16'b1100111101000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5011|biu/bus_unit/mmu/reg1_b59  (
    .a({_al_u2914_o,\biu/maddress [59]}),
    .b({_al_u2698_o,_al_u5011_o}),
    .c({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,_al_u2914_o}),
    .clk(clk_pad),
    .d({\biu/paddress [59],_al_u2698_o}),
    .sr(rst_pad),
    .f({_al_u5011_o,open_n29424}),
    .q({open_n29428,\biu/paddress [59]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~C*~A))"),
    //.LUT1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100100011001100),
    .INIT_LUT1(16'b1100111101000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5013|biu/bus_unit/mmu/reg1_b58  (
    .a({_al_u2914_o,\biu/maddress [58]}),
    .b({_al_u2698_o,_al_u5013_o}),
    .c({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,_al_u2914_o}),
    .clk(clk_pad),
    .d({\biu/paddress [58],_al_u2698_o}),
    .sr(rst_pad),
    .f({_al_u5013_o,open_n29442}),
    .q({open_n29446,\biu/paddress [58]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*~A))"),
    //.LUTF1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(B*~(D*~C*~A))"),
    //.LUTG1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100100011001100),
    .INIT_LUTF1(16'b1100111101000100),
    .INIT_LUTG0(16'b1100100011001100),
    .INIT_LUTG1(16'b1100111101000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5015|biu/bus_unit/mmu/reg1_b57  (
    .a({_al_u2914_o,\biu/maddress [57]}),
    .b({_al_u2698_o,_al_u5015_o}),
    .c({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,_al_u2914_o}),
    .clk(clk_pad),
    .d({\biu/paddress [57],_al_u2698_o}),
    .sr(rst_pad),
    .f({_al_u5015_o,open_n29464}),
    .q({open_n29468,\biu/paddress [57]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*~A))"),
    //.LUTF1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(B*~(D*~C*~A))"),
    //.LUTG1("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100100011001100),
    .INIT_LUTF1(16'b1100111101000100),
    .INIT_LUTG0(16'b1100100011001100),
    .INIT_LUTG1(16'b1100111101000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5017|biu/bus_unit/mmu/reg1_b56  (
    .a({_al_u2914_o,\biu/maddress [56]}),
    .b({_al_u2698_o,_al_u5017_o}),
    .c({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,_al_u2914_o}),
    .clk(clk_pad),
    .d({\biu/paddress [56],_al_u2698_o}),
    .sr(rst_pad),
    .f({_al_u5017_o,open_n29486}),
    .q({open_n29490,\biu/paddress [56]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5019|biu/cache_ctrl_logic/reg6_b55  (
    .a({\biu/maddress [55],open_n29491}),
    .b({_al_u2914_o,\biu/paddress [55]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [55]}),
    .clk(clk_pad),
    .d({\biu/paddress [55],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5019_o,open_n29509}),
    .q({open_n29513,\biu/cache_ctrl_logic/pa_temp [55]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5020|biu/bus_unit/mmu/reg3_b53  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [55],\biu/bus_unit/mmu_hwdata [53]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [53],hrdata_pad[53]}),
    .sr(rst_pad),
    .f({_al_u5020_o,open_n29527}),
    .q({open_n29531,\biu/bus_unit/mmu_hwdata [53]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5022|biu/cache_ctrl_logic/reg6_b54  (
    .a({\biu/maddress [54],open_n29532}),
    .b({_al_u2914_o,\biu/paddress [54]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [54]}),
    .clk(clk_pad),
    .d({\biu/paddress [54],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5022_o,open_n29546}),
    .q({open_n29550,\biu/cache_ctrl_logic/pa_temp [54]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5023|biu/bus_unit/mmu/reg3_b52  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [54],\biu/bus_unit/mmu_hwdata [52]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [52],hrdata_pad[52]}),
    .sr(rst_pad),
    .f({_al_u5023_o,open_n29564}),
    .q({open_n29568,\biu/bus_unit/mmu_hwdata [52]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5025|biu/cache_ctrl_logic/reg6_b53  (
    .a({\biu/maddress [53],open_n29569}),
    .b({_al_u2914_o,\biu/paddress [53]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [53]}),
    .clk(clk_pad),
    .d({\biu/paddress [53],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5025_o,open_n29583}),
    .q({open_n29587,\biu/cache_ctrl_logic/pa_temp [53]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5026|biu/bus_unit/mmu/reg3_b51  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [53],\biu/bus_unit/mmu_hwdata [51]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [51],hrdata_pad[51]}),
    .sr(rst_pad),
    .f({_al_u5026_o,open_n29605}),
    .q({open_n29609,\biu/bus_unit/mmu_hwdata [51]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5028|biu/cache_ctrl_logic/reg6_b52  (
    .a({\biu/maddress [52],open_n29610}),
    .b({_al_u2914_o,\biu/paddress [52]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [52]}),
    .clk(clk_pad),
    .d({\biu/paddress [52],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5028_o,open_n29624}),
    .q({open_n29628,\biu/cache_ctrl_logic/pa_temp [52]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5029|biu/bus_unit/mmu/reg3_b50  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [52],\biu/bus_unit/mmu_hwdata [50]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [50],hrdata_pad[50]}),
    .sr(rst_pad),
    .f({_al_u5029_o,open_n29646}),
    .q({open_n29650,\biu/bus_unit/mmu_hwdata [50]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5031|biu/cache_ctrl_logic/reg6_b51  (
    .a({\biu/maddress [51],open_n29651}),
    .b({_al_u2914_o,\biu/paddress [51]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [51]}),
    .clk(clk_pad),
    .d({\biu/paddress [51],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5031_o,open_n29669}),
    .q({open_n29673,\biu/cache_ctrl_logic/pa_temp [51]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5032|biu/bus_unit/mmu/reg3_b49  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [51],\biu/bus_unit/mmu_hwdata [49]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [49],hrdata_pad[49]}),
    .sr(rst_pad),
    .f({_al_u5032_o,open_n29687}),
    .q({open_n29691,\biu/bus_unit/mmu_hwdata [49]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5034|biu/cache_ctrl_logic/reg6_b50  (
    .a({\biu/maddress [50],open_n29692}),
    .b({_al_u2914_o,\biu/paddress [50]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [50]}),
    .clk(clk_pad),
    .d({\biu/paddress [50],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5034_o,open_n29710}),
    .q({open_n29714,\biu/cache_ctrl_logic/pa_temp [50]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5035|biu/bus_unit/mmu/reg3_b48  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [50],\biu/bus_unit/mmu_hwdata [48]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [48],hrdata_pad[48]}),
    .sr(rst_pad),
    .f({_al_u5035_o,open_n29728}),
    .q({open_n29732,\biu/bus_unit/mmu_hwdata [48]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5037|biu/cache_ctrl_logic/reg6_b49  (
    .a({\biu/maddress [49],open_n29733}),
    .b({_al_u2914_o,\biu/paddress [49]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [49]}),
    .clk(clk_pad),
    .d({\biu/paddress [49],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5037_o,open_n29751}),
    .q({open_n29755,\biu/cache_ctrl_logic/pa_temp [49]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5038|biu/bus_unit/mmu/reg3_b47  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [49],\biu/bus_unit/mmu_hwdata [47]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [47],hrdata_pad[47]}),
    .sr(rst_pad),
    .f({_al_u5038_o,open_n29773}),
    .q({open_n29777,\biu/bus_unit/mmu_hwdata [47]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5040|biu/cache_ctrl_logic/reg6_b48  (
    .a({\biu/maddress [48],open_n29778}),
    .b({_al_u2914_o,\biu/paddress [48]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [48]}),
    .clk(clk_pad),
    .d({\biu/paddress [48],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5040_o,open_n29796}),
    .q({open_n29800,\biu/cache_ctrl_logic/pa_temp [48]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5041|biu/bus_unit/mmu/reg3_b46  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [48],\biu/bus_unit/mmu_hwdata [46]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [46],hrdata_pad[46]}),
    .sr(rst_pad),
    .f({_al_u5041_o,open_n29818}),
    .q({open_n29822,\biu/bus_unit/mmu_hwdata [46]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5043|biu/cache_ctrl_logic/reg6_b47  (
    .a({\biu/maddress [47],open_n29823}),
    .b({_al_u2914_o,\biu/paddress [47]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [47]}),
    .clk(clk_pad),
    .d({\biu/paddress [47],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5043_o,open_n29837}),
    .q({open_n29841,\biu/cache_ctrl_logic/pa_temp [47]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5044|biu/bus_unit/mmu/reg3_b45  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [47],\biu/bus_unit/mmu_hwdata [45]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [45],hrdata_pad[45]}),
    .sr(rst_pad),
    .f({_al_u5044_o,open_n29855}),
    .q({open_n29859,\biu/bus_unit/mmu_hwdata [45]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5046|biu/cache_ctrl_logic/reg6_b46  (
    .a({\biu/maddress [46],open_n29860}),
    .b({_al_u2914_o,\biu/paddress [46]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [46]}),
    .clk(clk_pad),
    .d({\biu/paddress [46],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5046_o,open_n29874}),
    .q({open_n29878,\biu/cache_ctrl_logic/pa_temp [46]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5047|biu/bus_unit/mmu/reg3_b44  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [46],\biu/bus_unit/mmu_hwdata [44]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [44],hrdata_pad[44]}),
    .sr(rst_pad),
    .f({_al_u5047_o,open_n29892}),
    .q({open_n29896,\biu/bus_unit/mmu_hwdata [44]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5049|biu/cache_ctrl_logic/reg6_b45  (
    .a({\biu/maddress [45],open_n29897}),
    .b({_al_u2914_o,\biu/paddress [45]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [45]}),
    .clk(clk_pad),
    .d({\biu/paddress [45],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5049_o,open_n29915}),
    .q({open_n29919,\biu/cache_ctrl_logic/pa_temp [45]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5050|biu/bus_unit/mmu/reg3_b43  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [45],\biu/bus_unit/mmu_hwdata [43]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [43],hrdata_pad[43]}),
    .sr(rst_pad),
    .f({_al_u5050_o,open_n29937}),
    .q({open_n29941,\biu/bus_unit/mmu_hwdata [43]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5052|biu/cache_ctrl_logic/reg6_b44  (
    .a({\biu/maddress [44],open_n29942}),
    .b({_al_u2914_o,\biu/paddress [44]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [44]}),
    .clk(clk_pad),
    .d({\biu/paddress [44],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5052_o,open_n29956}),
    .q({open_n29960,\biu/cache_ctrl_logic/pa_temp [44]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5053|biu/bus_unit/mmu/reg3_b42  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [44],\biu/bus_unit/mmu_hwdata [42]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [42],hrdata_pad[42]}),
    .sr(rst_pad),
    .f({_al_u5053_o,open_n29978}),
    .q({open_n29982,\biu/bus_unit/mmu_hwdata [42]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5055|biu/cache_ctrl_logic/reg6_b43  (
    .a({\biu/maddress [43],open_n29983}),
    .b({_al_u2914_o,\biu/paddress [43]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [43]}),
    .clk(clk_pad),
    .d({\biu/paddress [43],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5055_o,open_n29997}),
    .q({open_n30001,\biu/cache_ctrl_logic/pa_temp [43]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5056|biu/bus_unit/mmu/reg3_b41  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [43],\biu/bus_unit/mmu_hwdata [41]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [41],hrdata_pad[41]}),
    .sr(rst_pad),
    .f({_al_u5056_o,open_n30015}),
    .q({open_n30019,\biu/bus_unit/mmu_hwdata [41]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5058|biu/cache_ctrl_logic/reg6_b42  (
    .a({\biu/maddress [42],open_n30020}),
    .b({_al_u2914_o,\biu/paddress [42]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [42]}),
    .clk(clk_pad),
    .d({\biu/paddress [42],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5058_o,open_n30038}),
    .q({open_n30042,\biu/cache_ctrl_logic/pa_temp [42]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5059|biu/bus_unit/mmu/reg3_b40  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [42],\biu/bus_unit/mmu_hwdata [40]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [40],hrdata_pad[40]}),
    .sr(rst_pad),
    .f({_al_u5059_o,open_n30056}),
    .q({open_n30060,\biu/bus_unit/mmu_hwdata [40]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5061|biu/cache_ctrl_logic/reg6_b41  (
    .a({\biu/maddress [41],open_n30061}),
    .b({_al_u2914_o,\biu/paddress [41]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [41]}),
    .clk(clk_pad),
    .d({\biu/paddress [41],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5061_o,open_n30075}),
    .q({open_n30079,\biu/cache_ctrl_logic/pa_temp [41]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5062|biu/bus_unit/mmu/reg3_b39  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [41],\biu/bus_unit/mmu_hwdata [39]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [39],hrdata_pad[39]}),
    .sr(rst_pad),
    .f({_al_u5062_o,open_n30097}),
    .q({open_n30101,\biu/bus_unit/mmu_hwdata [39]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5064|biu/cache_ctrl_logic/reg6_b40  (
    .a({\biu/maddress [40],open_n30102}),
    .b({_al_u2914_o,\biu/paddress [40]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [40]}),
    .clk(clk_pad),
    .d({\biu/paddress [40],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5064_o,open_n30116}),
    .q({open_n30120,\biu/cache_ctrl_logic/pa_temp [40]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5065|biu/bus_unit/mmu/reg3_b38  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [40],\biu/bus_unit/mmu_hwdata [38]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [38],hrdata_pad[38]}),
    .sr(rst_pad),
    .f({_al_u5065_o,open_n30138}),
    .q({open_n30142,\biu/bus_unit/mmu_hwdata [38]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5067|biu/cache_ctrl_logic/reg6_b39  (
    .a({\biu/maddress [39],open_n30143}),
    .b({_al_u2914_o,\biu/paddress [39]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [39]}),
    .clk(clk_pad),
    .d({\biu/paddress [39],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5067_o,open_n30161}),
    .q({open_n30165,\biu/cache_ctrl_logic/pa_temp [39]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5068|biu/bus_unit/mmu/reg3_b37  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [39],\biu/bus_unit/mmu_hwdata [37]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [37],hrdata_pad[37]}),
    .sr(rst_pad),
    .f({_al_u5068_o,open_n30179}),
    .q({open_n30183,\biu/bus_unit/mmu_hwdata [37]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5070|biu/cache_ctrl_logic/reg6_b38  (
    .a({\biu/maddress [38],open_n30184}),
    .b({_al_u2914_o,\biu/paddress [38]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [38]}),
    .clk(clk_pad),
    .d({\biu/paddress [38],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5070_o,open_n30202}),
    .q({open_n30206,\biu/cache_ctrl_logic/pa_temp [38]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5071|biu/bus_unit/mmu/reg3_b36  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [38],\biu/bus_unit/mmu_hwdata [36]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [36],hrdata_pad[36]}),
    .sr(rst_pad),
    .f({_al_u5071_o,open_n30220}),
    .q({open_n30224,\biu/bus_unit/mmu_hwdata [36]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5073|biu/cache_ctrl_logic/reg6_b37  (
    .a({\biu/maddress [37],open_n30225}),
    .b({_al_u2914_o,\biu/paddress [37]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [37]}),
    .clk(clk_pad),
    .d({\biu/paddress [37],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5073_o,open_n30239}),
    .q({open_n30243,\biu/cache_ctrl_logic/pa_temp [37]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5074|biu/bus_unit/mmu/reg3_b35  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [37],\biu/bus_unit/mmu_hwdata [35]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [35],hrdata_pad[35]}),
    .sr(rst_pad),
    .f({_al_u5074_o,open_n30261}),
    .q({open_n30265,\biu/bus_unit/mmu_hwdata [35]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5076|biu/cache_ctrl_logic/reg6_b36  (
    .a({\biu/maddress [36],open_n30266}),
    .b({_al_u2914_o,\biu/paddress [36]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [36]}),
    .clk(clk_pad),
    .d({\biu/paddress [36],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5076_o,open_n30280}),
    .q({open_n30284,\biu/cache_ctrl_logic/pa_temp [36]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5077|biu/bus_unit/mmu/reg3_b34  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [36],\biu/bus_unit/mmu_hwdata [34]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [34],hrdata_pad[34]}),
    .sr(rst_pad),
    .f({_al_u5077_o,open_n30302}),
    .q({open_n30306,\biu/bus_unit/mmu_hwdata [34]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5079|biu/cache_ctrl_logic/reg6_b35  (
    .a({\biu/maddress [35],open_n30307}),
    .b({_al_u2914_o,\biu/paddress [35]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [35]}),
    .clk(clk_pad),
    .d({\biu/paddress [35],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5079_o,open_n30325}),
    .q({open_n30329,\biu/cache_ctrl_logic/pa_temp [35]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5080|biu/bus_unit/mmu/reg3_b33  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [35],\biu/bus_unit/mmu_hwdata [33]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [33],hrdata_pad[33]}),
    .sr(rst_pad),
    .f({_al_u5080_o,open_n30343}),
    .q({open_n30347,\biu/bus_unit/mmu_hwdata [33]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5082|biu/cache_ctrl_logic/reg6_b34  (
    .a({\biu/maddress [34],open_n30348}),
    .b({_al_u2914_o,\biu/paddress [34]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [34]}),
    .clk(clk_pad),
    .d({\biu/paddress [34],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5082_o,open_n30366}),
    .q({open_n30370,\biu/cache_ctrl_logic/pa_temp [34]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5083|biu/bus_unit/mmu/reg3_b32  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [34],\biu/bus_unit/mmu_hwdata [32]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [32],hrdata_pad[32]}),
    .sr(rst_pad),
    .f({_al_u5083_o,open_n30384}),
    .q({open_n30388,\biu/bus_unit/mmu_hwdata [32]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5085|biu/cache_ctrl_logic/reg6_b33  (
    .a({\biu/maddress [33],open_n30389}),
    .b({_al_u2914_o,\biu/paddress [33]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [33]}),
    .clk(clk_pad),
    .d({\biu/paddress [33],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5085_o,open_n30403}),
    .q({open_n30407,\biu/cache_ctrl_logic/pa_temp [33]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5086|biu/bus_unit/mmu/reg3_b31  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [33],\biu/bus_unit/mmu_hwdata [31]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [31],hrdata_pad[31]}),
    .sr(rst_pad),
    .f({_al_u5086_o,open_n30425}),
    .q({open_n30429,\biu/bus_unit/mmu_hwdata [31]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5088|biu/cache_ctrl_logic/reg6_b32  (
    .a({\biu/maddress [32],open_n30430}),
    .b({_al_u2914_o,\biu/paddress [32]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [32]}),
    .clk(clk_pad),
    .d({\biu/paddress [32],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5088_o,open_n30444}),
    .q({open_n30448,\biu/cache_ctrl_logic/pa_temp [32]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5089|biu/bus_unit/mmu/reg3_b30  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [32],\biu/bus_unit/mmu_hwdata [30]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [30],hrdata_pad[30]}),
    .sr(rst_pad),
    .f({_al_u5089_o,open_n30466}),
    .q({open_n30470,\biu/bus_unit/mmu_hwdata [30]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5091|biu/cache_ctrl_logic/reg6_b31  (
    .a({\biu/maddress [31],open_n30471}),
    .b({_al_u2914_o,\biu/paddress [31]}),
    .c({_al_u2698_o,\biu/cache_ctrl_logic/pa_temp [31]}),
    .clk(clk_pad),
    .d({\biu/paddress [31],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5091_o,open_n30489}),
    .q({open_n30493,\biu/cache_ctrl_logic/pa_temp [31]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5092|biu/bus_unit/mmu/reg3_b29  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [31],\biu/bus_unit/mmu_hwdata [29]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [29],hrdata_pad[29]}),
    .sr(rst_pad),
    .f({_al_u5092_o,open_n30507}),
    .q({open_n30511,\biu/bus_unit/mmu_hwdata [29]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5094|biu/bus_unit/mmu/reg1_b30  (
    .a({\biu/maddress [30],open_n30512}),
    .b({_al_u2914_o,open_n30513}),
    .c({_al_u2698_o,_al_u5095_o}),
    .clk(clk_pad),
    .d({\biu/paddress [30],_al_u5094_o}),
    .sr(rst_pad),
    .f({_al_u5094_o,open_n30531}),
    .q({open_n30535,\biu/paddress [30]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5095|biu/bus_unit/mmu/reg3_b28  (
    .a({_al_u2698_o,_al_u2963_o}),
    .b({\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/paddress [30],\biu/bus_unit/mmu_hwdata [28]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [28],hrdata_pad[28]}),
    .sr(rst_pad),
    .f({_al_u5095_o,open_n30549}),
    .q({open_n30553,\biu/bus_unit/mmu_hwdata [28]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~B*~(D*C)))"),
    //.LUT1("(~A*~(D*~(C*~B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010001000100),
    .INIT_LUT1(16'b0001000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5099|exu/ins_page_fault_reg  (
    .a({\cu_ru/medeleg_exc_ctrl/iaf_target_m_lutinv ,\cu_ru/m_s_status/n5 [1]}),
    .b({priv[3],_al_u4119_o}),
    .c({\cu_ru/medeleg [12],\cu_ru/medeleg [12]}),
    .clk(clk_pad),
    .d({wb_ins_page_fault,wb_ins_page_fault}),
    .mi({open_n30565,ex_ins_page_fault}),
    .sr(\exu/n86 ),
    .f({_al_u5099_o,_al_u5154_o}),
    .q({open_n30569,wb_ins_page_fault}));  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*~(C*~B)))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001000001010101),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u5102|_al_u5100  (
    .a({open_n30570,\cu_ru/medeleg_exc_ctrl/lam_target_m_lutinv }),
    .b({_al_u5100_o,priv[3]}),
    .c({_al_u5101_o,\cu_ru/medeleg [3]}),
    .d({_al_u5099_o,wb_ebreak}),
    .f({_al_u5102_o,_al_u5100_o}));
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5103|cu_ru/medeleg_exc_ctrl/decu_reg  (
    .a({open_n30591,\cu_ru/read_mcause_sel_lutinv }),
    .b({\cu_ru/medeleg [8],\cu_ru/read_medeleg_sel_lutinv }),
    .c({wb_ecall,\cu_ru/mcause [8]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({priv[0],\cu_ru/medeleg [8]}),
    .mi({open_n30595,data_csr[8]}),
    .sr(rst_pad),
    .f({\cu_ru/medeleg_exc_ctrl/ecu_target_m ,_al_u7670_o}),
    .q({open_n30610,\cu_ru/medeleg [8]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~B*~(~D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000001100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5104|cu_ru/medeleg_exc_ctrl/decs_reg  (
    .a({_al_u4229_o,\cu_ru/read_mcause_sel_lutinv }),
    .b({\cu_ru/medeleg_exc_ctrl/iam_target_m_lutinv ,\cu_ru/read_medeleg_sel_lutinv }),
    .c({\cu_ru/medeleg_exc_ctrl/ecu_target_m ,\cu_ru/mcause [9]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/medeleg [9],\cu_ru/medeleg [9]}),
    .mi({open_n30621,data_csr[9]}),
    .sr(rst_pad),
    .f({_al_u5104_o,_al_u7810_o}),
    .q({open_n30625,\cu_ru/medeleg [9]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*~(C*~B)))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~A*~(D*~(C*~B)))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001000001010101),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001000001010101),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5107|_al_u5106  (
    .a({open_n30626,\cu_ru/medeleg_exc_ctrl/laf_target_m_lutinv }),
    .b({_al_u5105_o,priv[3]}),
    .c({_al_u5106_o,\cu_ru/medeleg [2]}),
    .d({_al_u5104_o,wb_ill_ins}),
    .f({_al_u5107_o,_al_u5106_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*C*~(B*~A))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1011000000000000),
    .MODE("LOGIC"))
    \_al_u5108|_al_u9188  (
    .a({\cu_ru/mideleg_int_ctrl/n28_lutinv ,open_n30651}),
    .b({_al_u5098_o,open_n30652}),
    .c({_al_u5102_o,wb_valid}),
    .d({_al_u5107_o,wb_gpr_write}),
    .f({_al_u5108_o,_al_u9188_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5112|biu/cache_ctrl_logic/reg2_b17  (
    .a({open_n30673,_al_u2705_o}),
    .b({_al_u5111_o,_al_u5110_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4205_o,\biu/cache_ctrl_logic/pte_temp [17]}),
    .mi({open_n30684,\biu/cache_ctrl_logic/pte_temp [17]}),
    .sr(rst_pad),
    .f({_al_u5112_o,_al_u5111_o}),
    .q({open_n30688,\biu/cache_ctrl_logic/l1i_pte [17]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5113|biu/bus_unit/mmu/reg3_b17  (
    .a({open_n30689,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [17],\biu/bus_unit/mmu_hwdata [17]}),
    .clk(clk_pad),
    .d({_al_u5112_o,hrdata_pad[17]}),
    .sr(rst_pad),
    .f({hwdata_pad[17],open_n30703}),
    .q({open_n30707,\biu/bus_unit/mmu_hwdata [17]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5115|biu/cache_ctrl_logic/reg2_b16  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u5114_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [16]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [16],\biu/cache_ctrl_logic/pte_temp [16]}),
    .mi({open_n30718,\biu/cache_ctrl_logic/pte_temp [16]}),
    .sr(rst_pad),
    .f({_al_u5115_o,_al_u5114_o}),
    .q({open_n30722,\biu/cache_ctrl_logic/l1i_pte [16]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5117|biu/bus_unit/mmu/reg3_b16  (
    .a({open_n30723,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [16],\biu/bus_unit/mmu_hwdata [16]}),
    .clk(clk_pad),
    .d({_al_u5116_o,hrdata_pad[16]}),
    .sr(rst_pad),
    .f({hwdata_pad[16],open_n30737}),
    .q({open_n30741,\biu/bus_unit/mmu_hwdata [16]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5120|biu/cache_ctrl_logic/reg5_b23  (
    .a({open_n30742,_al_u2705_o}),
    .b({_al_u5119_o,_al_u5118_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4211_o,\biu/cache_ctrl_logic/l1d_pte [23]}),
    .mi({open_n30753,\biu/cache_ctrl_logic/pte_temp [23]}),
    .sr(rst_pad),
    .f({_al_u5120_o,_al_u5119_o}),
    .q({open_n30757,\biu/cache_ctrl_logic/l1d_pte [23]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5121|biu/bus_unit/mmu/reg3_b23  (
    .a({open_n30758,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [23],\biu/bus_unit/mmu_hwdata [23]}),
    .clk(clk_pad),
    .d({_al_u5120_o,hrdata_pad[23]}),
    .sr(rst_pad),
    .f({hwdata_pad[23],open_n30776}),
    .q({open_n30780,\biu/bus_unit/mmu_hwdata [23]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5124|biu/cache_ctrl_logic/reg2_b22  (
    .a({open_n30781,_al_u2705_o}),
    .b({_al_u5123_o,_al_u5122_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4214_o,\biu/cache_ctrl_logic/pte_temp [22]}),
    .mi({open_n30792,\biu/cache_ctrl_logic/pte_temp [22]}),
    .sr(rst_pad),
    .f({_al_u5124_o,_al_u5123_o}),
    .q({open_n30796,\biu/cache_ctrl_logic/l1i_pte [22]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5125|biu/bus_unit/mmu/reg3_b22  (
    .a({open_n30797,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [22],\biu/bus_unit/mmu_hwdata [22]}),
    .clk(clk_pad),
    .d({_al_u5124_o,hrdata_pad[22]}),
    .sr(rst_pad),
    .f({hwdata_pad[22],open_n30815}),
    .q({open_n30819,\biu/bus_unit/mmu_hwdata [22]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5127|biu/cache_ctrl_logic/reg2_b21  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u5126_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [21]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [21],\biu/cache_ctrl_logic/pte_temp [21]}),
    .mi({open_n30823,\biu/cache_ctrl_logic/pte_temp [21]}),
    .sr(rst_pad),
    .f({_al_u5127_o,_al_u5126_o}),
    .q({open_n30838,\biu/cache_ctrl_logic/l1i_pte [21]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5129|biu/bus_unit/mmu/reg3_b21  (
    .a({open_n30839,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [21],\biu/bus_unit/mmu_hwdata [21]}),
    .clk(clk_pad),
    .d({_al_u5128_o,hrdata_pad[21]}),
    .sr(rst_pad),
    .f({hwdata_pad[21],open_n30853}),
    .q({open_n30857,\biu/bus_unit/mmu_hwdata [21]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5132|biu/cache_ctrl_logic/reg2_b20  (
    .a({open_n30858,_al_u2705_o}),
    .b({_al_u5131_o,_al_u5130_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4220_o,\biu/cache_ctrl_logic/pte_temp [20]}),
    .mi({open_n30862,\biu/cache_ctrl_logic/pte_temp [20]}),
    .sr(rst_pad),
    .f({_al_u5132_o,_al_u5131_o}),
    .q({open_n30877,\biu/cache_ctrl_logic/l1i_pte [20]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5133|biu/bus_unit/mmu/reg3_b20  (
    .a({open_n30878,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [20],\biu/bus_unit/mmu_hwdata [20]}),
    .clk(clk_pad),
    .d({_al_u5132_o,hrdata_pad[20]}),
    .sr(rst_pad),
    .f({hwdata_pad[20],open_n30892}),
    .q({open_n30896,\biu/bus_unit/mmu_hwdata [20]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5136|biu/cache_ctrl_logic/reg2_b19  (
    .a({open_n30897,_al_u2705_o}),
    .b({_al_u5135_o,_al_u5134_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4223_o,\biu/cache_ctrl_logic/pte_temp [19]}),
    .mi({open_n30901,\biu/cache_ctrl_logic/pte_temp [19]}),
    .sr(rst_pad),
    .f({_al_u5136_o,_al_u5135_o}),
    .q({open_n30916,\biu/cache_ctrl_logic/l1i_pte [19]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5137|biu/bus_unit/mmu/reg3_b19  (
    .a({open_n30917,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [19],\biu/bus_unit/mmu_hwdata [19]}),
    .clk(clk_pad),
    .d({_al_u5136_o,hrdata_pad[19]}),
    .sr(rst_pad),
    .f({hwdata_pad[19],open_n30935}),
    .q({open_n30939,\biu/bus_unit/mmu_hwdata [19]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5139|biu/cache_ctrl_logic/reg2_b18  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u5138_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [18]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [18],\biu/cache_ctrl_logic/pte_temp [18]}),
    .mi({open_n30950,\biu/cache_ctrl_logic/pte_temp [18]}),
    .sr(rst_pad),
    .f({_al_u5139_o,_al_u5138_o}),
    .q({open_n30954,\biu/cache_ctrl_logic/l1i_pte [18]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5141|biu/bus_unit/mmu/reg3_b18  (
    .a({open_n30955,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [18],\biu/bus_unit/mmu_hwdata [18]}),
    .clk(clk_pad),
    .d({_al_u5140_o,hrdata_pad[18]}),
    .sr(rst_pad),
    .f({hwdata_pad[18],open_n30973}),
    .q({open_n30977,\biu/bus_unit/mmu_hwdata [18]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*~B*~D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"))
    \_al_u5142|_al_u2675  (
    .b({id_ins[20],open_n30980}),
    .c({_al_u3392_o,\ins_fetch/ins_hold [24]}),
    .d({id_ins[22],1'b0}),
    .f({_al_u5142_o,_al_u2675_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u5143|_al_u5144  (
    .c({id_ins[21],_al_u5143_o}),
    .d({_al_u5142_o,_al_u4086_o}),
    .f({_al_u5143_o,_al_u5144_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B*~A))"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(D*~(C*B*~A))"),
    //.LUTG1("(C*~B*D)"),
    .INIT_LUTF0(16'b1011111100000000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b1011111100000000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5147|_al_u5157  (
    .a({open_n31025,_al_u5147_o}),
    .b({_al_u3250_o,_al_u5152_o}),
    .c({_al_u5098_o,_al_u5156_o}),
    .d({\cu_ru/mideleg_int_ctrl/n28_lutinv ,wb_valid}),
    .f({_al_u5147_o,_al_u5157_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~C*~A*~(D*B))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~C*~A*~(D*B))"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000100000101),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5149|_al_u5148  (
    .a({\cu_ru/medeleg_exc_ctrl/iam_target_s ,open_n31050}),
    .b({_al_u4229_o,\cu_ru/medeleg [8]}),
    .c({\cu_ru/medeleg_exc_ctrl/ecu_target_s ,wb_ecall}),
    .d({\cu_ru/medeleg [9],priv[0]}),
    .f({_al_u5149_o,\cu_ru/medeleg_exc_ctrl/ecu_target_s }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*~(C*~B)))"),
    //.LUT1("(~A*~(~B*~(D*C)))"),
    .INIT_LUT0(16'b0001000001010101),
    .INIT_LUT1(16'b0101010001000100),
    .MODE("LOGIC"))
    \_al_u5151|_al_u5105  (
    .a({\cu_ru/m_s_status/n5 [1],\cu_ru/medeleg_exc_ctrl/saf_target_m_lutinv }),
    .b({_al_u4108_o,priv[3]}),
    .c({\cu_ru/medeleg [13],\cu_ru/medeleg [13]}),
    .d({wb_ld_page_fault,wb_ld_page_fault}),
    .f({_al_u5151_o,_al_u5105_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~D)"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(C*B*~D)"),
    //.LUTG1("(~D*~C*~B*A)"),
    .INIT_LUTF0(16'b0000000011000000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000011000000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5152|_al_u5150  (
    .a({_al_u5149_o,open_n31095}),
    .b({\cu_ru/medeleg_exc_ctrl/laf_target_s ,\cu_ru/medeleg [2]}),
    .c({\cu_ru/medeleg_exc_ctrl/ii_target_s ,wb_ill_ins}),
    .d({_al_u5151_o,\cu_ru/m_s_status/n5 [1]}),
    .f({_al_u5152_o,\cu_ru/medeleg_exc_ctrl/ii_target_s }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*~(C*~B)))"),
    //.LUT1("(C*B*~D)"),
    .INIT_LUT0(16'b0001000001010101),
    .INIT_LUT1(16'b0000000011000000),
    .MODE("LOGIC"))
    \_al_u5153|_al_u5101  (
    .a({open_n31120,\cu_ru/medeleg_exc_ctrl/spf_target_m_lutinv }),
    .b({\cu_ru/medeleg [6],priv[3]}),
    .c({wb_st_addr_mis,\cu_ru/medeleg [6]}),
    .d({\cu_ru/m_s_status/n5 [1],wb_st_addr_mis}),
    .f({\cu_ru/medeleg_exc_ctrl/sam_target_s ,_al_u5101_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B*A))"),
    //.LUT1("(~A*~(~B*~(D*C)))"),
    .INIT_LUT0(16'b1101111100000000),
    .INIT_LUT1(16'b0101010001000100),
    .MODE("LOGIC"))
    \_al_u5155|_al_u4141  (
    .a({\cu_ru/m_s_status/n5 [1],\cu_ru/m_s_status/n5 [1]}),
    .b({_al_u4123_o,priv[3]}),
    .c({\cu_ru/medeleg [3],\cu_ru/medeleg [3]}),
    .d({wb_ebreak,wb_ebreak}),
    .f({_al_u5155_o,_al_u4141_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5156|_al_u7488  (
    .a({\cu_ru/medeleg_exc_ctrl/sam_target_s ,open_n31161}),
    .b({\cu_ru/medeleg_exc_ctrl/spf_target_s ,_al_u7487_o}),
    .c({_al_u5154_o,\biu/bus_unit/mmu_hwdata [2]}),
    .d({_al_u5155_o,_al_u7486_o}),
    .f({_al_u5156_o,_al_u7488_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5158|_al_u3206  (
    .b({open_n31188,csr_index[1]}),
    .c({_al_u3184_o,csr_index[2]}),
    .d({_al_u3420_o,_al_u3183_o}),
    .f({_al_u5158_o,_al_u3206_o}));
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5162|exu/reg5_b9  (
    .b({wb_ins_pc[9],addr_ex[9]}),
    .c({wb_exc_code[9],ex_exc_code[9]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [9],open_n31228}),
    .q({open_n31232,wb_exc_code[9]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5165|exu/reg5_b8  (
    .b({wb_ins_pc[8],addr_ex[8]}),
    .c({wb_exc_code[8],ex_exc_code[8]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [8],open_n31248}),
    .q({open_n31252,wb_exc_code[8]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5168|exu/reg5_b7  (
    .b({wb_ins_pc[7],addr_ex[7]}),
    .c({wb_exc_code[7],ex_exc_code[7]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [7],open_n31272}),
    .q({open_n31276,wb_exc_code[7]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5170|cu_ru/m_s_tval/reg0_b63  (
    .b({\cu_ru/stval [63],_al_u5170_o}),
    .c({data_csr[63],\cu_ru/m_s_tval/n3 [63]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5170_o,open_n31291}),
    .q({open_n31295,\cu_ru/stval [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5171|exu/reg5_b63  (
    .b({wb_ins_pc[63],open_n31298}),
    .c({wb_exc_code[63],addr_ex[63]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [63],open_n31316}),
    .q({open_n31320,wb_exc_code[63]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5174|exu/reg5_b62  (
    .b({wb_ins_pc[62],open_n31323}),
    .c({wb_exc_code[62],addr_ex[62]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [62],open_n31337}),
    .q({open_n31341,wb_exc_code[62]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5177|exu/reg5_b61  (
    .b({wb_ins_pc[61],open_n31344}),
    .c({wb_exc_code[61],addr_ex[61]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [61],open_n31358}),
    .q({open_n31362,wb_exc_code[61]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5180|exu/reg5_b60  (
    .b({wb_ins_pc[60],open_n31365}),
    .c({wb_exc_code[60],addr_ex[60]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [60],open_n31379}),
    .q({open_n31383,wb_exc_code[60]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5183|exu/reg5_b6  (
    .b({wb_ins_pc[6],addr_ex[6]}),
    .c({wb_exc_code[6],ex_exc_code[6]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [6],open_n31399}),
    .q({open_n31403,wb_exc_code[6]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5185|cu_ru/m_s_tval/reg0_b59  (
    .b({\cu_ru/stval [59],_al_u5185_o}),
    .c({data_csr[59],\cu_ru/m_s_tval/n3 [59]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5185_o,open_n31422}),
    .q({open_n31426,\cu_ru/stval [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5186|cu_ru/m_s_tval/reg1_b59  (
    .b({wb_ins_pc[59],\cu_ru/trap_target_m }),
    .c({wb_exc_code[59],\cu_ru/m_s_tval/n3 [59]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6459_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [59],open_n31446}),
    .q({open_n31450,\cu_ru/mtval [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5188|cu_ru/m_s_tval/reg0_b58  (
    .b({\cu_ru/stval [58],_al_u5188_o}),
    .c({data_csr[58],\cu_ru/m_s_tval/n3 [58]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5188_o,open_n31469}),
    .q({open_n31473,\cu_ru/stval [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5189|exu/reg5_b58  (
    .b({wb_ins_pc[58],open_n31476}),
    .c({wb_exc_code[58],addr_ex[58]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [58],open_n31494}),
    .q({open_n31498,wb_exc_code[58]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5191|cu_ru/m_s_tval/reg0_b57  (
    .b({\cu_ru/stval [57],_al_u5191_o}),
    .c({data_csr[57],\cu_ru/m_s_tval/n3 [57]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5191_o,open_n31513}),
    .q({open_n31517,\cu_ru/stval [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5192|cu_ru/m_s_tval/reg1_b57  (
    .b({wb_ins_pc[57],\cu_ru/trap_target_m }),
    .c({wb_exc_code[57],\cu_ru/m_s_tval/n3 [57]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6463_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [57],open_n31533}),
    .q({open_n31537,\cu_ru/mtval [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5194|cu_ru/m_s_tval/reg0_b56  (
    .b({\cu_ru/stval [56],_al_u5194_o}),
    .c({data_csr[56],\cu_ru/m_s_tval/n3 [56]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5194_o,open_n31552}),
    .q({open_n31556,\cu_ru/stval [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5195|exu/reg5_b56  (
    .b({wb_ins_pc[56],open_n31559}),
    .c({wb_exc_code[56],addr_ex[56]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [56],open_n31577}),
    .q({open_n31581,wb_exc_code[56]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5197|cu_ru/m_s_tval/reg0_b55  (
    .b({\cu_ru/stval [55],_al_u5197_o}),
    .c({data_csr[55],\cu_ru/m_s_tval/n3 [55]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5197_o,open_n31600}),
    .q({open_n31604,\cu_ru/stval [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5198|exu/reg5_b55  (
    .b({wb_ins_pc[55],open_n31607}),
    .c({wb_exc_code[55],addr_ex[55]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [55],open_n31625}),
    .q({open_n31629,wb_exc_code[55]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5200|cu_ru/m_s_tval/reg0_b54  (
    .b({\cu_ru/stval [54],_al_u5200_o}),
    .c({data_csr[54],\cu_ru/m_s_tval/n3 [54]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5200_o,open_n31648}),
    .q({open_n31652,\cu_ru/stval [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5201|exu/reg5_b54  (
    .b({wb_ins_pc[54],open_n31655}),
    .c({wb_exc_code[54],addr_ex[54]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [54],open_n31669}),
    .q({open_n31673,wb_exc_code[54]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5203|cu_ru/m_s_tval/reg0_b53  (
    .b({\cu_ru/stval [53],_al_u5203_o}),
    .c({data_csr[53],\cu_ru/m_s_tval/n3 [53]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5203_o,open_n31688}),
    .q({open_n31692,\cu_ru/stval [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5204|cu_ru/m_s_tval/reg1_b53  (
    .b({wb_ins_pc[53],\cu_ru/trap_target_m }),
    .c({wb_exc_code[53],\cu_ru/m_s_tval/n3 [53]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6471_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [53],open_n31708}),
    .q({open_n31712,\cu_ru/mtval [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5206|cu_ru/m_s_tval/reg0_b52  (
    .b({\cu_ru/stval [52],_al_u5206_o}),
    .c({data_csr[52],\cu_ru/m_s_tval/n3 [52]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5206_o,open_n31727}),
    .q({open_n31731,\cu_ru/stval [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5207|cu_ru/m_s_tval/reg1_b52  (
    .b({wb_ins_pc[52],\cu_ru/trap_target_m }),
    .c({wb_exc_code[52],\cu_ru/m_s_tval/n3 [52]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6473_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [52],open_n31751}),
    .q({open_n31755,\cu_ru/mtval [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5209|cu_ru/m_s_tval/reg0_b51  (
    .b({\cu_ru/stval [51],_al_u5209_o}),
    .c({data_csr[51],\cu_ru/m_s_tval/n3 [51]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5209_o,open_n31774}),
    .q({open_n31778,\cu_ru/stval [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5210|cu_ru/m_s_tval/reg1_b51  (
    .b({wb_ins_pc[51],\cu_ru/trap_target_m }),
    .c({wb_exc_code[51],\cu_ru/m_s_tval/n3 [51]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6475_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [51],open_n31798}),
    .q({open_n31802,\cu_ru/mtval [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5212|cu_ru/m_s_tval/reg0_b50  (
    .b({\cu_ru/stval [50],_al_u5212_o}),
    .c({data_csr[50],\cu_ru/m_s_tval/n3 [50]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5212_o,open_n31821}),
    .q({open_n31825,\cu_ru/stval [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5213|cu_ru/m_s_tval/reg1_b50  (
    .b({wb_ins_pc[50],\cu_ru/trap_target_m }),
    .c({wb_exc_code[50],\cu_ru/m_s_tval/n3 [50]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6477_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [50],open_n31841}),
    .q({open_n31845,\cu_ru/mtval [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5216|exu/reg5_b5  (
    .b({wb_ins_pc[5],addr_ex[5]}),
    .c({wb_exc_code[5],ex_exc_code[5]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [5],open_n31865}),
    .q({open_n31869,wb_exc_code[5]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5218|cu_ru/m_s_tval/reg0_b49  (
    .b({\cu_ru/stval [49],_al_u5218_o}),
    .c({data_csr[49],\cu_ru/m_s_tval/n3 [49]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5218_o,open_n31884}),
    .q({open_n31888,\cu_ru/stval [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5219|cu_ru/m_s_tval/reg1_b49  (
    .b({wb_ins_pc[49],\cu_ru/trap_target_m }),
    .c({wb_exc_code[49],\cu_ru/m_s_tval/n3 [49]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6481_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [49],open_n31908}),
    .q({open_n31912,\cu_ru/mtval [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5221|cu_ru/m_s_tval/reg0_b48  (
    .b({\cu_ru/stval [48],_al_u5221_o}),
    .c({data_csr[48],\cu_ru/m_s_tval/n3 [48]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5221_o,open_n31931}),
    .q({open_n31935,\cu_ru/stval [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5222|cu_ru/m_s_tval/reg1_b48  (
    .b({wb_ins_pc[48],\cu_ru/trap_target_m }),
    .c({wb_exc_code[48],\cu_ru/m_s_tval/n3 [48]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6483_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [48],open_n31955}),
    .q({open_n31959,\cu_ru/mtval [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5224|cu_ru/m_s_tval/reg0_b47  (
    .b({\cu_ru/stval [47],_al_u5224_o}),
    .c({data_csr[47],\cu_ru/m_s_tval/n3 [47]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5224_o,open_n31978}),
    .q({open_n31982,\cu_ru/stval [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5225|cu_ru/m_s_tval/reg1_b47  (
    .b({wb_ins_pc[47],\cu_ru/trap_target_m }),
    .c({wb_exc_code[47],\cu_ru/m_s_tval/n3 [47]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6485_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [47],open_n31998}),
    .q({open_n32002,\cu_ru/mtval [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5227|cu_ru/m_s_tval/reg0_b46  (
    .b({\cu_ru/stval [46],_al_u5227_o}),
    .c({data_csr[46],\cu_ru/m_s_tval/n3 [46]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5227_o,open_n32017}),
    .q({open_n32021,\cu_ru/stval [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5228|cu_ru/m_s_tval/reg1_b46  (
    .b({wb_ins_pc[46],\cu_ru/trap_target_m }),
    .c({wb_exc_code[46],\cu_ru/m_s_tval/n3 [46]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6487_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [46],open_n32037}),
    .q({open_n32041,\cu_ru/mtval [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5230|cu_ru/m_s_tval/reg0_b45  (
    .b({\cu_ru/stval [45],_al_u5230_o}),
    .c({data_csr[45],\cu_ru/m_s_tval/n3 [45]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5230_o,open_n32056}),
    .q({open_n32060,\cu_ru/stval [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5231|cu_ru/m_s_tval/reg1_b45  (
    .b({wb_ins_pc[45],\cu_ru/trap_target_m }),
    .c({wb_exc_code[45],\cu_ru/m_s_tval/n3 [45]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6489_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [45],open_n32080}),
    .q({open_n32084,\cu_ru/mtval [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5233|cu_ru/m_s_tval/reg0_b44  (
    .b({\cu_ru/stval [44],_al_u5233_o}),
    .c({data_csr[44],\cu_ru/m_s_tval/n3 [44]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5233_o,open_n32103}),
    .q({open_n32107,\cu_ru/stval [44]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5234|exu/reg5_b44  (
    .b({wb_ins_pc[44],open_n32110}),
    .c({wb_exc_code[44],addr_ex[44]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [44],open_n32128}),
    .q({open_n32132,wb_exc_code[44]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5237|cu_ru/m_s_tval/reg1_b43  (
    .b({wb_ins_pc[43],\cu_ru/trap_target_m }),
    .c({wb_exc_code[43],\cu_ru/m_s_tval/n3 [43]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6493_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [43],open_n32148}),
    .q({open_n32152,\cu_ru/mtval [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5240|cu_ru/m_s_tval/reg1_b42  (
    .b({wb_ins_pc[42],\cu_ru/trap_target_m }),
    .c({wb_exc_code[42],\cu_ru/m_s_tval/n3 [42]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6495_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [42],open_n32168}),
    .q({open_n32172,\cu_ru/mtval [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5243|cu_ru/m_s_tval/reg0_b41  (
    .b({wb_ins_pc[41],_al_u5242_o}),
    .c({wb_exc_code[41],\cu_ru/m_s_tval/n3 [41]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u5157_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [41],open_n32187}),
    .q({open_n32191,\cu_ru/stval [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5246|exu/reg5_b40  (
    .b({wb_ins_pc[40],open_n32194}),
    .c({wb_exc_code[40],addr_ex[40]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [40],open_n32208}),
    .q({open_n32212,wb_exc_code[40]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5249|exu/reg5_b4  (
    .b({wb_ins_pc[4],addr_ex[4]}),
    .c({wb_exc_code[4],ex_exc_code[4]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [4],open_n32228}),
    .q({open_n32232,wb_exc_code[4]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5252|cu_ru/m_s_tval/reg0_b39  (
    .b({wb_ins_pc[39],_al_u5251_o}),
    .c({wb_exc_code[39],\cu_ru/m_s_tval/n3 [39]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u5157_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [39],open_n32247}),
    .q({open_n32251,\cu_ru/stval [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5255|exu/reg5_b38  (
    .b({wb_ins_pc[38],open_n32254}),
    .c({wb_exc_code[38],addr_ex[38]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [38],open_n32272}),
    .q({open_n32276,wb_exc_code[38]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5258|exu/reg5_b37  (
    .b({wb_ins_pc[37],open_n32279}),
    .c({wb_exc_code[37],addr_ex[37]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [37],open_n32293}),
    .q({open_n32297,wb_exc_code[37]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5261|exu/reg5_b36  (
    .b({wb_ins_pc[36],open_n32300}),
    .c({wb_exc_code[36],addr_ex[36]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [36],open_n32318}),
    .q({open_n32322,wb_exc_code[36]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5264|cu_ru/m_s_tval/reg1_b35  (
    .b({wb_ins_pc[35],\cu_ru/trap_target_m }),
    .c({wb_exc_code[35],\cu_ru/m_s_tval/n3 [35]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6511_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [35],open_n32338}),
    .q({open_n32342,\cu_ru/mtval [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5267|exu/reg5_b34  (
    .b({wb_ins_pc[34],open_n32345}),
    .c({wb_exc_code[34],addr_ex[34]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [34],open_n32359}),
    .q({open_n32363,wb_exc_code[34]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5270|cu_ru/m_s_tval/reg1_b33  (
    .b({wb_ins_pc[33],\cu_ru/trap_target_m }),
    .c({wb_exc_code[33],\cu_ru/m_s_tval/n3 [33]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6515_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [33],open_n32383}),
    .q({open_n32387,\cu_ru/mtval [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5273|cu_ru/m_s_tval/reg1_b32  (
    .b({wb_ins_pc[32],\cu_ru/trap_target_m }),
    .c({wb_exc_code[32],\cu_ru/m_s_tval/n3 [32]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6517_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [32],open_n32403}),
    .q({open_n32407,\cu_ru/mtval [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5276|cu_ru/m_s_tval/reg0_b31  (
    .b({wb_ins_pc[31],_al_u5275_o}),
    .c({wb_exc_code[31],\cu_ru/m_s_tval/n3 [31]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u5157_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [31],open_n32422}),
    .q({open_n32426,\cu_ru/stval [31]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5279|cu_ru/m_s_tval/reg1_b30  (
    .b({wb_ins_pc[30],\cu_ru/trap_target_m }),
    .c({wb_exc_code[30],\cu_ru/m_s_tval/n3 [30]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6521_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [30],open_n32446}),
    .q({open_n32450,\cu_ru/mtval [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5281|cu_ru/m_s_tval/reg0_b3  (
    .b({\cu_ru/stval [3],_al_u5281_o}),
    .c({data_csr[3],\cu_ru/m_s_tval/n3 [3]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5281_o,open_n32469}),
    .q({open_n32473,\cu_ru/stval [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5282|exu/reg5_b3  (
    .b({wb_ins_pc[3],addr_ex[3]}),
    .c({wb_exc_code[3],ex_exc_code[3]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [3],open_n32493}),
    .q({open_n32497,wb_exc_code[3]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5285|exu/reg5_b29  (
    .b({wb_ins_pc[29],addr_ex[29]}),
    .c({wb_exc_code[29],ex_exc_code[29]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [29],open_n32513}),
    .q({open_n32517,wb_exc_code[29]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5288|cu_ru/m_s_tval/reg1_b28  (
    .b({wb_ins_pc[28],\cu_ru/trap_target_m }),
    .c({wb_exc_code[28],\cu_ru/m_s_tval/n3 [28]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6527_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [28],open_n32533}),
    .q({open_n32537,\cu_ru/mtval [28]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5291|cu_ru/m_s_tval/reg1_b27  (
    .b({wb_ins_pc[27],\cu_ru/trap_target_m }),
    .c({wb_exc_code[27],\cu_ru/m_s_tval/n3 [27]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6529_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [27],open_n32557}),
    .q({open_n32561,\cu_ru/mtval [27]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5294|exu/reg5_b26  (
    .b({wb_ins_pc[26],addr_ex[26]}),
    .c({wb_exc_code[26],ex_exc_code[26]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [26],open_n32577}),
    .q({open_n32581,wb_exc_code[26]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5297|exu/reg5_b25  (
    .b({wb_ins_pc[25],addr_ex[25]}),
    .c({wb_exc_code[25],ex_exc_code[25]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [25],open_n32597}),
    .q({open_n32601,wb_exc_code[25]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5300|exu/reg5_b24  (
    .b({wb_ins_pc[24],addr_ex[24]}),
    .c({wb_exc_code[24],ex_exc_code[24]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [24],open_n32621}),
    .q({open_n32625,wb_exc_code[24]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5303|exu/reg5_b23  (
    .b({wb_ins_pc[23],addr_ex[23]}),
    .c({wb_exc_code[23],ex_exc_code[23]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [23],open_n32641}),
    .q({open_n32645,wb_exc_code[23]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5306|cu_ru/m_s_tval/reg1_b22  (
    .b({wb_ins_pc[22],\cu_ru/trap_target_m }),
    .c({wb_exc_code[22],\cu_ru/m_s_tval/n3 [22]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6539_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [22],open_n32665}),
    .q({open_n32669,\cu_ru/mtval [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5309|cu_ru/m_s_tval/reg1_b21  (
    .b({wb_ins_pc[21],\cu_ru/trap_target_m }),
    .c({wb_exc_code[21],\cu_ru/m_s_tval/n3 [21]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6541_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [21],open_n32685}),
    .q({open_n32689,\cu_ru/mtval [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5312|cu_ru/m_s_tval/reg1_b20  (
    .b({wb_ins_pc[20],\cu_ru/trap_target_m }),
    .c({wb_exc_code[20],\cu_ru/m_s_tval/n3 [20]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6543_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [20],open_n32705}),
    .q({open_n32709,\cu_ru/mtval [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5314|cu_ru/m_s_tval/reg0_b2  (
    .b({\cu_ru/stval [2],_al_u5314_o}),
    .c({data_csr[2],\cu_ru/m_s_tval/n3 [2]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5314_o,open_n32724}),
    .q({open_n32728,\cu_ru/stval [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5315|exu/reg5_b2  (
    .b({wb_ins_pc[2],addr_ex[2]}),
    .c({wb_exc_code[2],ex_exc_code[2]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [2],open_n32748}),
    .q({open_n32752,wb_exc_code[2]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5318|cu_ru/m_s_tval/reg1_b19  (
    .b({wb_ins_pc[19],\cu_ru/trap_target_m }),
    .c({wb_exc_code[19],\cu_ru/m_s_tval/n3 [19]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6547_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [19],open_n32772}),
    .q({open_n32776,\cu_ru/mtval [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5321|exu/reg5_b18  (
    .b({wb_ins_pc[18],addr_ex[18]}),
    .c({wb_exc_code[18],ex_exc_code[18]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [18],open_n32792}),
    .q({open_n32796,wb_exc_code[18]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5324|cu_ru/m_s_tval/reg1_b17  (
    .b({wb_ins_pc[17],\cu_ru/trap_target_m }),
    .c({wb_exc_code[17],\cu_ru/m_s_tval/n3 [17]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6551_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [17],open_n32812}),
    .q({open_n32816,\cu_ru/mtval [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5327|cu_ru/m_s_tval/reg0_b16  (
    .b({wb_ins_pc[16],_al_u5326_o}),
    .c({wb_exc_code[16],\cu_ru/m_s_tval/n3 [16]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u5157_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [16],open_n32831}),
    .q({open_n32835,\cu_ru/stval [16]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5330|exu/reg5_b15  (
    .b({wb_ins_pc[15],addr_ex[15]}),
    .c({wb_exc_code[15],ex_exc_code[15]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [15],open_n32855}),
    .q({open_n32859,wb_exc_code[15]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5333|exu/reg5_b14  (
    .b({wb_ins_pc[14],addr_ex[14]}),
    .c({wb_exc_code[14],ex_exc_code[14]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [14],open_n32879}),
    .q({open_n32883,wb_exc_code[14]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5336|exu/reg5_b13  (
    .b({wb_ins_pc[13],addr_ex[13]}),
    .c({wb_exc_code[13],ex_exc_code[13]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [13],open_n32903}),
    .q({open_n32907,wb_exc_code[13]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5339|cu_ru/m_s_tval/reg1_b12  (
    .b({wb_ins_pc[12],\cu_ru/trap_target_m }),
    .c({wb_exc_code[12],\cu_ru/m_s_tval/n3 [12]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6561_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [12],open_n32927}),
    .q({open_n32931,\cu_ru/mtval [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5341|cu_ru/m_s_cause/reg0_b11  (
    .a({open_n32932,_al_u5157_o}),
    .b({\cu_ru/stval [11],\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({data_csr[11],\cu_ru/scause [11]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,data_csr[11]}),
    .sr(rst_pad),
    .f({_al_u5341_o,open_n32949}),
    .q({open_n32953,\cu_ru/scause [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5342|exu/reg5_b11  (
    .b({wb_ins_pc[11],addr_ex[11]}),
    .c({wb_exc_code[11],ex_exc_code[11]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [11],open_n32973}),
    .q({open_n32977,wb_exc_code[11]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5344|cu_ru/m_s_tval/reg0_b10  (
    .b({\cu_ru/stval [10],_al_u5344_o}),
    .c({data_csr[10],\cu_ru/m_s_tval/n3 [10]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5344_o,open_n32996}),
    .q({open_n33000,\cu_ru/stval [10]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5345|cu_ru/m_s_tval/reg1_b10  (
    .b({wb_ins_pc[10],\cu_ru/trap_target_m }),
    .c({wb_exc_code[10],\cu_ru/m_s_tval/n3 [10]}),
    .clk(clk_pad),
    .d({_al_u5161_o,_al_u6565_o}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [10],open_n33016}),
    .q({open_n33020,\cu_ru/mtval [10]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5348|exu/reg5_b1  (
    .b({wb_ins_pc[1],addr_ex[1]}),
    .c({wb_exc_code[1],ex_exc_code[1]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [1],open_n33036}),
    .q({open_n33040,wb_exc_code[1]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5350|cu_ru/m_s_tval/reg0_b0  (
    .b({\cu_ru/stval [0],_al_u5350_o}),
    .c({data_csr[0],\cu_ru/m_s_tval/n3 [0]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u5350_o,open_n33055}),
    .q({open_n33059,\cu_ru/stval [0]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5351|exu/reg5_b0  (
    .b({wb_ins_pc[0],addr_ex[0]}),
    .c({wb_exc_code[0],ex_exc_code[0]}),
    .clk(clk_pad),
    .d({_al_u5161_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_tval/n3 [0],open_n33079}),
    .q({open_n33083,wb_exc_code[0]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*D)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111111),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5354|exu/pc_jmp_reg  (
    .b({pc_jmp,open_n33086}),
    .c({new_pc[9],pc_jmp}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [7],_al_u6055_o}),
    .mi({open_n33098,jmp}),
    .sr(rst_pad),
    .f({_al_u5354_o,pip_flush}),
    .q({open_n33102,pc_jmp}));  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0000110000111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0000110000111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5359|_al_u5599  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[8],new_pc[10]}),
    .d({\cu_ru/m_s_epc/n0 [6],\cu_ru/m_s_epc/n0 [8]}),
    .f({_al_u5359_o,_al_u5599_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0000110000111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0000110000111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5363|_al_u5595  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[7],new_pc[11]}),
    .d({\cu_ru/m_s_epc/n0 [5],\cu_ru/m_s_epc/n0 [9]}),
    .f({_al_u5363_o,_al_u5595_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5367|exu/reg3_b63  (
    .a({open_n33155,\biu/cache_ctrl_logic/l1d_va [49]}),
    .b({pc_jmp,\biu/cache_ctrl_logic/l1d_va [63]}),
    .c({new_pc[63],addr_ex[49]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [61],addr_ex[63]}),
    .mi({open_n33160,addr_ex[63]}),
    .sr(rst_pad),
    .f({_al_u5367_o,_al_u6261_o}),
    .q({open_n33175,new_pc[63]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5369|cu_ru/m_s_epc/reg0_b63  (
    .b({\cu_ru/sepc [63],_al_u5157_o}),
    .c({data_csr[63],_al_u5369_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ,\cu_ru/m_s_epc/n2 [63]}),
    .sr(rst_pad),
    .f({_al_u5369_o,open_n33194}),
    .q({open_n33198,\cu_ru/sepc [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5371|exu/reg3_b62  (
    .a({open_n33199,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({pc_jmp,_al_u4399_o}),
    .c({new_pc[62],\biu/cache_ctrl_logic/n209 [62]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [60],addr_ex[62]}),
    .mi({open_n33204,addr_ex[62]}),
    .sr(rst_pad),
    .f({_al_u5371_o,_al_u4423_o}),
    .q({open_n33219,new_pc[62]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5375|exu/reg3_b61  (
    .a({open_n33220,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({pc_jmp,_al_u4399_o}),
    .c({new_pc[61],\biu/cache_ctrl_logic/n209 [61]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [59],addr_ex[61]}),
    .mi({open_n33225,addr_ex[61]}),
    .sr(rst_pad),
    .f({_al_u5375_o,_al_u4431_o}),
    .q({open_n33240,new_pc[61]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111000000010),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0000111000000010),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5379|exu/reg3_b60  (
    .a({open_n33241,_al_u9331_o}),
    .b({pc_jmp,_al_u6055_o}),
    .c({new_pc[60],_al_u2842_o}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [58],new_pc[60]}),
    .mi({open_n33246,addr_ex[60]}),
    .sr(rst_pad),
    .f({_al_u5379_o,_al_u9332_o}),
    .q({open_n33261,new_pc[60]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0000110000111111),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5383|_al_u5591  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[6],new_pc[12]}),
    .d({\cu_ru/m_s_epc/n0 [4],\cu_ru/m_s_epc/n0 [10]}),
    .f({_al_u5383_o,_al_u5591_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5387|exu/reg3_b59  (
    .a({open_n33284,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({pc_jmp,_al_u4399_o}),
    .c({new_pc[59],\biu/cache_ctrl_logic/n209 [59]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [57],addr_ex[59]}),
    .mi({open_n33296,addr_ex[59]}),
    .sr(rst_pad),
    .f({_al_u5387_o,_al_u4449_o}),
    .q({open_n33300,new_pc[59]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0000110000111111),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5391|_al_u5579  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[58],new_pc[15]}),
    .d({\cu_ru/m_s_epc/n0 [56],\cu_ru/m_s_epc/n0 [13]}),
    .f({_al_u5391_o,_al_u5579_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5395|exu/reg3_b57  (
    .a({open_n33323,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({pc_jmp,_al_u4399_o}),
    .c({new_pc[57],\biu/cache_ctrl_logic/n209 [57]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [55],addr_ex[57]}),
    .mi({open_n33328,addr_ex[57]}),
    .sr(rst_pad),
    .f({_al_u5395_o,_al_u4461_o}),
    .q({open_n33343,new_pc[57]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0000110000111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0000110000111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5399|_al_u5563  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[56],new_pc[19]}),
    .d({\cu_ru/m_s_epc/n0 [54],\cu_ru/m_s_epc/n0 [17]}),
    .f({_al_u5399_o,_al_u5563_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5403|exu/reg3_b55  (
    .a({open_n33370,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({pc_jmp,\biu/cache_ctrl_logic/n97_lutinv }),
    .c({new_pc[55],\biu/cache_ctrl_logic/n212 [55]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [53],addr_ex[55]}),
    .mi({open_n33375,addr_ex[55]}),
    .sr(rst_pad),
    .f({_al_u5403_o,_al_u4474_o}),
    .q({open_n33390,new_pc[55]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0000110000111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0000110000111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5407|_al_u5559  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[54],new_pc[2]}),
    .d({\cu_ru/m_s_epc/n0 [52],\cu_ru/m_s_epc/n0 [0]}),
    .f({_al_u5407_o,_al_u5559_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5411|exu/reg3_b53  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[53],new_pc[53]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [51],_al_u6055_o}),
    .mi({open_n33423,addr_ex[53]}),
    .sr(rst_pad),
    .f({_al_u5411_o,_al_u9373_o}),
    .q({open_n33438,new_pc[53]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0000110000111111),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5415|_al_u5543  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[52],new_pc[23]}),
    .d({\cu_ru/m_s_epc/n0 [50],\cu_ru/m_s_epc/n0 [21]}),
    .f({_al_u5415_o,_al_u5543_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0000110000111111),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5419|_al_u5487  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[51],new_pc[36]}),
    .d({\cu_ru/m_s_epc/n0 [49],\cu_ru/m_s_epc/n0 [34]}),
    .f({_al_u5419_o,_al_u5487_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0000110000111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0000110000111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5423|_al_u5471  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[50],new_pc[4]}),
    .d({\cu_ru/m_s_epc/n0 [48],\cu_ru/m_s_epc/n0 [2]}),
    .f({_al_u5423_o,_al_u5471_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0000110000111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0000110000111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5427|_al_u5467  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[5],new_pc[40]}),
    .d({\cu_ru/m_s_epc/n0 [3],\cu_ru/m_s_epc/n0 [38]}),
    .f({_al_u5427_o,_al_u5467_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0000110000111111),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5431|_al_u5455  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[49],new_pc[43]}),
    .d({\cu_ru/m_s_epc/n0 [47],\cu_ru/m_s_epc/n0 [41]}),
    .f({_al_u5431_o,_al_u5455_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0000110000111111),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5435|_al_u5443  (
    .b({pc_jmp,pc_jmp}),
    .c({new_pc[48],new_pc[46]}),
    .d({\cu_ru/m_s_epc/n0 [46],\cu_ru/m_s_epc/n0 [44]}),
    .f({_al_u5435_o,_al_u5443_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5439|exu/reg3_b47  (
    .a({open_n33579,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({pc_jmp,\biu/cache_ctrl_logic/n97_lutinv }),
    .c({new_pc[47],\biu/cache_ctrl_logic/n212 [47]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [45],addr_ex[47]}),
    .mi({open_n33591,addr_ex[47]}),
    .sr(rst_pad),
    .f({_al_u5439_o,_al_u4528_o}),
    .q({open_n33595,new_pc[47]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5447|_al_u9432  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[45],new_pc[45]}),
    .d({\cu_ru/m_s_epc/n0 [43],_al_u6055_o}),
    .f({_al_u5447_o,_al_u9432_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5451|exu/reg3_b44  (
    .a({open_n33622,\biu/cache_ctrl_logic/l1i_va [44]}),
    .b({pc_jmp,\biu/cache_ctrl_logic/l1i_va [46]}),
    .c({new_pc[44],addr_ex[44]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [42],addr_ex[46]}),
    .mi({open_n33634,addr_ex[44]}),
    .sr(rst_pad),
    .f({_al_u5451_o,_al_u6383_o}),
    .q({open_n33638,new_pc[44]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5459|_al_u9451  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[42],new_pc[42]}),
    .d({\cu_ru/m_s_epc/n0 [40],_al_u6055_o}),
    .f({_al_u5459_o,_al_u9451_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5463|_al_u9463  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[41],new_pc[41]}),
    .d({\cu_ru/m_s_epc/n0 [39],_al_u6055_o}),
    .f({_al_u5463_o,_al_u9463_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5475|_al_u9475  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[39],new_pc[39]}),
    .d({\cu_ru/m_s_epc/n0 [37],_al_u6055_o}),
    .f({_al_u5475_o,_al_u9475_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5479|_al_u9482  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[38],new_pc[38]}),
    .d({\cu_ru/m_s_epc/n0 [36],_al_u6055_o}),
    .f({_al_u5479_o,_al_u9482_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*A))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100110001),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5483|exu/reg3_b37  (
    .a({open_n33735,\biu/cache_ctrl_logic/l1d_va [30]}),
    .b({pc_jmp,\biu/cache_ctrl_logic/l1d_va [37]}),
    .c({new_pc[37],addr_ex[30]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [35],addr_ex[37]}),
    .mi({open_n33747,addr_ex[37]}),
    .sr(rst_pad),
    .f({_al_u5483_o,_al_u6302_o}),
    .q({open_n33751,new_pc[37]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5491|_al_u9501  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[35],new_pc[35]}),
    .d({\cu_ru/m_s_epc/n0 [33],_al_u6055_o}),
    .f({_al_u5491_o,_al_u9501_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5495|_al_u9508  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[34],new_pc[34]}),
    .d({\cu_ru/m_s_epc/n0 [32],_al_u6055_o}),
    .f({_al_u5495_o,_al_u9508_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5499|exu/reg3_b33  (
    .a({open_n33804,\biu/cache_ctrl_logic/l1d_va [33]}),
    .b({pc_jmp,\biu/cache_ctrl_logic/l1d_va [60]}),
    .c({new_pc[33],addr_ex[33]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [31],addr_ex[60]}),
    .mi({open_n33816,addr_ex[33]}),
    .sr(rst_pad),
    .f({_al_u5499_o,_al_u6259_o}),
    .q({open_n33820,new_pc[33]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5503|_al_u9520  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[32],new_pc[32]}),
    .d({\cu_ru/m_s_epc/n0 [30],_al_u6055_o}),
    .f({_al_u5503_o,_al_u9520_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5507|exu/reg3_b31  (
    .a({open_n33843,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({pc_jmp,\biu/cache_ctrl_logic/n97_lutinv }),
    .c({new_pc[31],\biu/cache_ctrl_logic/n212 [31]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [29],addr_ex[31]}),
    .mi({open_n33848,addr_ex[31]}),
    .sr(rst_pad),
    .f({_al_u5507_o,_al_u4630_o}),
    .q({open_n33863,new_pc[31]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5511|_al_u9539  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[30],new_pc[30]}),
    .d({\cu_ru/m_s_epc/n0 [28],_al_u6055_o}),
    .f({_al_u5511_o,_al_u9539_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5515|_al_u9600  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[3],new_pc[3]}),
    .d({\cu_ru/m_s_epc/n0 [1],_al_u6055_o}),
    .f({_al_u5515_o,_al_u9600_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5516|cu_ru/m_s_epc/reg0_b3  (
    .b({_al_u5515_o,_al_u5157_o}),
    .c({wb_ins_pc[3],_al_u5517_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u5353_o,\cu_ru/m_s_epc/n2 [3]}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [3],open_n33930}),
    .q({open_n33934,\cu_ru/sepc [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5519|exu/reg3_b29  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[29],new_pc[29]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [27],_al_u6055_o}),
    .mi({open_n33948,addr_ex[29]}),
    .sr(rst_pad),
    .f({_al_u5519_o,_al_u9546_o}),
    .q({open_n33952,new_pc[29]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5523|_al_u9553  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[28],new_pc[28]}),
    .d({\cu_ru/m_s_epc/n0 [26],_al_u6055_o}),
    .f({_al_u5523_o,_al_u9553_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5527|_al_u9560  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[27],new_pc[27]}),
    .d({\cu_ru/m_s_epc/n0 [25],_al_u6055_o}),
    .f({_al_u5527_o,_al_u9560_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5531|_al_u9567  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[26],new_pc[26]}),
    .d({\cu_ru/m_s_epc/n0 [24],_al_u6055_o}),
    .f({_al_u5531_o,_al_u9567_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5535|_al_u9574  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[25],new_pc[25]}),
    .d({\cu_ru/m_s_epc/n0 [23],_al_u6055_o}),
    .f({_al_u5535_o,_al_u9574_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5539|_al_u9581  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[24],new_pc[24]}),
    .d({\cu_ru/m_s_epc/n0 [22],_al_u6055_o}),
    .f({_al_u5539_o,_al_u9581_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5547|exu/reg3_b22  (
    .a({open_n34075,\biu/cache_ctrl_logic/n75_lutinv }),
    .b({pc_jmp,_al_u4399_o}),
    .c({new_pc[22],\biu/cache_ctrl_logic/n209 [22]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [20],addr_ex[22]}),
    .mi({open_n34087,addr_ex[22]}),
    .sr(rst_pad),
    .f({_al_u5547_o,_al_u4689_o}),
    .q({open_n34091,new_pc[22]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5551|exu/reg3_b21  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[21],new_pc[21]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [19],_al_u6055_o}),
    .mi({open_n34105,addr_ex[21]}),
    .sr(rst_pad),
    .f({_al_u5551_o,_al_u9607_o}),
    .q({open_n34109,new_pc[21]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5555|_al_u9614  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[20],new_pc[20]}),
    .d({\cu_ru/m_s_epc/n0 [18],_al_u6055_o}),
    .f({_al_u5555_o,_al_u9614_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5560|cu_ru/m_s_epc/reg0_b2  (
    .b({_al_u5559_o,_al_u5157_o}),
    .c({wb_ins_pc[2],_al_u5561_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u5353_o,\cu_ru/m_s_epc/n2 [2]}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [2],open_n34154}),
    .q({open_n34158,\cu_ru/sepc [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5567|_al_u9626  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[18],new_pc[18]}),
    .d({\cu_ru/m_s_epc/n0 [16],_al_u6055_o}),
    .f({_al_u5567_o,_al_u9626_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5571|_al_u9633  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[17],new_pc[17]}),
    .d({\cu_ru/m_s_epc/n0 [15],_al_u6055_o}),
    .f({_al_u5571_o,_al_u9633_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"))
    \_al_u5575|_al_u9640  (
    .b({pc_jmp,_al_u2844_o}),
    .c({new_pc[16],new_pc[16]}),
    .d({\cu_ru/m_s_epc/n0 [14],_al_u6055_o}),
    .f({_al_u5575_o,_al_u9640_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D@C))"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000001000),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5583|exu/reg3_b14  (
    .a({open_n34229,_al_u6244_o}),
    .b({pc_jmp,_al_u6245_o}),
    .c({new_pc[14],\biu/cache_ctrl_logic/l1d_va [14]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [12],addr_ex[14]}),
    .mi({open_n34241,addr_ex[14]}),
    .sr(rst_pad),
    .f({_al_u5583_o,_al_u6246_o}),
    .q({open_n34245,new_pc[14]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5587|exu/reg3_b13  (
    .b({pc_jmp,\biu/cache_ctrl_logic/l1d_va [13]}),
    .c({new_pc[13],addr_ex[13]}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/n0 [11],_al_u6293_o}),
    .mi({open_n34252,addr_ex[13]}),
    .sr(rst_pad),
    .f({_al_u5587_o,_al_u6294_o}),
    .q({open_n34267,new_pc[13]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5607|cu_ru/m_s_epc/reg0_b0  (
    .b({\cu_ru/sepc [0],_al_u5157_o}),
    .c({data_csr[0],_al_u5607_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ,\cu_ru/m_s_epc/n2 [0]}),
    .sr(rst_pad),
    .f({_al_u5607_o,open_n34286}),
    .q({open_n34290,\cu_ru/sepc [0]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5609|cu_ru/medeleg_exc_ctrl/dbk_reg  (
    .b({open_n34293,_al_u3206_o}),
    .c({_al_u3206_o,_al_u3184_o}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({_al_u5158_o,_al_u3195_o}),
    .mi({open_n34304,data_csr[3]}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ,\cu_ru/medeleg_exc_ctrl/n0 }),
    .q({open_n34308,\cu_ru/medeleg [3]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5613|cu_ru/m_s_cause/reg0_b63  (
    .c({_al_u4234_o,_al_u5614_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u5157_o,\cu_ru/n41 }),
    .sr(rst_pad),
    .f({\cu_ru/n41 ,open_n34325}),
    .q({open_n34329,\cu_ru/scause [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5614|cu_ru/m_s_cause/reg0_b7  (
    .a({_al_u5157_o,_al_u5157_o}),
    .b({\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [63],\cu_ru/scause [7]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({data_csr[63],data_csr[7]}),
    .sr(rst_pad),
    .f({_al_u5614_o,open_n34346}),
    .q({open_n34350,\cu_ru/scause [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5674|cu_ru/m_s_cause/reg0_b26  (
    .a({_al_u5157_o,_al_u5157_o}),
    .b({\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [0],\cu_ru/scause [26]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({data_csr[0],data_csr[26]}),
    .sr(rst_pad),
    .f({_al_u5674_o,open_n34367}),
    .q({open_n34371,\cu_ru/scause [26]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5678|biu/cache_ctrl_logic/reg2_b63  (
    .a({open_n34372,_al_u2705_o}),
    .b({_al_u5677_o,_al_u5676_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4238_o,\biu/cache_ctrl_logic/pte_temp [63]}),
    .mi({open_n34383,\biu/cache_ctrl_logic/pte_temp [63]}),
    .sr(rst_pad),
    .f({_al_u5678_o,_al_u5677_o}),
    .q({open_n34387,\biu/cache_ctrl_logic/l1i_pte [63]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5679|biu/bus_unit/mmu/reg3_b63  (
    .a({open_n34388,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [63],\biu/bus_unit/mmu_hwdata [63]}),
    .clk(clk_pad),
    .d({_al_u5678_o,hrdata_pad[63]}),
    .sr(rst_pad),
    .f({hwdata_pad[63],open_n34406}),
    .q({open_n34410,\biu/bus_unit/mmu_hwdata [63]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5682|biu/cache_ctrl_logic/reg2_b62  (
    .a({open_n34411,_al_u2705_o}),
    .b({_al_u5681_o,_al_u5680_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4242_o,\biu/cache_ctrl_logic/pte_temp [62]}),
    .mi({open_n34415,\biu/cache_ctrl_logic/pte_temp [62]}),
    .sr(rst_pad),
    .f({_al_u5682_o,_al_u5681_o}),
    .q({open_n34430,\biu/cache_ctrl_logic/l1i_pte [62]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5683|biu/bus_unit/mmu/reg3_b62  (
    .a({open_n34431,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [62],\biu/bus_unit/mmu_hwdata [62]}),
    .clk(clk_pad),
    .d({_al_u5682_o,hrdata_pad[62]}),
    .sr(rst_pad),
    .f({hwdata_pad[62],open_n34445}),
    .q({open_n34449,\biu/bus_unit/mmu_hwdata [62]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5686|biu/cache_ctrl_logic/reg5_b61  (
    .a({open_n34450,_al_u2705_o}),
    .b({_al_u5685_o,_al_u5684_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4246_o,\biu/cache_ctrl_logic/l1d_pte [61]}),
    .mi({open_n34454,\biu/cache_ctrl_logic/pte_temp [61]}),
    .sr(rst_pad),
    .f({_al_u5686_o,_al_u5685_o}),
    .q({open_n34469,\biu/cache_ctrl_logic/l1d_pte [61]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5687|biu/bus_unit/mmu/reg3_b61  (
    .a({open_n34470,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [61],\biu/bus_unit/mmu_hwdata [61]}),
    .clk(clk_pad),
    .d({_al_u5686_o,hrdata_pad[61]}),
    .sr(rst_pad),
    .f({hwdata_pad[61],open_n34484}),
    .q({open_n34488,\biu/bus_unit/mmu_hwdata [61]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5690|biu/cache_ctrl_logic/reg2_b60  (
    .a({open_n34489,_al_u2705_o}),
    .b({_al_u5689_o,_al_u5688_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4250_o,\biu/cache_ctrl_logic/pte_temp [60]}),
    .mi({open_n34493,\biu/cache_ctrl_logic/pte_temp [60]}),
    .sr(rst_pad),
    .f({_al_u5690_o,_al_u5689_o}),
    .q({open_n34508,\biu/cache_ctrl_logic/l1i_pte [60]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5691|biu/bus_unit/mmu/reg3_b60  (
    .a({open_n34509,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [60],\biu/bus_unit/mmu_hwdata [60]}),
    .clk(clk_pad),
    .d({_al_u5690_o,hrdata_pad[60]}),
    .sr(rst_pad),
    .f({hwdata_pad[60],open_n34527}),
    .q({open_n34531,\biu/bus_unit/mmu_hwdata [60]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5694|biu/cache_ctrl_logic/reg2_b59  (
    .a({open_n34532,_al_u2705_o}),
    .b({_al_u5693_o,_al_u5692_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4254_o,\biu/cache_ctrl_logic/pte_temp [59]}),
    .mi({open_n34543,\biu/cache_ctrl_logic/pte_temp [59]}),
    .sr(rst_pad),
    .f({_al_u5694_o,_al_u5693_o}),
    .q({open_n34547,\biu/cache_ctrl_logic/l1i_pte [59]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5695|biu/bus_unit/mmu/reg3_b59  (
    .a({open_n34548,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [59],\biu/bus_unit/mmu_hwdata [59]}),
    .clk(clk_pad),
    .d({_al_u5694_o,hrdata_pad[59]}),
    .sr(rst_pad),
    .f({hwdata_pad[59],open_n34566}),
    .q({open_n34570,\biu/bus_unit/mmu_hwdata [59]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5698|biu/cache_ctrl_logic/reg2_b58  (
    .a({open_n34571,_al_u2705_o}),
    .b({_al_u5697_o,_al_u5696_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4258_o,\biu/cache_ctrl_logic/pte_temp [58]}),
    .mi({open_n34575,\biu/cache_ctrl_logic/pte_temp [58]}),
    .sr(rst_pad),
    .f({_al_u5698_o,_al_u5697_o}),
    .q({open_n34590,\biu/cache_ctrl_logic/l1i_pte [58]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5699|biu/bus_unit/mmu/reg3_b58  (
    .a({open_n34591,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [58],\biu/bus_unit/mmu_hwdata [58]}),
    .clk(clk_pad),
    .d({_al_u5698_o,hrdata_pad[58]}),
    .sr(rst_pad),
    .f({hwdata_pad[58],open_n34605}),
    .q({open_n34609,\biu/bus_unit/mmu_hwdata [58]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5701|biu/cache_ctrl_logic/reg2_b57  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u5700_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [57]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [57],\biu/cache_ctrl_logic/pte_temp [57]}),
    .mi({open_n34620,\biu/cache_ctrl_logic/pte_temp [57]}),
    .sr(rst_pad),
    .f({_al_u5701_o,_al_u5700_o}),
    .q({open_n34624,\biu/cache_ctrl_logic/l1i_pte [57]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5703|biu/bus_unit/mmu/reg3_b57  (
    .a({open_n34625,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [57],\biu/bus_unit/mmu_hwdata [57]}),
    .clk(clk_pad),
    .d({_al_u5702_o,hrdata_pad[57]}),
    .sr(rst_pad),
    .f({hwdata_pad[57],open_n34639}),
    .q({open_n34643,\biu/bus_unit/mmu_hwdata [57]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5706|biu/cache_ctrl_logic/reg2_b56  (
    .a({open_n34644,_al_u2705_o}),
    .b({_al_u5705_o,_al_u5704_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4266_o,\biu/cache_ctrl_logic/pte_temp [56]}),
    .mi({open_n34648,\biu/cache_ctrl_logic/pte_temp [56]}),
    .sr(rst_pad),
    .f({_al_u5706_o,_al_u5705_o}),
    .q({open_n34663,\biu/cache_ctrl_logic/l1i_pte [56]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5707|biu/bus_unit/mmu/reg3_b56  (
    .a({open_n34664,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [56],\biu/bus_unit/mmu_hwdata [56]}),
    .clk(clk_pad),
    .d({_al_u5706_o,hrdata_pad[56]}),
    .sr(rst_pad),
    .f({hwdata_pad[56],open_n34682}),
    .q({open_n34686,\biu/bus_unit/mmu_hwdata [56]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5709|biu/cache_ctrl_logic/reg2_b55  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u5708_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [55]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [55],\biu/cache_ctrl_logic/pte_temp [55]}),
    .mi({open_n34697,\biu/cache_ctrl_logic/pte_temp [55]}),
    .sr(rst_pad),
    .f({_al_u5709_o,_al_u5708_o}),
    .q({open_n34701,\biu/cache_ctrl_logic/l1i_pte [55]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5711|biu/bus_unit/mmu/reg3_b55  (
    .a({open_n34702,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [55],\biu/bus_unit/mmu_hwdata [55]}),
    .clk(clk_pad),
    .d({_al_u5710_o,hrdata_pad[55]}),
    .sr(rst_pad),
    .f({hwdata_pad[55],open_n34720}),
    .q({open_n34724,\biu/bus_unit/mmu_hwdata [55]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5714|biu/cache_ctrl_logic/reg5_b54  (
    .a({open_n34725,_al_u2705_o}),
    .b({_al_u5713_o,_al_u5712_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4274_o,\biu/cache_ctrl_logic/l1d_pte [54]}),
    .mi({open_n34729,\biu/cache_ctrl_logic/pte_temp [54]}),
    .sr(rst_pad),
    .f({_al_u5714_o,_al_u5713_o}),
    .q({open_n34744,\biu/cache_ctrl_logic/l1d_pte [54]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5715|biu/bus_unit/mmu/reg3_b54  (
    .a({open_n34745,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [54],\biu/bus_unit/mmu_hwdata [54]}),
    .clk(clk_pad),
    .d({_al_u5714_o,hrdata_pad[54]}),
    .sr(rst_pad),
    .f({hwdata_pad[54],open_n34759}),
    .q({open_n34763,\biu/bus_unit/mmu_hwdata [54]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5718|biu/cache_ctrl_logic/reg5_b53  (
    .a({open_n34764,_al_u2705_o}),
    .b({_al_u5717_o,_al_u5716_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4278_o,\biu/cache_ctrl_logic/l1d_pte [53]}),
    .mi({open_n34775,\biu/cache_ctrl_logic/pte_temp [53]}),
    .sr(rst_pad),
    .f({_al_u5718_o,_al_u5717_o}),
    .q({open_n34779,\biu/cache_ctrl_logic/l1d_pte [53]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5719|biu/bus_unit/mmu/reg2_b55  (
    .b({_al_u2705_o,open_n34782}),
    .c({\biu/bus_unit/mmu_hwdata [53],_al_u3044_o}),
    .clk(clk_pad),
    .d({_al_u5718_o,_al_u3043_o}),
    .sr(rst_pad),
    .f({hwdata_pad[53],open_n34800}),
    .q({open_n34804,\biu/paddress [119]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5722|biu/cache_ctrl_logic/reg2_b52  (
    .a({open_n34805,_al_u2705_o}),
    .b({_al_u5721_o,_al_u5720_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4282_o,\biu/cache_ctrl_logic/pte_temp [52]}),
    .mi({open_n34816,\biu/cache_ctrl_logic/pte_temp [52]}),
    .sr(rst_pad),
    .f({_al_u5722_o,_al_u5721_o}),
    .q({open_n34820,\biu/cache_ctrl_logic/l1i_pte [52]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5726|biu/cache_ctrl_logic/reg5_b51  (
    .a({open_n34821,_al_u2705_o}),
    .b({_al_u5725_o,_al_u5724_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4286_o,\biu/cache_ctrl_logic/l1d_pte [51]}),
    .mi({open_n34832,\biu/cache_ctrl_logic/pte_temp [51]}),
    .sr(rst_pad),
    .f({_al_u5726_o,_al_u5725_o}),
    .q({open_n34836,\biu/cache_ctrl_logic/l1d_pte [51]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5729|biu/cache_ctrl_logic/reg2_b50  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u5728_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [50]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [50],\biu/cache_ctrl_logic/pte_temp [50]}),
    .mi({open_n34840,\biu/cache_ctrl_logic/pte_temp [50]}),
    .sr(rst_pad),
    .f({_al_u5729_o,_al_u5728_o}),
    .q({open_n34855,\biu/cache_ctrl_logic/l1i_pte [50]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5731|biu/bus_unit/mmu/reg1_b52  (
    .b({_al_u2705_o,open_n34858}),
    .c({\biu/bus_unit/mmu_hwdata [50],_al_u5029_o}),
    .clk(clk_pad),
    .d({_al_u5730_o,_al_u5028_o}),
    .sr(rst_pad),
    .f({hwdata_pad[50],open_n34872}),
    .q({open_n34876,\biu/paddress [52]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5734|biu/cache_ctrl_logic/reg2_b49  (
    .a({open_n34877,_al_u2705_o}),
    .b({_al_u5733_o,_al_u5732_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4294_o,\biu/cache_ctrl_logic/pte_temp [49]}),
    .mi({open_n34881,\biu/cache_ctrl_logic/pte_temp [49]}),
    .sr(rst_pad),
    .f({_al_u5734_o,_al_u5733_o}),
    .q({open_n34896,\biu/cache_ctrl_logic/l1i_pte [49]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5738|biu/cache_ctrl_logic/reg2_b48  (
    .a({open_n34897,_al_u2705_o}),
    .b({_al_u5737_o,_al_u5736_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4298_o,\biu/cache_ctrl_logic/pte_temp [48]}),
    .mi({open_n34901,\biu/cache_ctrl_logic/pte_temp [48]}),
    .sr(rst_pad),
    .f({_al_u5738_o,_al_u5737_o}),
    .q({open_n34916,\biu/cache_ctrl_logic/l1i_pte [48]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5739|biu/bus_unit/mmu/reg1_b50  (
    .b({_al_u2705_o,open_n34919}),
    .c({\biu/bus_unit/mmu_hwdata [48],_al_u5035_o}),
    .clk(clk_pad),
    .d({_al_u5738_o,_al_u5034_o}),
    .sr(rst_pad),
    .f({hwdata_pad[48],open_n34937}),
    .q({open_n34941,\biu/paddress [50]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5741|biu/cache_ctrl_logic/reg2_b47  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u5740_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [47]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [47],\biu/cache_ctrl_logic/pte_temp [47]}),
    .mi({open_n34945,\biu/cache_ctrl_logic/pte_temp [47]}),
    .sr(rst_pad),
    .f({_al_u5741_o,_al_u5740_o}),
    .q({open_n34960,\biu/cache_ctrl_logic/l1i_pte [47]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u5742|_al_u5743  (
    .b({_al_u5741_o,_al_u2705_o}),
    .c({_al_u3222_o,\biu/bus_unit/mmu_hwdata [47]}),
    .d({_al_u4302_o,_al_u5742_o}),
    .f({_al_u5742_o,hwdata_pad[47]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5746|biu/cache_ctrl_logic/reg2_b46  (
    .a({open_n34983,_al_u2705_o}),
    .b({_al_u5745_o,_al_u5744_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4306_o,\biu/cache_ctrl_logic/pte_temp [46]}),
    .mi({open_n34994,\biu/cache_ctrl_logic/pte_temp [46]}),
    .sr(rst_pad),
    .f({_al_u5746_o,_al_u5745_o}),
    .q({open_n34998,\biu/cache_ctrl_logic/l1i_pte [46]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5749|biu/cache_ctrl_logic/reg2_b45  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u5748_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [45]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [45],\biu/cache_ctrl_logic/pte_temp [45]}),
    .mi({open_n35009,\biu/cache_ctrl_logic/pte_temp [45]}),
    .sr(rst_pad),
    .f({_al_u5749_o,_al_u5748_o}),
    .q({open_n35013,\biu/cache_ctrl_logic/l1i_pte [45]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5750|_al_u5751  (
    .b({_al_u5749_o,_al_u2705_o}),
    .c({_al_u3222_o,\biu/bus_unit/mmu_hwdata [45]}),
    .d({_al_u4310_o,_al_u5750_o}),
    .f({_al_u5750_o,hwdata_pad[45]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5754|biu/cache_ctrl_logic/reg5_b44  (
    .a({open_n35040,_al_u2705_o}),
    .b({_al_u5753_o,_al_u5752_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4314_o,\biu/cache_ctrl_logic/l1d_pte [44]}),
    .mi({open_n35044,\biu/cache_ctrl_logic/pte_temp [44]}),
    .sr(rst_pad),
    .f({_al_u5754_o,_al_u5753_o}),
    .q({open_n35059,\biu/cache_ctrl_logic/l1d_pte [44]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5758|biu/cache_ctrl_logic/reg2_b43  (
    .a({open_n35060,_al_u2705_o}),
    .b({_al_u5757_o,_al_u5756_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4318_o,\biu/cache_ctrl_logic/pte_temp [43]}),
    .mi({open_n35071,\biu/cache_ctrl_logic/pte_temp [43]}),
    .sr(rst_pad),
    .f({_al_u5758_o,_al_u5757_o}),
    .q({open_n35075,\biu/cache_ctrl_logic/l1i_pte [43]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5762|biu/cache_ctrl_logic/reg2_b42  (
    .a({open_n35076,_al_u2705_o}),
    .b({_al_u5761_o,_al_u5760_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4322_o,\biu/cache_ctrl_logic/pte_temp [42]}),
    .mi({open_n35080,\biu/cache_ctrl_logic/pte_temp [42]}),
    .sr(rst_pad),
    .f({_al_u5762_o,_al_u5761_o}),
    .q({open_n35095,\biu/cache_ctrl_logic/l1i_pte [42]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5766|biu/cache_ctrl_logic/reg2_b41  (
    .a({open_n35096,_al_u2705_o}),
    .b({_al_u5765_o,_al_u5764_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4326_o,\biu/cache_ctrl_logic/pte_temp [41]}),
    .mi({open_n35100,\biu/cache_ctrl_logic/pte_temp [41]}),
    .sr(rst_pad),
    .f({_al_u5766_o,_al_u5765_o}),
    .q({open_n35115,\biu/cache_ctrl_logic/l1i_pte [41]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5770|biu/cache_ctrl_logic/reg5_b40  (
    .a({open_n35116,_al_u2705_o}),
    .b({_al_u5769_o,_al_u5768_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4330_o,\biu/cache_ctrl_logic/l1d_pte [40]}),
    .mi({open_n35120,\biu/cache_ctrl_logic/pte_temp [40]}),
    .sr(rst_pad),
    .f({_al_u5770_o,_al_u5769_o}),
    .q({open_n35135,\biu/cache_ctrl_logic/l1d_pte [40]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5774|biu/cache_ctrl_logic/reg2_b39  (
    .a({open_n35136,_al_u2705_o}),
    .b({_al_u5773_o,_al_u5772_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4334_o,\biu/cache_ctrl_logic/pte_temp [39]}),
    .mi({open_n35147,\biu/cache_ctrl_logic/pte_temp [39]}),
    .sr(rst_pad),
    .f({_al_u5774_o,_al_u5773_o}),
    .q({open_n35151,\biu/cache_ctrl_logic/l1i_pte [39]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5775|biu/bus_unit/mmu/reg1_b41  (
    .b({_al_u2705_o,open_n35154}),
    .c({\biu/bus_unit/mmu_hwdata [39],_al_u5062_o}),
    .clk(clk_pad),
    .d({_al_u5774_o,_al_u5061_o}),
    .sr(rst_pad),
    .f({hwdata_pad[39],open_n35168}),
    .q({open_n35172,\biu/paddress [41]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5778|biu/cache_ctrl_logic/reg2_b38  (
    .a({open_n35173,_al_u2705_o}),
    .b({_al_u5777_o,_al_u5776_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4338_o,\biu/cache_ctrl_logic/pte_temp [38]}),
    .mi({open_n35184,\biu/cache_ctrl_logic/pte_temp [38]}),
    .sr(rst_pad),
    .f({_al_u5778_o,_al_u5777_o}),
    .q({open_n35188,\biu/cache_ctrl_logic/l1i_pte [38]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5779|biu/bus_unit/mmu/reg1_b40  (
    .b({_al_u2705_o,open_n35191}),
    .c({\biu/bus_unit/mmu_hwdata [38],_al_u5065_o}),
    .clk(clk_pad),
    .d({_al_u5778_o,_al_u5064_o}),
    .sr(rst_pad),
    .f({hwdata_pad[38],open_n35205}),
    .q({open_n35209,\biu/paddress [40]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5782|biu/cache_ctrl_logic/reg2_b37  (
    .a({open_n35210,_al_u2705_o}),
    .b({_al_u5781_o,_al_u5780_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4342_o,\biu/cache_ctrl_logic/pte_temp [37]}),
    .mi({open_n35214,\biu/cache_ctrl_logic/pte_temp [37]}),
    .sr(rst_pad),
    .f({_al_u5782_o,_al_u5781_o}),
    .q({open_n35229,\biu/cache_ctrl_logic/l1i_pte [37]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5786|biu/cache_ctrl_logic/reg5_b36  (
    .a({open_n35230,_al_u2705_o}),
    .b({_al_u5785_o,_al_u5784_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4346_o,\biu/cache_ctrl_logic/l1d_pte [36]}),
    .mi({open_n35241,\biu/cache_ctrl_logic/pte_temp [36]}),
    .sr(rst_pad),
    .f({_al_u5786_o,_al_u5785_o}),
    .q({open_n35245,\biu/cache_ctrl_logic/l1d_pte [36]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5790|biu/cache_ctrl_logic/reg5_b35  (
    .a({open_n35246,_al_u2705_o}),
    .b({_al_u5789_o,_al_u5788_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4350_o,\biu/cache_ctrl_logic/l1d_pte [35]}),
    .mi({open_n35257,\biu/cache_ctrl_logic/pte_temp [35]}),
    .sr(rst_pad),
    .f({_al_u5790_o,_al_u5789_o}),
    .q({open_n35261,\biu/cache_ctrl_logic/l1d_pte [35]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5791|biu/bus_unit/mmu/reg1_b37  (
    .b({_al_u2705_o,open_n35264}),
    .c({\biu/bus_unit/mmu_hwdata [35],_al_u5074_o}),
    .clk(clk_pad),
    .d({_al_u5790_o,_al_u5073_o}),
    .sr(rst_pad),
    .f({hwdata_pad[35],open_n35278}),
    .q({open_n35282,\biu/paddress [37]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5794|biu/cache_ctrl_logic/reg2_b34  (
    .a({open_n35283,_al_u2705_o}),
    .b({_al_u5793_o,_al_u5792_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4354_o,\biu/cache_ctrl_logic/pte_temp [34]}),
    .mi({open_n35287,\biu/cache_ctrl_logic/pte_temp [34]}),
    .sr(rst_pad),
    .f({_al_u5794_o,_al_u5793_o}),
    .q({open_n35302,\biu/cache_ctrl_logic/l1i_pte [34]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5795|biu/bus_unit/mmu/reg1_b36  (
    .b({_al_u2705_o,open_n35305}),
    .c({\biu/bus_unit/mmu_hwdata [34],_al_u5077_o}),
    .clk(clk_pad),
    .d({_al_u5794_o,_al_u5076_o}),
    .sr(rst_pad),
    .f({hwdata_pad[34],open_n35319}),
    .q({open_n35323,\biu/paddress [36]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5798|biu/cache_ctrl_logic/reg2_b33  (
    .a({open_n35324,_al_u2705_o}),
    .b({_al_u5797_o,_al_u5796_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4358_o,\biu/cache_ctrl_logic/pte_temp [33]}),
    .mi({open_n35335,\biu/cache_ctrl_logic/pte_temp [33]}),
    .sr(rst_pad),
    .f({_al_u5798_o,_al_u5797_o}),
    .q({open_n35339,\biu/cache_ctrl_logic/l1i_pte [33]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5799|biu/bus_unit/mmu/reg1_b35  (
    .b({_al_u2705_o,open_n35342}),
    .c({\biu/bus_unit/mmu_hwdata [33],_al_u5080_o}),
    .clk(clk_pad),
    .d({_al_u5798_o,_al_u5079_o}),
    .sr(rst_pad),
    .f({hwdata_pad[33],open_n35360}),
    .q({open_n35364,\biu/paddress [35]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5802|biu/cache_ctrl_logic/reg5_b32  (
    .a({open_n35365,_al_u2705_o}),
    .b({_al_u5801_o,_al_u5800_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4362_o,\biu/cache_ctrl_logic/l1d_pte [32]}),
    .mi({open_n35369,\biu/cache_ctrl_logic/pte_temp [32]}),
    .sr(rst_pad),
    .f({_al_u5802_o,_al_u5801_o}),
    .q({open_n35384,\biu/cache_ctrl_logic/l1d_pte [32]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5805|biu/cache_ctrl_logic/reg2_b31  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u5804_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [31]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [31],\biu/cache_ctrl_logic/pte_temp [31]}),
    .mi({open_n35395,\biu/cache_ctrl_logic/pte_temp [31]}),
    .sr(rst_pad),
    .f({_al_u5805_o,_al_u5804_o}),
    .q({open_n35399,\biu/cache_ctrl_logic/l1i_pte [31]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5807|biu/bus_unit/mmu/reg1_b33  (
    .b({_al_u2705_o,open_n35402}),
    .c({\biu/bus_unit/mmu_hwdata [31],_al_u5086_o}),
    .clk(clk_pad),
    .d({_al_u5806_o,_al_u5085_o}),
    .sr(rst_pad),
    .f({hwdata_pad[31],open_n35416}),
    .q({open_n35420,\biu/paddress [33]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5810|biu/cache_ctrl_logic/reg2_b30  (
    .a({open_n35421,_al_u2705_o}),
    .b({_al_u5809_o,_al_u5808_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4370_o,\biu/cache_ctrl_logic/pte_temp [30]}),
    .mi({open_n35432,\biu/cache_ctrl_logic/pte_temp [30]}),
    .sr(rst_pad),
    .f({_al_u5810_o,_al_u5809_o}),
    .q({open_n35436,\biu/cache_ctrl_logic/l1i_pte [30]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5811|biu/bus_unit/mmu/reg1_b32  (
    .b({_al_u2705_o,open_n35439}),
    .c({\biu/bus_unit/mmu_hwdata [30],_al_u5089_o}),
    .clk(clk_pad),
    .d({_al_u5810_o,_al_u5088_o}),
    .sr(rst_pad),
    .f({hwdata_pad[30],open_n35453}),
    .q({open_n35457,\biu/paddress [32]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5814|biu/cache_ctrl_logic/reg2_b29  (
    .a({open_n35458,_al_u2705_o}),
    .b({_al_u5813_o,_al_u5812_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4374_o,\biu/cache_ctrl_logic/pte_temp [29]}),
    .mi({open_n35462,\biu/cache_ctrl_logic/pte_temp [29]}),
    .sr(rst_pad),
    .f({_al_u5814_o,_al_u5813_o}),
    .q({open_n35477,\biu/cache_ctrl_logic/l1i_pte [29]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5815|biu/bus_unit/mmu/reg1_b31  (
    .b({_al_u2705_o,open_n35480}),
    .c({\biu/bus_unit/mmu_hwdata [29],_al_u5092_o}),
    .clk(clk_pad),
    .d({_al_u5814_o,_al_u5091_o}),
    .sr(rst_pad),
    .f({hwdata_pad[29],open_n35494}),
    .q({open_n35498,\biu/paddress [31]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5817|biu/cache_ctrl_logic/reg2_b28  (
    .a({_al_u2705_o,_al_u3945_o}),
    .b({_al_u5816_o,_al_u3947_o}),
    .c({_al_u3950_o,\biu/cache_ctrl_logic/l1d_pte [28]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_pte [28],\biu/cache_ctrl_logic/pte_temp [28]}),
    .mi({open_n35502,\biu/cache_ctrl_logic/pte_temp [28]}),
    .sr(rst_pad),
    .f({_al_u5817_o,_al_u5816_o}),
    .q({open_n35517,\biu/cache_ctrl_logic/l1i_pte [28]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(B*~(~C*~D))"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"))
    \_al_u5818|_al_u5819  (
    .b({_al_u5817_o,_al_u2705_o}),
    .c({_al_u3222_o,\biu/bus_unit/mmu_hwdata [28]}),
    .d({_al_u4378_o,_al_u5818_o}),
    .f({_al_u5818_o,hwdata_pad[28]}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5822|biu/cache_ctrl_logic/reg2_b27  (
    .a({open_n35540,_al_u2705_o}),
    .b({_al_u5821_o,_al_u5820_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4382_o,\biu/cache_ctrl_logic/pte_temp [27]}),
    .mi({open_n35544,\biu/cache_ctrl_logic/pte_temp [27]}),
    .sr(rst_pad),
    .f({_al_u5822_o,_al_u5821_o}),
    .q({open_n35559,\biu/cache_ctrl_logic/l1i_pte [27]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5823|biu/bus_unit/mmu/reg3_b27  (
    .a({open_n35560,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [27],\biu/bus_unit/mmu_hwdata [27]}),
    .clk(clk_pad),
    .d({_al_u5822_o,hrdata_pad[27]}),
    .sr(rst_pad),
    .f({hwdata_pad[27],open_n35578}),
    .q({open_n35582,\biu/bus_unit/mmu_hwdata [27]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*C))"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(B*~A*~(D*C))"),
    //.LUTG1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010001000100),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000010001000100),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5826|biu/cache_ctrl_logic/reg5_b26  (
    .a({open_n35583,_al_u2705_o}),
    .b({_al_u5825_o,_al_u5824_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4386_o,\biu/cache_ctrl_logic/l1d_pte [26]}),
    .mi({open_n35587,\biu/cache_ctrl_logic/pte_temp [26]}),
    .sr(rst_pad),
    .f({_al_u5826_o,_al_u5825_o}),
    .q({open_n35602,\biu/cache_ctrl_logic/l1d_pte [26]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111010111010),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111111010111010),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5827|biu/bus_unit/mmu/reg3_b26  (
    .a({open_n35603,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [26],\biu/bus_unit/mmu_hwdata [26]}),
    .clk(clk_pad),
    .d({_al_u5826_o,hrdata_pad[26]}),
    .sr(rst_pad),
    .f({hwdata_pad[26],open_n35621}),
    .q({open_n35625,\biu/bus_unit/mmu_hwdata [26]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5830|biu/cache_ctrl_logic/reg5_b25  (
    .a({open_n35626,_al_u2705_o}),
    .b({_al_u5829_o,_al_u5828_o}),
    .c({_al_u3222_o,_al_u3947_o}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u4390_o,\biu/cache_ctrl_logic/l1d_pte [25]}),
    .mi({open_n35637,\biu/cache_ctrl_logic/pte_temp [25]}),
    .sr(rst_pad),
    .f({_al_u5830_o,_al_u5829_o}),
    .q({open_n35641,\biu/cache_ctrl_logic/l1d_pte [25]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5831|biu/bus_unit/mmu/reg3_b25  (
    .a({open_n35642,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [25],\biu/bus_unit/mmu_hwdata [25]}),
    .clk(clk_pad),
    .d({_al_u5830_o,hrdata_pad[25]}),
    .sr(rst_pad),
    .f({hwdata_pad[25],open_n35656}),
    .q({open_n35660,\biu/bus_unit/mmu_hwdata [25]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(D*C))"),
    //.LUT1("(B*~(~C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010001000100),
    .INIT_LUT1(16'b1100110011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5834|biu/cache_ctrl_logic/reg2_b24  (
    .a({open_n35661,_al_u2705_o}),
    .b({_al_u5833_o,_al_u5832_o}),
    .c({_al_u3222_o,_al_u3945_o}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({_al_u4394_o,\biu/cache_ctrl_logic/pte_temp [24]}),
    .mi({open_n35672,\biu/cache_ctrl_logic/pte_temp [24]}),
    .sr(rst_pad),
    .f({_al_u5834_o,_al_u5833_o}),
    .q({open_n35676,\biu/cache_ctrl_logic/l1i_pte [24]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111010111010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5835|biu/bus_unit/mmu/reg3_b24  (
    .a({open_n35677,_al_u2963_o}),
    .b({_al_u2705_o,\biu/bus_unit/mmu/mux34_b0_sel_is_3_o }),
    .c({\biu/bus_unit/mmu_hwdata [24],\biu/bus_unit/mmu_hwdata [24]}),
    .clk(clk_pad),
    .d({_al_u5834_o,hrdata_pad[24]}),
    .sr(rst_pad),
    .f({hwdata_pad[24],open_n35691}),
    .q({open_n35695,\biu/bus_unit/mmu_hwdata [24]}));  // ../../RTL/CPU/BIU/mmu.v(218)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(~B*~(D*~C*A))"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(~B*~(D*~C*A))"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0011000100110011),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b0011000100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5836|_al_u4800  (
    .a({_al_u4092_o,_al_u4092_o}),
    .b({\ins_dec/ins_srai ,_al_u3216_o}),
    .c({_al_u3217_o,_al_u3217_o}),
    .d({_al_u3384_o,_al_u3384_o}),
    .f({\ins_dec/n57_neg_lutinv ,\ins_dec/ins_srli }));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5837|_al_u5847  (
    .a({_al_u5144_o,_al_u5144_o}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_005 ,\cu_ru/al_ram_gpr_al_u0_do_i0_000 }),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_005 ,\cu_ru/al_ram_gpr_al_u0_do_i1_000 }),
    .d({\cu_ru/n49 [4],\cu_ru/n49 [4]}),
    .f({_al_u5837_o,_al_u5847_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5839|_al_u5845  (
    .a({_al_u5144_o,_al_u5144_o}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_004 ,\cu_ru/al_ram_gpr_al_u0_do_i0_001 }),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_004 ,\cu_ru/al_ram_gpr_al_u0_do_i1_001 }),
    .d({\cu_ru/n49 [4],\cu_ru/n49 [4]}),
    .f({_al_u5839_o,_al_u5845_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"))
    \_al_u5841|_al_u5843  (
    .a({_al_u5144_o,_al_u5144_o}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_003 ,\cu_ru/al_ram_gpr_al_u0_do_i0_002 }),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_003 ,\cu_ru/al_ram_gpr_al_u0_do_i1_002 }),
    .d({\cu_ru/n49 [4],\cu_ru/n49 [4]}),
    .f({_al_u5841_o,_al_u5843_o}));
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5849|ins_dec/csr_write_reg  (
    .b({open_n35790,_al_u3217_o}),
    .c({_al_u3216_o,_al_u3384_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/n239 ,id_system}),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/mux19_b10_sel_is_2_o ,\ins_dec/n239 }),
    .q({open_n35806,ex_csr_write}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A*~(~C*~B))"),
    //.LUT1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010100),
    .INIT_LUT1(16'b0000011111110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5850|ins_dec/reg5_b9  (
    .a({rs1_data[9],_al_u7891_o}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,rs1_data[9]}),
    .c({_al_u3927_o,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[29],\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u5850_o,open_n35819}),
    .q({open_n35823,ds1[9]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011111100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0000110011111100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5851|ins_dec/reg6_b9  (
    .a({_al_u5143_o,open_n35824}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_009 ,_al_u5851_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_009 ,_al_u4086_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5850_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5851_o,open_n35841}),
    .q({open_n35845,ds2[9]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A*~(~C*~B))"),
    //.LUT1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010100),
    .INIT_LUT1(16'b0000011111110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5853|ins_dec/reg5_b8  (
    .a({rs1_data[8],_al_u7871_o}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,rs1_data[8]}),
    .c({_al_u3927_o,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[28],\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u5853_o,open_n35858}),
    .q({open_n35862,ds1[8]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011111100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5854|ins_dec/reg6_b8  (
    .a({_al_u5143_o,open_n35863}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_008 ,_al_u5854_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_008 ,_al_u4086_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5853_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5854_o,open_n35876}),
    .q({open_n35880,ds2[8]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A*~(~C*~B))"),
    //.LUT1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010100),
    .INIT_LUT1(16'b0000011111110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5856|ins_dec/reg5_b7  (
    .a({rs1_data[7],_al_u7836_o}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,rs1_data[7]}),
    .c({_al_u3927_o,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[27],\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u5856_o,open_n35893}),
    .q({open_n35897,ds1[7]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5858|_al_u7353  (
    .c({id_ins[31],id_ins[31]}),
    .d({_al_u3955_o,\ins_dec/op_lui_lutinv }),
    .f({_al_u5858_o,_al_u7353_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u5859|_al_u6100  (
    .b({_al_u5858_o,_al_u5858_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,\ins_dec/mux19_b10_sel_is_2_o }),
    .d({rs1_data[63],rs1_data[43]}),
    .f({_al_u5859_o,_al_u6100_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5860|ins_dec/reg6_b63  (
    .a({_al_u5144_o,open_n35944}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_063 ,open_n35945}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_063 ,_al_u5860_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5859_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5860_o,open_n35958}),
    .q({open_n35962,ds2[63]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u5862|_al_u5868  (
    .b({_al_u5858_o,_al_u5858_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,\ins_dec/mux19_b10_sel_is_2_o }),
    .d({rs1_data[62],rs1_data[60]}),
    .f({_al_u5862_o,_al_u5868_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5863|ins_dec/reg6_b62  (
    .a({_al_u5144_o,open_n35985}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_062 ,open_n35986}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_062 ,_al_u5863_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5862_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5863_o,open_n36003}),
    .q({open_n36007,ds2[62]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5866|ins_dec/reg6_b61  (
    .a({_al_u5144_o,open_n36008}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_061 ,open_n36009}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_061 ,_al_u5866_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5865_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5866_o,open_n36022}),
    .q({open_n36026,ds2[61]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5869|ins_dec/reg6_b60  (
    .a({_al_u5144_o,open_n36027}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_060 ,open_n36028}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_060 ,_al_u5869_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5868_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5869_o,open_n36041}),
    .q({open_n36045,ds2[60]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~A*~(~C*~B))"),
    //.LUTF1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    //.LUTG0("(~D*~A*~(~C*~B))"),
    //.LUTG1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000001010100),
    .INIT_LUTF1(16'b0000011111110111),
    .INIT_LUTG0(16'b0000000001010100),
    .INIT_LUTG1(16'b0000011111110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5871|ins_dec/reg5_b6  (
    .a({rs1_data[6],_al_u7814_o}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,rs1_data[6]}),
    .c({_al_u3927_o,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[26],\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u5871_o,open_n36062}),
    .q({open_n36066,ds1[6]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5873|ins_dec/reg7_b59  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[59]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[59],rs1_data[59]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5873_o,open_n36081}),
    .q({open_n36085,as1[59]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5874|ins_dec/reg6_b59  (
    .a({_al_u5144_o,open_n36086}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_059 ,open_n36087}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_059 ,_al_u5874_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5873_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5874_o,open_n36104}),
    .q({open_n36108,ds2[59]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5876|ins_dec/reg7_b58  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[58]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[58],rs1_data[58]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5876_o,open_n36127}),
    .q({open_n36131,as1[58]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5877|ins_dec/reg6_b58  (
    .a({_al_u5144_o,open_n36132}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_058 ,open_n36133}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_058 ,_al_u5877_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5876_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5877_o,open_n36150}),
    .q({open_n36154,ds2[58]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5879|ins_dec/reg7_b57  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[57]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[57],rs1_data[57]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5879_o,open_n36173}),
    .q({open_n36177,as1[57]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5880|ins_dec/reg6_b57  (
    .a({_al_u5144_o,open_n36178}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_057 ,open_n36179}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_057 ,_al_u5880_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5879_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5880_o,open_n36192}),
    .q({open_n36196,ds2[57]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5882|ins_dec/reg7_b56  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[56]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[56],rs1_data[56]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5882_o,open_n36211}),
    .q({open_n36215,as1[56]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5883|ins_dec/reg6_b56  (
    .a({_al_u5144_o,open_n36216}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_056 ,open_n36217}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_056 ,_al_u5883_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5882_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5883_o,open_n36230}),
    .q({open_n36234,ds2[56]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~A*~(~C*~B))"),
    //.LUTF1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    //.LUTG0("(~D*~A*~(~C*~B))"),
    //.LUTG1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000001010100),
    .INIT_LUTF1(16'b0000011111110111),
    .INIT_LUTG0(16'b0000000001010100),
    .INIT_LUTG1(16'b0000011111110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5885|ins_dec/reg5_b5  (
    .a({rs1_data[5],_al_u7895_o}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,rs1_data[5]}),
    .c({_al_u3927_o,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[25],\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u5885_o,open_n36251}),
    .q({open_n36255,ds1[5]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~A*~(~C*~B))"),
    //.LUTF1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    //.LUTG0("(~D*~A*~(~C*~B))"),
    //.LUTG1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000001010100),
    .INIT_LUTF1(16'b0000011111110111),
    .INIT_LUTG0(16'b0000000001010100),
    .INIT_LUTG1(16'b0000011111110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5887|ins_dec/reg5_b11  (
    .a({rs1_data[11],_al_u7834_o}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,rs1_data[11]}),
    .c({_al_u3927_o,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[31],\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u5887_o,open_n36272}),
    .q({open_n36276,ds1[11]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUT1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011111100),
    .INIT_LUT1(16'b0101000001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5888|ins_dec/reg6_b11  (
    .a({_al_u5143_o,open_n36277}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_011 ,_al_u5888_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_011 ,_al_u4086_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5887_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5888_o,open_n36290}),
    .q({open_n36294,ds2[11]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~A*~(~C*~B))"),
    //.LUTF1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    //.LUTG0("(~D*~A*~(~C*~B))"),
    //.LUTG1("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000001010100),
    .INIT_LUTF1(16'b0000011111110111),
    .INIT_LUTG0(16'b0000000001010100),
    .INIT_LUTG1(16'b0000011111110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5890|ins_dec/reg5_b10  (
    .a({rs1_data[10],_al_u7710_o}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,rs1_data[10]}),
    .c({_al_u3927_o,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[30],\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u5890_o,open_n36311}),
    .q({open_n36315,ds1[10]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTF1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG1("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011111100),
    .INIT_LUTF1(16'b0101000001000100),
    .INIT_LUTG0(16'b0000110011111100),
    .INIT_LUTG1(16'b0101000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5891|ins_dec/reg6_b10  (
    .a({_al_u5143_o,open_n36316}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_010 ,_al_u5891_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_010 ,_al_u4086_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u5890_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u5891_o,open_n36333}),
    .q({open_n36337,ds2[10]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0100110001111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0100110001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5893|biu/cache_ctrl_logic/reg6_b29  (
    .a({\biu/bus_unit/mmu/i [0],open_n36338}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [29]}),
    .c({\biu/paddress [29],\biu/cache_ctrl_logic/pa_temp [29]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [27],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5893_o,open_n36356}),
    .q({open_n36360,\biu/cache_ctrl_logic/pa_temp [29]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUTF1("(B*~(D*~C*A))"),
    //.LUTG0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUTG1("(B*~(D*~C*A))"),
    .INIT_LUTF0(16'b0010000000100011),
    .INIT_LUTF1(16'b1100010011001100),
    .INIT_LUTG0(16'b0010000000100011),
    .INIT_LUTG1(16'b1100010011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5894|_al_u5895  (
    .a({\biu/maddress [29],_al_u5894_o}),
    .b({_al_u5893_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [29]}),
    .f({_al_u5894_o,_al_u5895_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5896|biu/bus_unit/mmu/reg1_b29  (
    .a({\biu/maddress [29],open_n36385}),
    .b({_al_u2914_o,open_n36386}),
    .c({_al_u2698_o,_al_u5896_o}),
    .clk(clk_pad),
    .d({\biu/paddress [29],_al_u5895_o}),
    .sr(rst_pad),
    .f({_al_u5896_o,open_n36404}),
    .q({open_n36408,\biu/paddress [29]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0100110001111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0100110001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5898|biu/cache_ctrl_logic/reg6_b28  (
    .a({\biu/bus_unit/mmu/i [0],open_n36409}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [28]}),
    .c({\biu/paddress [28],\biu/cache_ctrl_logic/pa_temp [28]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [26],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5898_o,open_n36427}),
    .q({open_n36431,\biu/cache_ctrl_logic/pa_temp [28]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUT1("(B*~(D*~C*A))"),
    .INIT_LUT0(16'b0010000000100011),
    .INIT_LUT1(16'b1100010011001100),
    .MODE("LOGIC"))
    \_al_u5899|_al_u5900  (
    .a({\biu/maddress [28],_al_u5899_o}),
    .b({_al_u5898_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [28]}),
    .f({_al_u5899_o,_al_u5900_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5901|biu/bus_unit/mmu/reg1_b28  (
    .a({\biu/maddress [28],open_n36452}),
    .b({_al_u2914_o,open_n36453}),
    .c({_al_u2698_o,_al_u5901_o}),
    .clk(clk_pad),
    .d({\biu/paddress [28],_al_u5900_o}),
    .sr(rst_pad),
    .f({_al_u5901_o,open_n36471}),
    .q({open_n36475,\biu/paddress [28]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0100110001111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5903|biu/cache_ctrl_logic/reg6_b27  (
    .a({\biu/bus_unit/mmu/i [0],open_n36476}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [27]}),
    .c({\biu/paddress [27],\biu/cache_ctrl_logic/pa_temp [27]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [25],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5903_o,open_n36490}),
    .q({open_n36494,\biu/cache_ctrl_logic/pa_temp [27]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUT1("(B*~(D*~C*A))"),
    .INIT_LUT0(16'b0010000000100011),
    .INIT_LUT1(16'b1100010011001100),
    .MODE("LOGIC"))
    \_al_u5904|_al_u5905  (
    .a({\biu/maddress [27],_al_u5904_o}),
    .b({_al_u5903_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [27]}),
    .f({_al_u5904_o,_al_u5905_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5906|biu/bus_unit/mmu/reg1_b27  (
    .a({\biu/maddress [27],open_n36515}),
    .b({_al_u2914_o,open_n36516}),
    .c({_al_u2698_o,_al_u5906_o}),
    .clk(clk_pad),
    .d({\biu/paddress [27],_al_u5905_o}),
    .sr(rst_pad),
    .f({_al_u5906_o,open_n36530}),
    .q({open_n36534,\biu/paddress [27]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0100110001111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5908|biu/cache_ctrl_logic/reg6_b26  (
    .a({\biu/bus_unit/mmu/i [0],open_n36535}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [26]}),
    .c({\biu/paddress [26],\biu/cache_ctrl_logic/pa_temp [26]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [24],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5908_o,open_n36549}),
    .q({open_n36553,\biu/cache_ctrl_logic/pa_temp [26]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUTF1("(B*~(D*~C*A))"),
    //.LUTG0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUTG1("(B*~(D*~C*A))"),
    .INIT_LUTF0(16'b0010000000100011),
    .INIT_LUTF1(16'b1100010011001100),
    .INIT_LUTG0(16'b0010000000100011),
    .INIT_LUTG1(16'b1100010011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5909|_al_u5910  (
    .a({\biu/maddress [26],_al_u5909_o}),
    .b({_al_u5908_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [26]}),
    .f({_al_u5909_o,_al_u5910_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5911|biu/bus_unit/mmu/reg1_b26  (
    .a({\biu/maddress [26],open_n36578}),
    .b({_al_u2914_o,open_n36579}),
    .c({_al_u2698_o,_al_u5911_o}),
    .clk(clk_pad),
    .d({\biu/paddress [26],_al_u5910_o}),
    .sr(rst_pad),
    .f({_al_u5911_o,open_n36593}),
    .q({open_n36597,\biu/paddress [26]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0100110001111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0100110001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5913|biu/cache_ctrl_logic/reg6_b25  (
    .a({\biu/bus_unit/mmu/i [0],open_n36598}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [25]}),
    .c({\biu/paddress [25],\biu/cache_ctrl_logic/pa_temp [25]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [23],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5913_o,open_n36616}),
    .q({open_n36620,\biu/cache_ctrl_logic/pa_temp [25]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUTF1("(B*~(D*~C*A))"),
    //.LUTG0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUTG1("(B*~(D*~C*A))"),
    .INIT_LUTF0(16'b0010000000100011),
    .INIT_LUTF1(16'b1100010011001100),
    .INIT_LUTG0(16'b0010000000100011),
    .INIT_LUTG1(16'b1100010011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5914|_al_u5915  (
    .a({\biu/maddress [25],_al_u5914_o}),
    .b({_al_u5913_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [25]}),
    .f({_al_u5914_o,_al_u5915_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5916|biu/bus_unit/mmu/reg1_b25  (
    .a({\biu/maddress [25],open_n36645}),
    .b({_al_u2914_o,open_n36646}),
    .c({_al_u2698_o,_al_u5916_o}),
    .clk(clk_pad),
    .d({\biu/paddress [25],_al_u5915_o}),
    .sr(rst_pad),
    .f({_al_u5916_o,open_n36664}),
    .q({open_n36668,\biu/paddress [25]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0100110001111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0100110001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5918|biu/cache_ctrl_logic/reg6_b24  (
    .a({\biu/bus_unit/mmu/i [0],open_n36669}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [24]}),
    .c({\biu/paddress [24],\biu/cache_ctrl_logic/pa_temp [24]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [22],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5918_o,open_n36687}),
    .q({open_n36691,\biu/cache_ctrl_logic/pa_temp [24]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUT1("(B*~(D*~C*A))"),
    .INIT_LUT0(16'b0010000000100011),
    .INIT_LUT1(16'b1100010011001100),
    .MODE("LOGIC"))
    \_al_u5919|_al_u5920  (
    .a({\biu/maddress [24],_al_u5919_o}),
    .b({_al_u5918_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [24]}),
    .f({_al_u5919_o,_al_u5920_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5921|biu/bus_unit/mmu/reg1_b24  (
    .a({\biu/maddress [24],open_n36712}),
    .b({_al_u2914_o,open_n36713}),
    .c({_al_u2698_o,_al_u5921_o}),
    .clk(clk_pad),
    .d({\biu/paddress [24],_al_u5920_o}),
    .sr(rst_pad),
    .f({_al_u5921_o,open_n36731}),
    .q({open_n36735,\biu/paddress [24]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0100110001111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5923|biu/cache_ctrl_logic/reg6_b23  (
    .a({\biu/bus_unit/mmu/i [0],open_n36736}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [23]}),
    .c({\biu/paddress [23],\biu/cache_ctrl_logic/pa_temp [23]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [21],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5923_o,open_n36750}),
    .q({open_n36754,\biu/cache_ctrl_logic/pa_temp [23]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUT1("(B*~(D*~C*A))"),
    .INIT_LUT0(16'b0010000000100011),
    .INIT_LUT1(16'b1100010011001100),
    .MODE("LOGIC"))
    \_al_u5924|_al_u5925  (
    .a({\biu/maddress [23],_al_u5924_o}),
    .b({_al_u5923_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [23]}),
    .f({_al_u5924_o,_al_u5925_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5926|biu/bus_unit/mmu/reg1_b23  (
    .a({\biu/maddress [23],open_n36775}),
    .b({_al_u2914_o,open_n36776}),
    .c({_al_u2698_o,_al_u5926_o}),
    .clk(clk_pad),
    .d({\biu/paddress [23],_al_u5925_o}),
    .sr(rst_pad),
    .f({_al_u5926_o,open_n36790}),
    .q({open_n36794,\biu/paddress [23]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0100110001111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5928|biu/cache_ctrl_logic/reg6_b22  (
    .a({\biu/bus_unit/mmu/i [0],open_n36795}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [22]}),
    .c({\biu/paddress [22],\biu/cache_ctrl_logic/pa_temp [22]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [20],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5928_o,open_n36809}),
    .q({open_n36813,\biu/cache_ctrl_logic/pa_temp [22]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUTF1("(B*~(D*~C*A))"),
    //.LUTG0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUTG1("(B*~(D*~C*A))"),
    .INIT_LUTF0(16'b0010000000100011),
    .INIT_LUTF1(16'b1100010011001100),
    .INIT_LUTG0(16'b0010000000100011),
    .INIT_LUTG1(16'b1100010011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5929|_al_u5930  (
    .a({\biu/maddress [22],_al_u5929_o}),
    .b({_al_u5928_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [22]}),
    .f({_al_u5929_o,_al_u5930_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5931|biu/bus_unit/mmu/reg1_b22  (
    .a({\biu/maddress [22],open_n36838}),
    .b({_al_u2914_o,open_n36839}),
    .c({_al_u2698_o,_al_u5931_o}),
    .clk(clk_pad),
    .d({\biu/paddress [22],_al_u5930_o}),
    .sr(rst_pad),
    .f({_al_u5931_o,open_n36853}),
    .q({open_n36857,\biu/paddress [22]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0100110001111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0100110001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5933|biu/cache_ctrl_logic/reg6_b21  (
    .a({\biu/bus_unit/mmu/i [0],open_n36858}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [21]}),
    .c({\biu/paddress [21],\biu/cache_ctrl_logic/pa_temp [21]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [19],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5933_o,open_n36876}),
    .q({open_n36880,\biu/cache_ctrl_logic/pa_temp [21]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUTF1("(B*~(D*~C*A))"),
    //.LUTG0("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    //.LUTG1("(B*~(D*~C*A))"),
    .INIT_LUTF0(16'b0010000000100011),
    .INIT_LUTF1(16'b1100010011001100),
    .INIT_LUTG0(16'b0010000000100011),
    .INIT_LUTG1(16'b1100010011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5934|_al_u5935  (
    .a({\biu/maddress [21],_al_u5934_o}),
    .b({_al_u5933_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [21]}),
    .f({_al_u5934_o,_al_u5935_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5936|biu/bus_unit/mmu/reg1_b21  (
    .a({\biu/maddress [21],open_n36905}),
    .b({_al_u2914_o,open_n36906}),
    .c({_al_u2698_o,_al_u5936_o}),
    .clk(clk_pad),
    .d({\biu/paddress [21],_al_u5935_o}),
    .sr(rst_pad),
    .f({_al_u5936_o,open_n36924}),
    .q({open_n36928,\biu/paddress [21]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000001010011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5938|biu/bus_unit/mmu/reg1_b20  (
    .a({open_n36929,_al_u5938_o}),
    .b({_al_u2914_o,_al_u5941_o}),
    .c({\biu/paddress [20],_al_u2698_o}),
    .clk(clk_pad),
    .d({\biu/maddress [20],_al_u5942_o}),
    .sr(rst_pad),
    .f({_al_u5938_o,open_n36943}),
    .q({open_n36947,\biu/paddress [20]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0110111001111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0110111001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5939|biu/cache_ctrl_logic/reg6_b20  (
    .a({\biu/bus_unit/mmu/i [0],open_n36948}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [20]}),
    .c({\biu/paddress [20],\biu/cache_ctrl_logic/pa_temp [20]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [18],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5939_o,open_n36966}),
    .q({open_n36970,\biu/cache_ctrl_logic/pa_temp [20]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(A*(D@C)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~(A*(D@C)))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100010001001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100010001001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5940|_al_u5941  (
    .a({open_n36971,\biu/maddress [20]}),
    .b({open_n36972,_al_u5940_o}),
    .c({_al_u5939_o,\biu/bus_unit/mmu/i [0]}),
    .d({_al_u2915_o,\biu/bus_unit/mmu/i [1]}),
    .f({_al_u5940_o,_al_u5941_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5942|_al_u5990  (
    .c({\biu/paddress [20],\biu/paddress [12]}),
    .d({_al_u2915_o,_al_u2915_o}),
    .f({_al_u5942_o,_al_u5990_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0101000001010011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5944|biu/bus_unit/mmu/reg1_b19  (
    .a({open_n37025,_al_u5944_o}),
    .b({_al_u2914_o,_al_u5947_o}),
    .c({\biu/paddress [19],_al_u2698_o}),
    .clk(clk_pad),
    .d({\biu/maddress [19],_al_u5948_o}),
    .sr(rst_pad),
    .f({_al_u5944_o,open_n37043}),
    .q({open_n37047,\biu/paddress [19]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0110111001111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5945|biu/cache_ctrl_logic/reg6_b19  (
    .a({\biu/bus_unit/mmu/i [0],open_n37048}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [19]}),
    .c({\biu/paddress [19],\biu/cache_ctrl_logic/pa_temp [19]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [17],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5945_o,open_n37062}),
    .q({open_n37066,\biu/cache_ctrl_logic/pa_temp [19]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*(D@C)))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100010001001100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5946|_al_u5947  (
    .a({open_n37067,\biu/maddress [19]}),
    .b({open_n37068,_al_u5946_o}),
    .c({_al_u5945_o,\biu/bus_unit/mmu/i [0]}),
    .d({_al_u2915_o,\biu/bus_unit/mmu/i [1]}),
    .f({_al_u5946_o,_al_u5947_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u5948|_al_u5978  (
    .c({\biu/paddress [19],\biu/paddress [14]}),
    .d({_al_u2915_o,_al_u2915_o}),
    .f({_al_u5948_o,_al_u5978_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0101000001010011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5950|biu/bus_unit/mmu/reg1_b18  (
    .a({open_n37113,_al_u5950_o}),
    .b({_al_u2914_o,_al_u5953_o}),
    .c({\biu/paddress [18],_al_u2698_o}),
    .clk(clk_pad),
    .d({\biu/maddress [18],_al_u5954_o}),
    .sr(rst_pad),
    .f({_al_u5950_o,open_n37131}),
    .q({open_n37135,\biu/paddress [18]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0110111001111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5951|biu/cache_ctrl_logic/reg6_b18  (
    .a({\biu/bus_unit/mmu/i [0],open_n37136}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [18]}),
    .c({\biu/paddress [18],\biu/cache_ctrl_logic/pa_temp [18]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [16],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5951_o,open_n37150}),
    .q({open_n37154,\biu/cache_ctrl_logic/pa_temp [18]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*(D@C)))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100010001001100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5952|_al_u5953  (
    .a({open_n37155,\biu/maddress [18]}),
    .b({open_n37156,_al_u5952_o}),
    .c({_al_u5951_o,\biu/bus_unit/mmu/i [0]}),
    .d({_al_u2915_o,\biu/bus_unit/mmu/i [1]}),
    .f({_al_u5952_o,_al_u5953_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u5954|_al_u5966  (
    .c({\biu/paddress [18],\biu/paddress [16]}),
    .d({_al_u2915_o,_al_u2915_o}),
    .f({_al_u5954_o,_al_u5966_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000001010011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5956|biu/bus_unit/mmu/reg1_b17  (
    .a({open_n37201,_al_u5956_o}),
    .b({_al_u2914_o,_al_u5959_o}),
    .c({\biu/paddress [17],_al_u2698_o}),
    .clk(clk_pad),
    .d({\biu/maddress [17],_al_u5960_o}),
    .sr(rst_pad),
    .f({_al_u5956_o,open_n37215}),
    .q({open_n37219,\biu/paddress [17]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0110111001111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0110111001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5957|biu/cache_ctrl_logic/reg6_b17  (
    .a({\biu/bus_unit/mmu/i [0],open_n37220}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [17]}),
    .c({\biu/paddress [17],\biu/cache_ctrl_logic/pa_temp [17]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [15],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5957_o,open_n37238}),
    .q({open_n37242,\biu/cache_ctrl_logic/pa_temp [17]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(A*(D@C)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~(A*(D@C)))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100010001001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100010001001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5958|_al_u5959  (
    .a({open_n37243,\biu/maddress [17]}),
    .b({open_n37244,_al_u5958_o}),
    .c({_al_u5957_o,\biu/bus_unit/mmu/i [0]}),
    .d({_al_u2915_o,\biu/bus_unit/mmu/i [1]}),
    .f({_al_u5958_o,_al_u5959_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUT1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000001010011),
    .INIT_LUT1(16'b0000110000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5962|biu/bus_unit/mmu/reg1_b16  (
    .a({open_n37269,_al_u5962_o}),
    .b({_al_u2914_o,_al_u5965_o}),
    .c({\biu/paddress [16],_al_u2698_o}),
    .clk(clk_pad),
    .d({\biu/maddress [16],_al_u5966_o}),
    .sr(rst_pad),
    .f({_al_u5962_o,open_n37283}),
    .q({open_n37287,\biu/paddress [16]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0110111001111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0110111001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5963|biu/cache_ctrl_logic/reg6_b16  (
    .a({\biu/bus_unit/mmu/i [0],open_n37288}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [16]}),
    .c({\biu/paddress [16],\biu/cache_ctrl_logic/pa_temp [16]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [14],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5963_o,open_n37306}),
    .q({open_n37310,\biu/cache_ctrl_logic/pa_temp [16]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(A*(D@C)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~(A*(D@C)))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1100010001001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1100010001001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5964|_al_u5965  (
    .a({open_n37311,\biu/maddress [16]}),
    .b({open_n37312,_al_u5964_o}),
    .c({_al_u5963_o,\biu/bus_unit/mmu/i [0]}),
    .d({_al_u2915_o,\biu/bus_unit/mmu/i [1]}),
    .f({_al_u5964_o,_al_u5965_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0110111001111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5968|biu/cache_ctrl_logic/reg6_b15  (
    .a({\biu/bus_unit/mmu/i [0],open_n37337}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [15]}),
    .c({\biu/paddress [15],\biu/cache_ctrl_logic/pa_temp [15]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [13],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5968_o,open_n37351}),
    .q({open_n37355,\biu/cache_ctrl_logic/pa_temp [15]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5969|_al_u5960  (
    .c({_al_u5968_o,\biu/paddress [17]}),
    .d({_al_u2915_o,_al_u2915_o}),
    .f({_al_u5969_o,_al_u5960_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~A*~(~D*~C)))"),
    //.LUT1("(B*~(A*(D@C)))"),
    .INIT_LUT0(16'b0010001000100011),
    .INIT_LUT1(16'b1100010001001100),
    .MODE("LOGIC"))
    \_al_u5970|_al_u5971  (
    .a({\biu/maddress [15],_al_u5970_o}),
    .b({_al_u5969_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [15]}),
    .f({_al_u5970_o,_al_u5971_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001000011010000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5972|biu/bus_unit/mmu/reg1_b15  (
    .a({\biu/maddress [15],open_n37404}),
    .b({_al_u2914_o,open_n37405}),
    .c({_al_u2698_o,_al_u5972_o}),
    .clk(clk_pad),
    .d({\biu/paddress [15],_al_u5971_o}),
    .sr(rst_pad),
    .f({_al_u5972_o,open_n37423}),
    .q({open_n37427,\biu/paddress [15]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0101000001010011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5974|biu/bus_unit/mmu/reg1_b14  (
    .a({open_n37428,_al_u5974_o}),
    .b({_al_u2914_o,_al_u5977_o}),
    .c({\biu/paddress [14],_al_u2698_o}),
    .clk(clk_pad),
    .d({\biu/maddress [14],_al_u5978_o}),
    .sr(rst_pad),
    .f({_al_u5974_o,open_n37446}),
    .q({open_n37450,\biu/paddress [14]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b0110111001111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5975|biu/cache_ctrl_logic/reg6_b14  (
    .a({\biu/bus_unit/mmu/i [0],open_n37451}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [14]}),
    .c({\biu/paddress [14],\biu/cache_ctrl_logic/pa_temp [14]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [12],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5975_o,open_n37465}),
    .q({open_n37469,\biu/cache_ctrl_logic/pa_temp [14]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*(D@C)))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100010001001100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5976|_al_u5977  (
    .a({open_n37470,\biu/maddress [14]}),
    .b({open_n37471,_al_u5976_o}),
    .c({_al_u5975_o,\biu/bus_unit/mmu/i [0]}),
    .d({_al_u2915_o,\biu/bus_unit/mmu/i [1]}),
    .f({_al_u5976_o,_al_u5977_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0110111001111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0110111001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5980|biu/cache_ctrl_logic/reg6_b13  (
    .a({\biu/bus_unit/mmu/i [0],open_n37492}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [13]}),
    .c({\biu/paddress [13],\biu/cache_ctrl_logic/pa_temp [13]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [11],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5980_o,open_n37510}),
    .q({open_n37514,\biu/cache_ctrl_logic/pa_temp [13]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~A*~(~D*~C)))"),
    //.LUT1("(B*~(A*(D@C)))"),
    .INIT_LUT0(16'b0010001000100011),
    .INIT_LUT1(16'b1100010001001100),
    .MODE("LOGIC"))
    \_al_u5982|_al_u5983  (
    .a({\biu/maddress [13],_al_u5982_o}),
    .b({_al_u5981_o,_al_u2698_o}),
    .c({\biu/bus_unit/mmu/i [0],_al_u2915_o}),
    .d({\biu/bus_unit/mmu/i [1],\biu/paddress [13]}),
    .f({_al_u5982_o,_al_u5983_o}));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001000011010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5984|biu/bus_unit/mmu/reg1_b13  (
    .a({\biu/maddress [13],open_n37535}),
    .b({_al_u2914_o,open_n37536}),
    .c({_al_u2698_o,_al_u5984_o}),
    .clk(clk_pad),
    .d({\biu/paddress [13],_al_u5983_o}),
    .sr(rst_pad),
    .f({_al_u5984_o,open_n37550}),
    .q({open_n37554,\biu/paddress [13]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010011),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0101000001010011),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5986|biu/bus_unit/mmu/reg1_b12  (
    .a({open_n37555,_al_u5986_o}),
    .b({_al_u2914_o,_al_u5989_o}),
    .c({\biu/paddress [12],_al_u2698_o}),
    .clk(clk_pad),
    .d({\biu/maddress [12],_al_u5990_o}),
    .sr(rst_pad),
    .f({_al_u5986_o,open_n37573}),
    .q({open_n37577,\biu/paddress [12]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b0110111001111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b0110111001111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5987|biu/cache_ctrl_logic/reg6_b12  (
    .a({\biu/bus_unit/mmu/i [0],open_n37578}),
    .b({\biu/bus_unit/mmu/i [1],\biu/paddress [12]}),
    .c({\biu/paddress [12],\biu/cache_ctrl_logic/pa_temp [12]}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [10],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u5987_o,open_n37596}),
    .q({open_n37600,\biu/cache_ctrl_logic/pa_temp [12]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*(D@C)))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100010001001100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u5988|_al_u5989  (
    .a({open_n37601,\biu/maddress [12]}),
    .b({open_n37602,_al_u5988_o}),
    .c({_al_u5987_o,\biu/bus_unit/mmu/i [0]}),
    .d({_al_u2915_o,\biu/bus_unit/mmu/i [1]}),
    .f({_al_u5988_o,_al_u5989_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u5994|_al_u5109  (
    .c({_al_u5108_o,wb_valid}),
    .d({_al_u5157_o,_al_u5108_o}),
    .f({\cu_ru/m_s_status/u14_sel_is_2_o ,\cu_ru/trap_target_m }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000001001100),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b0100000001001100),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5995|cu_ru/m_s_tvec/reg0_b9  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[9]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [9],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [9],id_ins_pc[9]}),
    .mi({open_n37654,csr_data[9]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [9],_al_u7891_o}),
    .q({open_n37669,\cu_ru/stvec [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000001001100),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5996|cu_ru/m_s_tvec/reg0_b8  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[8]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [8],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [8],id_ins_pc[8]}),
    .mi({open_n37680,csr_data[8]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [8],_al_u7871_o}),
    .q({open_n37684,\cu_ru/stvec [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000001001100),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u5997|cu_ru/m_s_tvec/reg0_b7  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[7]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [7],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [7],id_ins_pc[7]}),
    .mi({open_n37695,csr_data[7]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [7],_al_u7836_o}),
    .q({open_n37699,\cu_ru/stvec [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6000|cu_ru/m_cycle_event/reg0_b61  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6763_o}),
    .b({\cu_ru/trap_target_m ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/stvec [61],\cu_ru/minstret [61]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [61],\cu_ru/stvec [61]}),
    .mi({open_n37710,\cu_ru/m_cycle_event/n4 [61]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [61],_al_u6974_o}),
    .q({open_n37714,\cu_ru/minstret [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000001001100),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b0100000001001100),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6002|cu_ru/m_s_tvec/reg0_b6  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[6]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [6],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [6],id_ins_pc[6]}),
    .mi({open_n37718,csr_data[6]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [6],_al_u7814_o}),
    .q({open_n37733,\cu_ru/stvec [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6003|cu_ru/m_s_tvec/reg1_b59  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6785_o}),
    .b({\cu_ru/trap_target_m ,_al_u6790_o}),
    .c({\cu_ru/stvec [59],\cu_ru/read_mtvec_sel_lutinv }),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [59],\cu_ru/mtvec [59]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [59],csr_data[59]}),
    .q({open_n37753,\cu_ru/mtvec [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6007|cu_ru/m_s_tvec/reg1_b55  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6828_o}),
    .b({\cu_ru/trap_target_m ,_al_u6829_o}),
    .c({\cu_ru/stvec [55],\cu_ru/read_mtvec_sel_lutinv }),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [55],\cu_ru/mtvec [55]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [55],csr_data[55]}),
    .q({open_n37773,\cu_ru/mtvec [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6008|cu_ru/m_cycle_event/reg0_b54  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6763_o}),
    .b({\cu_ru/trap_target_m ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/stvec [54],\cu_ru/minstret [54]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [54],\cu_ru/stvec [54]}),
    .mi({open_n37777,\cu_ru/m_cycle_event/n4 [54]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [54],_al_u6838_o}),
    .q({open_n37792,\cu_ru/minstret [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6010|cu_ru/m_cycle_event/reg0_b52  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6763_o}),
    .b({\cu_ru/trap_target_m ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/stvec [52],\cu_ru/minstret [52]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [52],\cu_ru/stvec [52]}),
    .mi({open_n37803,\cu_ru/m_cycle_event/n4 [52]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [52],_al_u6857_o}),
    .q({open_n37807,\cu_ru/minstret [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6011|cu_ru/m_cycle_event/reg0_b51  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6763_o}),
    .b({\cu_ru/trap_target_m ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/stvec [51],\cu_ru/minstret [51]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [51],\cu_ru/stvec [51]}),
    .mi({open_n37818,\cu_ru/m_cycle_event/n4 [51]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [51],_al_u6867_o}),
    .q({open_n37822,\cu_ru/minstret [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000001001100),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6013|cu_ru/m_s_tvec/reg0_b5  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[5]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [5],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [5],id_ins_pc[5]}),
    .mi({open_n37833,csr_data[5]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [5],_al_u7895_o}),
    .q({open_n37837,\cu_ru/stvec [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*A*~(D*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011101110111),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6015|cu_ru/m_s_tvec/reg1_b48  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6896_o}),
    .b({\cu_ru/trap_target_m ,_al_u6897_o}),
    .c({\cu_ru/stvec [48],\cu_ru/read_mtvec_sel_lutinv }),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [48],\cu_ru/mtvec [48]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [48],csr_data[48]}),
    .q({open_n37853,\cu_ru/mtvec [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6017|cu_ru/m_cycle_event/reg0_b46  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6763_o}),
    .b({\cu_ru/trap_target_m ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/stvec [46],\cu_ru/minstret [46]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [46],\cu_ru/stvec [46]}),
    .mi({open_n37857,\cu_ru/m_cycle_event/n4 [46]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [46],_al_u6910_o}),
    .q({open_n37872,\cu_ru/minstret [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6021|cu_ru/m_s_tvec/reg0_b42  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[42]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [42],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [42],id_ins_pc[42]}),
    .mi({open_n37883,csr_data[42]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [42],_al_u7530_o}),
    .q({open_n37887,\cu_ru/stvec [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000001001100),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6024|cu_ru/m_s_tvec/reg0_b4  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[4]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [4],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [4],id_ins_pc[4]}),
    .mi({open_n37898,csr_data[4]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [4],_al_u7838_o}),
    .q({open_n37902,\cu_ru/stvec [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6028|cu_ru/m_cycle_event/reg0_b36  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6763_o}),
    .b({\cu_ru/trap_target_m ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/stvec [36],\cu_ru/minstret [36]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [36],\cu_ru/stvec [36]}),
    .mi({open_n37913,\cu_ru/m_cycle_event/n4 [36]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [36],_al_u7065_o}),
    .q({open_n37917,\cu_ru/minstret [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6029|cu_ru/m_cycle_event/reg0_b35  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6763_o}),
    .b({\cu_ru/trap_target_m ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/stvec [35],\cu_ru/minstret [35]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [35],\cu_ru/stvec [35]}),
    .mi({open_n37921,\cu_ru/m_cycle_event/n4 [35]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [35],_al_u7223_o}),
    .q({open_n37936,\cu_ru/minstret [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6031|cu_ru/m_s_tvec/reg0_b33  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[33]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [33],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [33],id_ins_pc[33]}),
    .mi({open_n37940,csr_data[33]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [33],_al_u7816_o}),
    .q({open_n37955,\cu_ru/stvec [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6032|cu_ru/m_s_tvec/reg0_b32  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[32]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [32],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [32],id_ins_pc[32]}),
    .mi({open_n37966,csr_data[32]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [32],_al_u7819_o}),
    .q({open_n37970,\cu_ru/stvec [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6034|cu_ru/m_s_tvec/reg0_b30  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[30]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [30],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [30],id_ins_pc[30]}),
    .mi({open_n37981,csr_data[30]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [30],_al_u7822_o}),
    .q({open_n37985,\cu_ru/stvec [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6035|cu_ru/m_s_tvec/reg0_b29  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[29]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [29],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [29],id_ins_pc[29]}),
    .mi({open_n37989,csr_data[29]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [29],_al_u7585_o}),
    .q({open_n38004,\cu_ru/stvec [29]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6036|cu_ru/m_s_tvec/reg0_b28  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[28]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [28],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [28],id_ins_pc[28]}),
    .mi({open_n38015,csr_data[28]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [28],_al_u7825_o}),
    .q({open_n38019,\cu_ru/stvec [28]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6037|cu_ru/m_s_tvec/reg0_b27  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[27]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [27],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [27],id_ins_pc[27]}),
    .mi({open_n38030,csr_data[27]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [27],_al_u7588_o}),
    .q({open_n38034,\cu_ru/stvec [27]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6038|cu_ru/m_s_tvec/reg0_b26  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[26]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [26],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [26],id_ins_pc[26]}),
    .mi({open_n38038,csr_data[26]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [26],_al_u7591_o}),
    .q({open_n38053,\cu_ru/stvec [26]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6039|cu_ru/m_s_tvec/reg0_b25  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[25]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [25],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [25],id_ins_pc[25]}),
    .mi({open_n38057,csr_data[25]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [25],_al_u7685_o}),
    .q({open_n38072,\cu_ru/stvec [25]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6040|cu_ru/m_s_tvec/reg0_b24  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[24]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [24],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [24],id_ins_pc[24]}),
    .mi({open_n38083,csr_data[24]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [24],_al_u7594_o}),
    .q({open_n38087,\cu_ru/stvec [24]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6041|cu_ru/m_s_tvec/reg0_b23  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[23]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [23],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [23],id_ins_pc[23]}),
    .mi({open_n38098,csr_data[23]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [23],_al_u7597_o}),
    .q({open_n38102,\cu_ru/stvec [23]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6042|cu_ru/m_s_tvec/reg0_b22  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[22]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [22],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [22],id_ins_pc[22]}),
    .mi({open_n38106,csr_data[22]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [22],_al_u7842_o}),
    .q({open_n38121,\cu_ru/stvec [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6043|cu_ru/m_s_tvec/reg0_b21  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[21]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [21],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [21],id_ins_pc[21]}),
    .mi({open_n38125,csr_data[21]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [21],_al_u7689_o}),
    .q({open_n38140,\cu_ru/stvec [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6044|cu_ru/m_s_tvec/reg0_b20  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[20]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [20],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [20],id_ins_pc[20]}),
    .mi({open_n38151,csr_data[20]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [20],_al_u7845_o}),
    .q({open_n38155,\cu_ru/stvec [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6045|cu_ru/m_s_tvec/reg0_b19  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[19]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [19],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [19],id_ins_pc[19]}),
    .mi({open_n38166,csr_data[19]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [19],_al_u7828_o}),
    .q({open_n38170,\cu_ru/stvec [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6046|cu_ru/m_s_tvec/reg0_b18  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[18]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [18],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [18],id_ins_pc[18]}),
    .mi({open_n38174,csr_data[18]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [18],_al_u7848_o}),
    .q({open_n38189,\cu_ru/stvec [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6047|cu_ru/m_s_tvec/reg0_b17  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[17]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [17],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [17],id_ins_pc[17]}),
    .mi({open_n38193,csr_data[17]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [17],_al_u7851_o}),
    .q({open_n38208,\cu_ru/stvec [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6048|cu_ru/m_s_tvec/reg0_b16  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[16]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [16],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [16],id_ins_pc[16]}),
    .mi({open_n38219,csr_data[16]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [16],_al_u7649_o}),
    .q({open_n38223,\cu_ru/stvec [16]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6049|cu_ru/m_s_tvec/reg0_b15  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[15]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [15],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [15],id_ins_pc[15]}),
    .mi({open_n38234,csr_data[15]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [15],_al_u7705_o}),
    .q({open_n38238,\cu_ru/stvec [15]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6050|cu_ru/m_s_tvec/reg0_b14  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[14]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [14],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [14],id_ins_pc[14]}),
    .mi({open_n38242,csr_data[14]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [14],_al_u7831_o}),
    .q({open_n38257,\cu_ru/stvec [14]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("~(~(D*B)*~(C*A))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b1110110010100000),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b1110110010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6051|cu_ru/m_s_tvec/reg0_b13  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[13]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [13],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [13],id_ins_pc[13]}),
    .mi({open_n38261,csr_data[13]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [13],_al_u7707_o}),
    .q({open_n38276,\cu_ru/stvec [13]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6052|cu_ru/m_s_tvec/reg0_b12  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[12]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [12],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [12],id_ins_pc[12]}),
    .mi({open_n38287,csr_data[12]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [12],_al_u7854_o}),
    .q({open_n38291,\cu_ru/stvec [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("~(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000001001100),
    .INIT_LUT1(16'b1110110010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6053|cu_ru/m_s_tvec/reg0_b11  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,csr_data[11]}),
    .b({\cu_ru/trap_target_m ,_al_u7141_o}),
    .c({\cu_ru/stvec [11],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [11],id_ins_pc[11]}),
    .mi({open_n38302,csr_data[11]}),
    .sr(rst_pad),
    .f({\cu_ru/tvec [11],_al_u7834_o}),
    .q({open_n38306,\cu_ru/stvec [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/ID/ins_dec.v(674)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(C*~B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100111111111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6058|ins_dec/unsign_reg  (
    .b({id_ins[31],_al_u6058_o}),
    .c({id_ins[30],_al_u6061_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3939_o,_al_u4806_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6058_o,open_n38325}),
    .q({open_n38329,unsign}));  // ../../RTL/CPU/ID/ins_dec.v(674)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*C*B))"),
    //.LUT1("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT_LUT0(16'b0010101010101010),
    .INIT_LUT1(16'b1100010010000000),
    .MODE("LOGIC"))
    \_al_u6060|_al_u6059  (
    .a({_al_u4064_o,\ins_dec/op_load }),
    .b({_al_u3216_o,_al_u3216_o}),
    .c({_al_u3217_o,_al_u3217_o}),
    .d({_al_u6059_o,_al_u3384_o}),
    .f({\ins_dec/n198_lutinv ,_al_u6059_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6061|_al_u4801  (
    .a({open_n38350,_al_u3925_o}),
    .b({\ins_dec/funct7_32_lutinv ,_al_u3216_o}),
    .c({_al_u4801_o,_al_u3217_o}),
    .d({\ins_dec/n198_lutinv ,_al_u3384_o}),
    .f({_al_u6061_o,_al_u4801_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6063|ins_dec/reg7_b55  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[55]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[55],rs1_data[55]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6063_o,open_n38389}),
    .q({open_n38393,as1[55]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6064|ins_dec/reg6_b55  (
    .a({_al_u5144_o,open_n38394}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_055 ,_al_u6064_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_055 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6063_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6064_o,open_n38411}),
    .q({open_n38415,ds2[55]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6067|ins_dec/reg7_b54  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[54]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[54],rs1_data[54]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6067_o,open_n38434}),
    .q({open_n38438,as1[54]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6068|ins_dec/reg6_b54  (
    .a({_al_u5144_o,open_n38439}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_054 ,_al_u6068_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_054 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6067_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6068_o,open_n38452}),
    .q({open_n38456,ds2[54]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6070|ins_dec/reg7_b53  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[53]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[53],rs1_data[53]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6070_o,open_n38475}),
    .q({open_n38479,as1[53]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6071|ins_dec/reg6_b53  (
    .a({_al_u5144_o,open_n38480}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_053 ,_al_u6071_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_053 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6070_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6071_o,open_n38493}),
    .q({open_n38497,ds2[53]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6073|ins_dec/reg7_b52  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[52]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[52],rs1_data[52]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6073_o,open_n38512}),
    .q({open_n38516,as1[52]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6074|ins_dec/reg6_b52  (
    .a({_al_u5144_o,open_n38517}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_052 ,_al_u6074_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_052 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6073_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6074_o,open_n38534}),
    .q({open_n38538,ds2[52]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6076|ins_dec/reg7_b51  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[51]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[51],rs1_data[51]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6076_o,open_n38553}),
    .q({open_n38557,as1[51]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6077|ins_dec/reg6_b51  (
    .a({_al_u5144_o,open_n38558}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_051 ,_al_u6077_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_051 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6076_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6077_o,open_n38575}),
    .q({open_n38579,ds2[51]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6079|ins_dec/reg7_b50  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[50]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[50],rs1_data[50]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6079_o,open_n38598}),
    .q({open_n38602,as1[50]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6080|ins_dec/reg6_b50  (
    .a({_al_u5144_o,open_n38603}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_050 ,_al_u6080_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_050 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6079_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6080_o,open_n38616}),
    .q({open_n38620,ds2[50]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6082|ins_dec/reg7_b49  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[49]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[49],rs1_data[49]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6082_o,open_n38635}),
    .q({open_n38639,as1[49]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6083|ins_dec/reg6_b49  (
    .a({_al_u5144_o,open_n38640}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_049 ,_al_u6083_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_049 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6082_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6083_o,open_n38653}),
    .q({open_n38657,ds2[49]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6085|ins_dec/reg7_b48  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[48]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[48],rs1_data[48]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6085_o,open_n38672}),
    .q({open_n38676,as1[48]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6086|ins_dec/reg6_b48  (
    .a({_al_u5144_o,open_n38677}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_048 ,_al_u6086_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_048 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6085_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6086_o,open_n38694}),
    .q({open_n38698,ds2[48]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6088|ins_dec/reg7_b47  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[47]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[47],rs1_data[47]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6088_o,open_n38717}),
    .q({open_n38721,as1[47]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6089|ins_dec/reg6_b47  (
    .a({_al_u5144_o,open_n38722}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_047 ,_al_u6089_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_047 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6088_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6089_o,open_n38739}),
    .q({open_n38743,ds2[47]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6091|ins_dec/reg7_b46  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[46]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[46],rs1_data[46]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6091_o,open_n38762}),
    .q({open_n38766,as1[46]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6092|ins_dec/reg6_b46  (
    .a({_al_u5144_o,open_n38767}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_046 ,_al_u6092_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_046 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6091_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6092_o,open_n38780}),
    .q({open_n38784,ds2[46]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6094|ins_dec/reg7_b45  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[45]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[45],rs1_data[45]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6094_o,open_n38799}),
    .q({open_n38803,as1[45]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6095|ins_dec/reg6_b45  (
    .a({_al_u5144_o,open_n38804}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_045 ,_al_u6095_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_045 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6094_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6095_o,open_n38817}),
    .q({open_n38821,ds2[45]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6097|ins_dec/reg7_b44  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[44]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[44],rs1_data[44]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6097_o,open_n38836}),
    .q({open_n38840,as1[44]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6098|ins_dec/reg6_b44  (
    .a({_al_u5144_o,open_n38841}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_044 ,_al_u6098_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_044 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6097_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6098_o,open_n38858}),
    .q({open_n38862,ds2[44]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6101|ins_dec/reg6_b43  (
    .a({_al_u5144_o,open_n38863}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_043 ,_al_u6101_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_043 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6100_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6101_o,open_n38880}),
    .q({open_n38884,ds2[43]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6103|ins_dec/reg7_b42  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[42]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[42],rs1_data[42]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6103_o,open_n38903}),
    .q({open_n38907,as1[42]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6104|ins_dec/reg6_b42  (
    .a({_al_u5144_o,open_n38908}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_042 ,_al_u6104_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_042 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6103_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6104_o,open_n38921}),
    .q({open_n38925,ds2[42]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6106|_al_u4929  (
    .a({open_n38926,\cu_ru/n45_lutinv }),
    .b({_al_u5858_o,\cu_ru/al_ram_gpr_do_i0_041 }),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,\cu_ru/al_ram_gpr_do_i1_041 }),
    .d({rs1_data[41],\cu_ru/n46 [4]}),
    .f({_al_u6106_o,rs1_data[41]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6107|ins_dec/reg6_b41  (
    .a({_al_u5144_o,open_n38951}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_041 ,_al_u6107_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_041 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6106_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6107_o,open_n38964}),
    .q({open_n38968,ds2[41]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6109|_al_u4931  (
    .a({open_n38969,\cu_ru/n45_lutinv }),
    .b({_al_u5858_o,\cu_ru/al_ram_gpr_do_i0_040 }),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,\cu_ru/al_ram_gpr_do_i1_040 }),
    .d({rs1_data[40],\cu_ru/n46 [4]}),
    .f({_al_u6109_o,rs1_data[40]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6110|ins_dec/reg6_b40  (
    .a({_al_u5144_o,open_n38994}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_040 ,_al_u6110_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_040 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6109_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6110_o,open_n39011}),
    .q({open_n39015,ds2[40]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001110100111111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001110100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6113|ins_dec/reg10_b11  (
    .a({_al_u6112_o,open_n39016}),
    .b({_al_u3927_o,open_n39017}),
    .c({id_ins[24],id_ins[11]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[11],id_ill_ins}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6113_o,open_n39034}),
    .q({open_n39038,ex_exc_code[11]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A*~(~C*~B))"),
    //.LUT1("(C*~(B*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010100),
    .INIT_LUT1(16'b0011000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6114|ins_dec/reg5_b4  (
    .a({open_n39039,_al_u7838_o}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,rs1_data[4]}),
    .c({_al_u6113_o,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[4],\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u6114_o,open_n39052}),
    .q({open_n39056,ds1[4]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u6116|_al_u4935  (
    .a({open_n39057,\cu_ru/n45_lutinv }),
    .b({_al_u5858_o,\cu_ru/al_ram_gpr_do_i0_039 }),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,\cu_ru/al_ram_gpr_do_i1_039 }),
    .d({rs1_data[39],\cu_ru/n46 [4]}),
    .f({_al_u6116_o,rs1_data[39]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6117|ins_dec/reg6_b39  (
    .a({_al_u5144_o,open_n39078}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_039 ,_al_u6117_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_039 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6116_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6117_o,open_n39095}),
    .q({open_n39099,ds2[39]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u6119|_al_u4937  (
    .a({open_n39100,\cu_ru/n45_lutinv }),
    .b({_al_u5858_o,\cu_ru/al_ram_gpr_do_i0_038 }),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,\cu_ru/al_ram_gpr_do_i1_038 }),
    .d({rs1_data[38],\cu_ru/n46 [4]}),
    .f({_al_u6119_o,rs1_data[38]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6120|ins_dec/reg6_b38  (
    .a({_al_u5144_o,open_n39121}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_038 ,_al_u6120_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_038 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6119_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6120_o,open_n39134}),
    .q({open_n39138,ds2[38]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6122|_al_u4939  (
    .a({open_n39139,\cu_ru/n45_lutinv }),
    .b({_al_u5858_o,\cu_ru/al_ram_gpr_do_i0_037 }),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,\cu_ru/al_ram_gpr_do_i1_037 }),
    .d({rs1_data[37],\cu_ru/n46 [4]}),
    .f({_al_u6122_o,rs1_data[37]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6123|ins_dec/reg6_b37  (
    .a({_al_u5144_o,open_n39164}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_037 ,_al_u6123_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_037 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6122_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6123_o,open_n39177}),
    .q({open_n39181,ds2[37]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0101000001000100),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0101000001000100),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6125|_al_u4941  (
    .a({open_n39182,\cu_ru/n45_lutinv }),
    .b({_al_u5858_o,\cu_ru/al_ram_gpr_do_i0_036 }),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,\cu_ru/al_ram_gpr_do_i1_036 }),
    .d({rs1_data[36],\cu_ru/n46 [4]}),
    .f({_al_u6125_o,rs1_data[36]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6126|ins_dec/reg6_b36  (
    .a({_al_u5144_o,open_n39207}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_036 ,_al_u6126_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_036 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6125_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6126_o,open_n39224}),
    .q({open_n39228,ds2[36]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6128|ins_dec/reg7_b35  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[35]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[35],rs1_data[35]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6128_o,open_n39243}),
    .q({open_n39247,as1[35]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6129|ins_dec/reg6_b35  (
    .a({_al_u5144_o,open_n39248}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_035 ,_al_u6129_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_035 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6128_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6129_o,open_n39265}),
    .q({open_n39269,ds2[35]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u6131|_al_u4945  (
    .a({open_n39270,\cu_ru/n45_lutinv }),
    .b({_al_u5858_o,\cu_ru/al_ram_gpr_do_i0_034 }),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,\cu_ru/al_ram_gpr_do_i1_034 }),
    .d({rs1_data[34],\cu_ru/n46 [4]}),
    .f({_al_u6131_o,rs1_data[34]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6132|ins_dec/reg6_b34  (
    .a({_al_u5144_o,open_n39291}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_034 ,_al_u6132_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_034 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6131_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6132_o,open_n39304}),
    .q({open_n39308,ds2[34]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6134|ins_dec/reg7_b33  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[33]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[33],rs1_data[33]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6134_o,open_n39323}),
    .q({open_n39327,as1[33]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6135|ins_dec/reg6_b33  (
    .a({_al_u5144_o,open_n39328}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_033 ,_al_u6135_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_033 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6134_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6135_o,open_n39341}),
    .q({open_n39345,ds2[33]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6137|ins_dec/reg7_b32  (
    .b({_al_u5858_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[32]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[32],rs1_data[32]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6137_o,open_n39364}),
    .q({open_n39368,as1[32]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6138|ins_dec/reg6_b32  (
    .a({_al_u5144_o,open_n39369}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_032 ,_al_u6138_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_032 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6137_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6138_o,open_n39386}),
    .q({open_n39390,ds2[32]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0101000001000100),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u6140|_al_u4951  (
    .a({open_n39391,\cu_ru/n45_lutinv }),
    .b({_al_u5858_o,\cu_ru/al_ram_gpr_do_i0_031 }),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,\cu_ru/al_ram_gpr_do_i1_031 }),
    .d({rs1_data[31],\cu_ru/n46 [4]}),
    .f({_al_u6140_o,rs1_data[31]}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6141|ins_dec/reg6_b31  (
    .a({_al_u5144_o,open_n39412}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_031 ,_al_u6141_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_031 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6140_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6141_o,open_n39429}),
    .q({open_n39433,ds2[31]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0100011101110111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0100011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6143|ins_dec/reg7_b30  (
    .a({rs1_data[30],open_n39434}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[30]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[30],rs1_data[30]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6143_o,open_n39451}),
    .q({open_n39455,as1[30]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6144|ins_dec/reg6_b30  (
    .a({_al_u5144_o,open_n39456}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_030 ,_al_u6144_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_030 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6143_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6144_o,open_n39469}),
    .q({open_n39473,ds2[30]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0001110100111111),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0001110100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6146|ins_dec/reg8_b3  (
    .a({_al_u6112_o,open_n39474}),
    .b({_al_u3927_o,open_n39475}),
    .c({id_ins[23],_al_u4073_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[10],_al_u4072_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6146_o,open_n39492}),
    .q({open_n39496,as2[3]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A*~(~C*~B))"),
    //.LUT1("(C*~(B*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010100),
    .INIT_LUT1(16'b0011000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6147|ins_dec/reg5_b3  (
    .a({open_n39497,_al_u7840_o}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,rs1_data[3]}),
    .c({_al_u6146_o,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[3],\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u6147_o,open_n39510}),
    .q({open_n39514,ds1[3]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0100011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6149|ins_dec/reg7_b29  (
    .a({rs1_data[29],open_n39515}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[29]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[29],rs1_data[29]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6149_o,open_n39528}),
    .q({open_n39532,as1[29]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6150|ins_dec/reg6_b29  (
    .a({_al_u5144_o,open_n39533}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_029 ,_al_u6150_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_029 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6149_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6150_o,open_n39546}),
    .q({open_n39550,ds2[29]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0100011101110111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0100011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6152|ins_dec/reg7_b28  (
    .a({rs1_data[28],open_n39551}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[28]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[28],rs1_data[28]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6152_o,open_n39568}),
    .q({open_n39572,as1[28]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6153|ins_dec/reg6_b28  (
    .a({_al_u5144_o,open_n39573}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_028 ,_al_u6153_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_028 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6152_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6153_o,open_n39590}),
    .q({open_n39594,ds2[28]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0100011101110111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0100011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6155|ins_dec/reg7_b27  (
    .a({rs1_data[27],open_n39595}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[27]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[27],rs1_data[27]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6155_o,open_n39612}),
    .q({open_n39616,as1[27]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6156|ins_dec/reg6_b27  (
    .a({_al_u5144_o,open_n39617}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_027 ,_al_u6156_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_027 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6155_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6156_o,open_n39634}),
    .q({open_n39638,ds2[27]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0100011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6158|ins_dec/reg7_b26  (
    .a({rs1_data[26],open_n39639}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[26]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[26],rs1_data[26]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6158_o,open_n39652}),
    .q({open_n39656,as1[26]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6159|ins_dec/reg6_b26  (
    .a({_al_u5144_o,open_n39657}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_026 ,_al_u6159_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_026 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6158_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6159_o,open_n39670}),
    .q({open_n39674,ds2[26]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0100011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6161|ins_dec/reg7_b25  (
    .a({rs1_data[25],open_n39675}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[25]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[25],rs1_data[25]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6161_o,open_n39688}),
    .q({open_n39692,as1[25]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6162|ins_dec/reg6_b25  (
    .a({_al_u5144_o,open_n39693}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_025 ,_al_u6162_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_025 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6161_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6162_o,open_n39706}),
    .q({open_n39710,ds2[25]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0100011101110111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0100011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6164|ins_dec/reg7_b24  (
    .a({rs1_data[24],open_n39711}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[24]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[24],rs1_data[24]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6164_o,open_n39728}),
    .q({open_n39732,as1[24]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6165|ins_dec/reg6_b24  (
    .a({_al_u5144_o,open_n39733}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_024 ,_al_u6165_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_024 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6164_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6165_o,open_n39750}),
    .q({open_n39754,ds2[24]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0100011101110111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0100011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6167|ins_dec/reg7_b23  (
    .a({rs1_data[23],open_n39755}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[23]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[23],rs1_data[23]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6167_o,open_n39772}),
    .q({open_n39776,as1[23]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6168|ins_dec/reg6_b23  (
    .a({_al_u5144_o,open_n39777}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_023 ,_al_u6168_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_023 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6167_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6168_o,open_n39794}),
    .q({open_n39798,ds2[23]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0100011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6170|ins_dec/reg7_b22  (
    .a({rs1_data[22],open_n39799}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[22]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[22],rs1_data[22]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6170_o,open_n39812}),
    .q({open_n39816,as1[22]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6171|ins_dec/reg6_b22  (
    .a({_al_u5144_o,open_n39817}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_022 ,_al_u6171_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_022 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6170_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6171_o,open_n39830}),
    .q({open_n39834,ds2[22]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0100011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6173|ins_dec/reg7_b21  (
    .a({rs1_data[21],open_n39835}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[21]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[21],rs1_data[21]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6173_o,open_n39848}),
    .q({open_n39852,as1[21]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6174|ins_dec/reg6_b21  (
    .a({_al_u5144_o,open_n39853}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_021 ,_al_u6174_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_021 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6173_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6174_o,open_n39866}),
    .q({open_n39870,ds2[21]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0100011101110111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0100011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6176|ins_dec/reg7_b20  (
    .a({rs1_data[20],open_n39871}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[20]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[20],rs1_data[20]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6176_o,open_n39888}),
    .q({open_n39892,as1[20]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6177|ins_dec/reg6_b20  (
    .a({_al_u5144_o,open_n39893}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_020 ,_al_u6177_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_020 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6176_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6177_o,open_n39910}),
    .q({open_n39914,ds2[20]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~A*~(~C*~B))"),
    //.LUTF1("~(~C*~((~D*A))*~(B)+~C*(~D*A)*~(B)+~(~C)*(~D*A)*B+~C*(~D*A)*B)"),
    //.LUTG0("(~D*~A*~(~C*~B))"),
    //.LUTG1("~(~C*~((~D*A))*~(B)+~C*(~D*A)*~(B)+~(~C)*(~D*A)*B+~C*(~D*A)*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000001010100),
    .INIT_LUTF1(16'b1111110001110100),
    .INIT_LUTG0(16'b0000000001010100),
    .INIT_LUTG1(16'b1111110001110100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6179|ins_dec/reg5_b2  (
    .a({rs1_data[2],_al_u7887_o}),
    .b({\ins_dec/n239 ,rs1_data[2]}),
    .c({_al_u3955_o,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3216_o,\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u6179_o,open_n39931}),
    .q({open_n39935,ds1[2]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A*~(~D*C))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0100010000000100),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u6180|_al_u6181  (
    .a({open_n39936,_al_u6180_o}),
    .b({_al_u6112_o,_al_u4086_o}),
    .c({id_ins[9],_al_u3927_o}),
    .d({_al_u6179_o,id_ins[22]}),
    .f({_al_u6180_o,_al_u6181_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0100011101110111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0100011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6183|ins_dec/reg7_b19  (
    .a({rs1_data[19],open_n39957}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[19]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[19],rs1_data[19]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6183_o,open_n39974}),
    .q({open_n39978,as1[19]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6184|ins_dec/reg6_b19  (
    .a({_al_u5144_o,open_n39979}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_019 ,_al_u6184_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_019 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6183_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6184_o,open_n39996}),
    .q({open_n40000,ds2[19]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0100011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6186|ins_dec/reg7_b18  (
    .a({rs1_data[18],open_n40001}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[18]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[18],rs1_data[18]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6186_o,open_n40014}),
    .q({open_n40018,as1[18]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6187|ins_dec/reg6_b18  (
    .a({_al_u5144_o,open_n40019}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_018 ,_al_u6187_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_018 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6186_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6187_o,open_n40032}),
    .q({open_n40036,ds2[18]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0100011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6189|ins_dec/reg7_b17  (
    .a({rs1_data[17],open_n40037}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[17]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[17],rs1_data[17]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6189_o,open_n40050}),
    .q({open_n40054,as1[17]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6190|ins_dec/reg6_b17  (
    .a({_al_u5144_o,open_n40055}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_017 ,_al_u6190_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_017 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6189_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6190_o,open_n40068}),
    .q({open_n40072,ds2[17]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0100011101110111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0100011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6192|ins_dec/reg7_b16  (
    .a({rs1_data[16],open_n40073}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[16]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[16],rs1_data[16]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6192_o,open_n40090}),
    .q({open_n40094,as1[16]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6193|ins_dec/reg6_b16  (
    .a({_al_u5144_o,open_n40095}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_016 ,_al_u6193_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_016 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6192_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6193_o,open_n40112}),
    .q({open_n40116,ds2[16]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0100011101110111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0100011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6195|ins_dec/reg7_b15  (
    .a({rs1_data[15],open_n40117}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[15]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({id_ins[15],rs1_data[15]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6195_o,open_n40134}),
    .q({open_n40138,as1[15]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6196|ins_dec/reg6_b15  (
    .a({_al_u5144_o,open_n40139}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_015 ,_al_u6196_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_015 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6195_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6196_o,open_n40156}),
    .q({open_n40160,ds2[15]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("~((B*A)*~(C)*~(D)+(B*A)*C*~(D)+~((B*A))*C*D+(B*A)*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0000111101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6198|ins_dec/reg7_b14  (
    .a({rs1_data[14],open_n40161}),
    .b({\ins_dec/n239 ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[14]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3216_o,rs1_data[14]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6198_o,open_n40174}),
    .q({open_n40178,as1[14]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6199|ins_dec/reg6_b14  (
    .a({_al_u5144_o,open_n40179}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_014 ,_al_u6199_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_014 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6198_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6199_o,open_n40192}),
    .q({open_n40196,ds2[14]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0100011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6201|ins_dec/reg7_b13  (
    .a({rs1_data[13],open_n40197}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[13]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3217_o,rs1_data[13]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6201_o,open_n40210}),
    .q({open_n40214,as1[13]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~B*D)"),
    //.LUT1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011111111),
    .INIT_LUT1(16'b1010000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6202|ins_dec/reg6_b13  (
    .a({_al_u5144_o,open_n40215}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_013 ,_al_u6202_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_013 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6201_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6202_o,open_n40228}),
    .q({open_n40232,ds2[13]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0100011101110111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0100011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6204|ins_dec/reg7_b12  (
    .a({rs1_data[12],open_n40233}),
    .b({\ins_dec/mux19_b10_sel_is_2_o ,_al_u4875_o}),
    .c({_al_u3955_o,id_ins_pc[12]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3384_o,rs1_data[12]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6204_o,open_n40250}),
    .q({open_n40254,as1[12]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*D)"),
    //.LUTF1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG0("~(~C*~B*D)"),
    //.LUTG1("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110011111111),
    .INIT_LUTF1(16'b1010000010001000),
    .INIT_LUTG0(16'b1111110011111111),
    .INIT_LUTG1(16'b1010000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6205|ins_dec/reg6_b12  (
    .a({_al_u5144_o,open_n40255}),
    .b({\cu_ru/al_ram_gpr_al_u0_do_i0_012 ,_al_u6205_o}),
    .c({\cu_ru/al_ram_gpr_al_u0_do_i1_012 ,_al_u6065_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\cu_ru/n49 [4],_al_u6204_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6205_o,open_n40272}),
    .q({open_n40276,ds2[12]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6208|_al_u5865  (
    .b({_al_u6207_o,_al_u5858_o}),
    .c({id_ins[8],\ins_dec/mux19_b10_sel_is_2_o }),
    .d({_al_u6112_o,rs1_data[61]}),
    .f({_al_u6208_o,_al_u5865_o}));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~A*~(~C*~B))"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(~D*~A*~(~C*~B))"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000001010100),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000000001010100),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6209|ins_dec/reg5_b1  (
    .a({open_n40303,_al_u7893_o}),
    .b({_al_u6208_o,rs1_data[1]}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,_al_u7141_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[1],\ins_dec/op_lui_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({_al_u6209_o,open_n40320}),
    .q({open_n40324,ds1[1]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u6212|_al_u9203  (
    .b({_al_u6211_o,open_n40327}),
    .c({id_ins[7],\ins_dec/n107 }),
    .d({_al_u6112_o,id_hold}),
    .f({_al_u6212_o,\ins_dec/mux13_b0_sel_is_0_o }));
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6213|ins_dec/reg7_b0  (
    .b({_al_u6212_o,_al_u4875_o}),
    .c({\ins_dec/mux19_b10_sel_is_2_o ,id_ins_pc[0]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[0],rs1_data[0]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u6213_o,open_n40366}),
    .q({open_n40370,as1[0]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6215|biu/bus_unit/mmu/reg2_b11  (
    .a({open_n40371,_al_u6215_o}),
    .b({\biu/bus_unit/mmu/i [0],_al_u6216_o}),
    .c({\biu/bus_unit/mmu/i [1],_al_u3034_o}),
    .clk(clk_pad),
    .d({\biu/maddress [20],\biu/paddress [75]}),
    .sr(rst_pad),
    .f({_al_u6215_o,open_n40389}),
    .q({open_n40393,\biu/paddress [75]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6218|biu/bus_unit/mmu/reg2_b10  (
    .a({open_n40394,_al_u6218_o}),
    .b({\biu/bus_unit/mmu/i [0],_al_u6219_o}),
    .c({\biu/bus_unit/mmu/i [1],_al_u3034_o}),
    .clk(clk_pad),
    .d({\biu/maddress [19],\biu/paddress [74]}),
    .sr(rst_pad),
    .f({_al_u6218_o,open_n40412}),
    .q({open_n40416,\biu/paddress [74]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6221|biu/bus_unit/mmu/reg2_b9  (
    .a({open_n40417,_al_u6221_o}),
    .b({\biu/bus_unit/mmu/i [0],_al_u6222_o}),
    .c({\biu/bus_unit/mmu/i [1],_al_u3034_o}),
    .clk(clk_pad),
    .d({\biu/maddress [18],\biu/paddress [73]}),
    .sr(rst_pad),
    .f({_al_u6221_o,open_n40435}),
    .q({open_n40439,\biu/paddress [73]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6224|biu/bus_unit/mmu/reg2_b8  (
    .a({open_n40440,_al_u6224_o}),
    .b({\biu/bus_unit/mmu/i [0],_al_u6225_o}),
    .c({\biu/bus_unit/mmu/i [1],_al_u3034_o}),
    .clk(clk_pad),
    .d({\biu/maddress [17],\biu/paddress [72]}),
    .sr(rst_pad),
    .f({_al_u6224_o,open_n40454}),
    .q({open_n40458,\biu/paddress [72]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6227|biu/bus_unit/mmu/reg2_b7  (
    .a({open_n40459,_al_u6227_o}),
    .b({\biu/bus_unit/mmu/i [0],_al_u6228_o}),
    .c({\biu/bus_unit/mmu/i [1],_al_u3034_o}),
    .clk(clk_pad),
    .d({\biu/maddress [16],\biu/paddress [71]}),
    .sr(rst_pad),
    .f({_al_u6227_o,open_n40473}),
    .q({open_n40477,\biu/paddress [71]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6230|biu/bus_unit/mmu/reg2_b6  (
    .a({open_n40478,_al_u6230_o}),
    .b({\biu/bus_unit/mmu/i [0],_al_u6231_o}),
    .c({\biu/bus_unit/mmu/i [1],_al_u3034_o}),
    .clk(clk_pad),
    .d({\biu/maddress [15],\biu/paddress [70]}),
    .sr(rst_pad),
    .f({_al_u6230_o,open_n40496}),
    .q({open_n40500,\biu/paddress [70]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6233|biu/bus_unit/mmu/reg2_b5  (
    .a({open_n40501,_al_u6233_o}),
    .b({\biu/bus_unit/mmu/i [0],_al_u6234_o}),
    .c({\biu/bus_unit/mmu/i [1],_al_u3034_o}),
    .clk(clk_pad),
    .d({\biu/maddress [14],\biu/paddress [69]}),
    .sr(rst_pad),
    .f({_al_u6233_o,open_n40519}),
    .q({open_n40523,\biu/paddress [69]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6236|biu/bus_unit/mmu/reg2_b4  (
    .a({open_n40524,_al_u6236_o}),
    .b({\biu/bus_unit/mmu/i [0],_al_u6237_o}),
    .c({\biu/bus_unit/mmu/i [1],_al_u3034_o}),
    .clk(clk_pad),
    .d({\biu/maddress [13],\biu/paddress [68]}),
    .sr(rst_pad),
    .f({_al_u6236_o,open_n40538}),
    .q({open_n40542,\biu/paddress [68]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6239|biu/bus_unit/mmu/reg2_b3  (
    .a({open_n40543,_al_u6239_o}),
    .b({\biu/bus_unit/mmu/i [0],_al_u6240_o}),
    .c({\biu/bus_unit/mmu/i [1],_al_u3034_o}),
    .clk(clk_pad),
    .d({\biu/maddress [12],\biu/paddress [67]}),
    .sr(rst_pad),
    .f({_al_u6239_o,open_n40557}),
    .q({open_n40561,\biu/paddress [67]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6243|biu/cache_ctrl_logic/reg3_b37  (
    .a({\biu/cache_ctrl_logic/l1d_va [37],\biu/cache_ctrl_logic/l1i_va [37]}),
    .b({\biu/cache_ctrl_logic/l1d_va [56],\biu/cache_ctrl_logic/l1i_va [61]}),
    .c({addr_ex[37],addr_ex[37]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[56],addr_ex[61]}),
    .mi({open_n40572,addr_ex[37]}),
    .sr(rst_pad),
    .f({_al_u6243_o,_al_u6396_o}),
    .q({open_n40576,\biu/cache_ctrl_logic/l1d_va [37]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6245|biu/cache_ctrl_logic/reg3_b20  (
    .a({\biu/cache_ctrl_logic/l1d_va [12],\biu/cache_ctrl_logic/l1i_va [20]}),
    .b({\biu/cache_ctrl_logic/l1d_va [20],\biu/cache_ctrl_logic/l1i_va [52]}),
    .c({addr_ex[12],addr_ex[20]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[20],addr_ex[52]}),
    .mi({open_n40580,addr_ex[20]}),
    .sr(rst_pad),
    .f({_al_u6245_o,_al_u6394_o}),
    .q({open_n40595,\biu/cache_ctrl_logic/l1d_va [20]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6251|biu/cache_ctrl_logic/reg3_b22  (
    .a({_al_u6246_o,open_n40596}),
    .b({_al_u6248_o,\biu/cache_ctrl_logic/l1d_va [22]}),
    .c({_al_u6249_o,addr_ex[22]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6250_o,_al_u6247_o}),
    .mi({open_n40600,addr_ex[22]}),
    .sr(rst_pad),
    .f({_al_u6251_o,_al_u6248_o}),
    .q({open_n40615,\biu/cache_ctrl_logic/l1d_va [22]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A*(D@B))"),
    //.LUT1("(~D*C*~B*~A)"),
    .INIT_LUT0(16'b0000000100000100),
    .INIT_LUT1(16'b0000000000010000),
    .MODE("LOGIC"))
    \_al_u6254|_al_u6252  (
    .a({\exu/main_state [0],\exu/main_state [0]}),
    .b({\exu/main_state [1],\exu/main_state [1]}),
    .c({\exu/main_state [2],\exu/main_state [2]}),
    .d({\exu/main_state [3],\exu/main_state [3]}),
    .f({_al_u6254_o,\exu/n59_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*A*(D@B))"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(~C*A*(D@B))"),
    //.LUTG1("(D*~C*B*A)"),
    .INIT_LUTF0(16'b0000001000001000),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b0000001000001000),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6255|_al_u7903  (
    .a({\exu/main_state [0],\exu/main_state [0]}),
    .b({\exu/main_state [1],\exu/main_state [1]}),
    .c({\exu/main_state [2],\exu/main_state [2]}),
    .d({\exu/main_state [3],\exu/main_state [3]}),
    .f({_al_u6255_o,\exu/n60_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6257|_al_u6253  (
    .c({write,load}),
    .d({read,\exu/n59_lutinv }),
    .f({_al_u6257_o,read}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(D*~(~C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6258|biu/cache_ctrl_logic/reg3_b44  (
    .a({open_n40684,\biu/cache_ctrl_logic/l1i_va [44]}),
    .b({\biu/cache_ctrl_logic/l1d_va [44],\biu/cache_ctrl_logic/l1i_va [52]}),
    .c({addr_ex[44],addr_ex[44]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_value ,addr_ex[52]}),
    .mi({open_n40695,addr_ex[44]}),
    .sr(rst_pad),
    .f({_al_u6258_o,_al_u6403_o}),
    .q({open_n40699,\biu/cache_ctrl_logic/l1d_va [44]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6265|biu/cache_ctrl_logic/reg3_b52  (
    .a({_al_u6261_o,\biu/cache_ctrl_logic/l1d_va [52]}),
    .b({_al_u6262_o,\biu/cache_ctrl_logic/l1d_va [57]}),
    .c({_al_u6263_o,addr_ex[52]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6264_o,addr_ex[57]}),
    .mi({open_n40703,addr_ex[52]}),
    .sr(rst_pad),
    .f({_al_u6265_o,_al_u6263_o}),
    .q({open_n40718,\biu/cache_ctrl_logic/l1d_va [52]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(D*C*B*~A)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(D*C*B*~A)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0100000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6270|_al_u9223  (
    .a({\biu/cache_ctrl_logic/eq1/xor_i0[4]_i1[4]_o_lutinv ,_al_u9219_o}),
    .b({_al_u6267_o,_al_u9220_o}),
    .c({_al_u6268_o,_al_u9221_o}),
    .d({_al_u6269_o,_al_u9222_o}),
    .f({_al_u6270_o,_al_u9223_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D@C))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000001000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6271|biu/cache_ctrl_logic/reg3_b55  (
    .a({open_n40743,_al_u6258_o}),
    .b({_al_u6265_o,_al_u6259_o}),
    .c({_al_u6270_o,\biu/cache_ctrl_logic/l1d_va [55]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6260_o,addr_ex[55]}),
    .mi({open_n40754,addr_ex[55]}),
    .sr(rst_pad),
    .f({_al_u6271_o,_al_u6260_o}),
    .q({open_n40758,\biu/cache_ctrl_logic/l1d_va [55]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6276|exu/reg3_b15  (
    .a({_al_u6272_o,\biu/cache_ctrl_logic/l1d_va [15]}),
    .b({_al_u6273_o,\biu/cache_ctrl_logic/l1d_va [25]}),
    .c({_al_u6274_o,addr_ex[15]}),
    .clk(clk_pad),
    .d({_al_u6275_o,addr_ex[25]}),
    .mi({open_n40770,addr_ex[15]}),
    .sr(rst_pad),
    .f({_al_u6276_o,_al_u6273_o}),
    .q({open_n40774,new_pc[15]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*A))"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100110001),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6278|biu/cache_ctrl_logic/reg3_b32  (
    .a({\biu/cache_ctrl_logic/l1d_va [28],\biu/cache_ctrl_logic/l1i_va [26]}),
    .b({\biu/cache_ctrl_logic/l1d_va [32],\biu/cache_ctrl_logic/l1i_va [32]}),
    .c({addr_ex[28],addr_ex[26]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[32],addr_ex[32]}),
    .mi({open_n40785,addr_ex[32]}),
    .sr(rst_pad),
    .f({_al_u6278_o,_al_u6410_o}),
    .q({open_n40789,\biu/cache_ctrl_logic/l1d_va [32]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6280|_al_u6308  (
    .a({open_n40790,_al_u6300_o}),
    .b({_al_u6278_o,_al_u6305_o}),
    .c({_al_u6279_o,_al_u6306_o}),
    .d({_al_u6277_o,_al_u6307_o}),
    .f({_al_u6280_o,_al_u6308_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6285|exu/reg3_b56  (
    .a({_al_u6281_o,\biu/cache_ctrl_logic/l1d_va [44]}),
    .b({_al_u6282_o,\biu/cache_ctrl_logic/l1d_va [56]}),
    .c({_al_u6283_o,addr_ex[44]}),
    .clk(clk_pad),
    .d({_al_u6284_o,addr_ex[56]}),
    .mi({open_n40815,addr_ex[56]}),
    .sr(rst_pad),
    .f({_al_u6285_o,_al_u6282_o}),
    .q({open_n40830,new_pc[56]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D@C))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000001000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6290|biu/cache_ctrl_logic/reg3_b59  (
    .a({_al_u6286_o,_al_u6380_o}),
    .b({_al_u6287_o,_al_u6381_o}),
    .c({_al_u6288_o,\biu/cache_ctrl_logic/l1i_va [59]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6289_o,addr_ex[59]}),
    .mi({open_n40841,addr_ex[59]}),
    .sr(rst_pad),
    .f({_al_u6290_o,_al_u6382_o}),
    .q({open_n40845,\biu/cache_ctrl_logic/l1d_va [59]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B*~A))"),
    //.LUTF1("(C*B*~D)"),
    //.LUTG0("(~D*~(C*~B*~A))"),
    //.LUTG1("(C*B*~D)"),
    .INIT_LUTF0(16'b0000000011101111),
    .INIT_LUTF1(16'b0000000011000000),
    .INIT_LUTG0(16'b0000000011101111),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6292|_al_u7159  (
    .a({open_n40846,_al_u7149_o}),
    .b({_al_u6271_o,_al_u6257_o}),
    .c({_al_u6291_o,\biu/cache_ctrl_logic/l1d_wr_sel_lutinv }),
    .d({_al_u6257_o,\biu/cache_ctrl_logic/n75_lutinv }),
    .f({_al_u6292_o,_al_u7159_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6298|biu/cache_ctrl_logic/reg3_b41  (
    .a({_al_u6294_o,\biu/cache_ctrl_logic/l1d_va [15]}),
    .b({_al_u6295_o,\biu/cache_ctrl_logic/l1d_va [41]}),
    .c({_al_u6296_o,addr_ex[15]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6297_o,addr_ex[41]}),
    .mi({open_n40874,addr_ex[41]}),
    .sr(rst_pad),
    .f({_al_u6298_o,_al_u6297_o}),
    .q({open_n40889,\biu/cache_ctrl_logic/l1d_va [41]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6305|exu/reg3_b26  (
    .a({_al_u6301_o,\biu/cache_ctrl_logic/l1d_va [17]}),
    .b({_al_u6302_o,\biu/cache_ctrl_logic/l1d_va [26]}),
    .c({_al_u6303_o,addr_ex[17]}),
    .clk(clk_pad),
    .d({_al_u6304_o,addr_ex[26]}),
    .mi({open_n40894,addr_ex[26]}),
    .sr(rst_pad),
    .f({_al_u6305_o,_al_u6301_o}),
    .q({open_n40909,new_pc[26]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6309|_al_u6421  (
    .a({_al_u6251_o,_al_u6388_o}),
    .b({_al_u6292_o,_al_u6400_o}),
    .c({_al_u6298_o,_al_u6420_o}),
    .d({_al_u6308_o,_al_u6257_o}),
    .f({_al_u6309_o,\biu/cache_ctrl_logic/ex_l1i_hit }));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(D*C)))"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100100010001000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6311|biu/cache_ctrl_logic/reg5_b2  (
    .a({open_n40934,\biu/cache_ctrl_logic/n34 }),
    .b({write,\biu/cache_ctrl_logic/n30 }),
    .c({\biu/cache_ctrl_logic/l1d_pte [2],write}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/n42 ,\biu/cache_ctrl_logic/l1d_pte [2]}),
    .mi({open_n40945,\biu/cache_ctrl_logic/pte_temp [2]}),
    .sr(rst_pad),
    .f({_al_u6311_o,\biu/cache_ctrl_logic/n36 }),
    .q({open_n40949,\biu/cache_ctrl_logic/l1d_pte [2]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6314|_al_u6313  (
    .c({priv[0],priv[3]}),
    .d({_al_u6313_o,priv[1]}),
    .f({\biu/bus_unit/mmu/n7_lutinv ,_al_u6313_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*B*~D)"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000000000001100),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6319|_al_u2963  (
    .b({\cu_ru/m_s_status/n5 [1],_al_u2698_o}),
    .c({priv[3],\biu/bus_unit/mmu/n31_lutinv }),
    .d({\biu/bus_unit/mmu/n31_lutinv ,_al_u2914_o}),
    .f({_al_u6319_o,_al_u2963_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(D*~B*~(C*~A))"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(D*~B*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0010001100000000),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0010001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6320|biu/cache_ctrl_logic/reg5_b4  (
    .a({_al_u6311_o,open_n41004}),
    .b({\biu/cache_ctrl_logic/n36 ,\biu/cache_ctrl_logic/l1d_pte [4]}),
    .c({\biu/cache_ctrl_logic/n40 ,sum}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6319_o,\biu/bus_unit/mmu/n8_lutinv }),
    .mi({open_n41008,\biu/cache_ctrl_logic/pte_temp [4]}),
    .sr(rst_pad),
    .f({_al_u6320_o,\biu/cache_ctrl_logic/n40 }),
    .q({open_n41023,\biu/cache_ctrl_logic/l1d_pte [4]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u6321|_al_u9283  (
    .b({open_n41026,_al_u6257_o}),
    .c({_al_u6320_o,\biu/cache_ctrl_logic/n55_lutinv }),
    .d({_al_u6309_o,_al_u6309_o}),
    .f({_al_u6321_o,_al_u9283_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0001001111011111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0001001111011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6323|_al_u7197  (
    .a({_al_u6321_o,open_n41047}),
    .b({\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ,open_n41048}),
    .c({write,write}),
    .d({\biu/cache_write_lutinv ,\biu/cache_ctrl_logic/n75_lutinv }),
    .f({_al_u6323_o,\biu/bus_unit/mmu/n12_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6326|_al_u6332  (
    .b({open_n41075,\exu/lsu/n8_lutinv }),
    .c({\biu/cache_ctrl_logic/n174_lutinv ,addr_ex[2]}),
    .d({\biu/cache_ctrl_logic/n176_lutinv ,\biu/cache_ctrl_logic/n176_lutinv }),
    .f({_al_u6326_o,\biu/cache_ctrl_logic/n189 [2]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~A*~(~D*C*B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~A*~(~D*C*B))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0101010100010101),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0101010100010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6331|_al_u6330  (
    .a({\biu/cache_ctrl_logic/n189 [6],open_n41096}),
    .b({\biu/cache_ctrl_logic/n176_lutinv ,open_n41097}),
    .c({\exu/lsu/n5_lutinv ,addr_ex[1]}),
    .d({addr_ex[2],addr_ex[0]}),
    .f({_al_u6331_o,\exu/lsu/n5_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*~A)"),
    //.LUT1("(~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"))
    \_al_u6333|_al_u6325  (
    .a({ex_size[0],ex_size[0]}),
    .b({ex_size[1],ex_size[1]}),
    .c({ex_size[2],ex_size[2]}),
    .d({ex_size[3],ex_size[3]}),
    .f({\biu/cache_ctrl_logic/n173_lutinv ,\biu/cache_ctrl_logic/n174_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*A*~(D*C))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000001000100010),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u6334|_al_u8944  (
    .a({open_n41142,_al_u8941_o}),
    .b({open_n41143,_al_u8943_o}),
    .c({\biu/cache_ctrl_logic/n173_lutinv ,_al_u8779_o}),
    .d({\biu/cache_ctrl_logic/n174_lutinv ,\exu/lsu/n5_lutinv }),
    .f({_al_u6334_o,_al_u8944_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~D)"),
    //.LUT1("(~D*~C*B*~A)"),
    .INIT_LUT0(16'b0000000011000000),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("LOGIC"))
    \_al_u6336|_al_u6327  (
    .a({\biu/cache_ctrl_logic/n185 [3],open_n41164}),
    .b({_al_u6331_o,\exu/lsu/n0_lutinv }),
    .c({\biu/cache_ctrl_logic/n189 [2],addr_ex[2]}),
    .d({\biu/cache_ctrl_logic/n182 [4],_al_u6326_o}),
    .f({_al_u6336_o,\biu/cache_ctrl_logic/n185 [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u6337|_al_u6430  (
    .b({\biu/cache_ctrl_logic/n55_lutinv ,\biu/cache_ctrl_logic/n55_lutinv }),
    .c({_al_u6336_o,_al_u6336_o}),
    .d({_al_u6323_o,\biu/l1i_write_lutinv }),
    .f({\biu/cache/n11 ,\biu/cache/n27 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000011000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6339|_al_u6335  (
    .b({open_n41209,\exu/lsu/n2_lutinv }),
    .c({_al_u6334_o,addr_ex[2]}),
    .d({\biu/cache_ctrl_logic/n176_lutinv ,_al_u6334_o}),
    .f({_al_u6339_o,\biu/cache_ctrl_logic/n182 [4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*B*~(D)+~(A)*~(B)*D+A*~(B)*D))"),
    //.LUTF1("(~B*A*~(D*~C))"),
    //.LUTG0("(~C*(A*B*~(D)+~(A)*~(B)*D+A*~(B)*D))"),
    //.LUTG1("(~B*A*~(D*~C))"),
    .INIT_LUTF0(16'b0000001100001000),
    .INIT_LUTF1(16'b0010000000100010),
    .INIT_LUTG0(16'b0000001100001000),
    .INIT_LUTG1(16'b0010000000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6341|_al_u6340  (
    .a({_al_u6331_o,\biu/cache_ctrl_logic/n176_lutinv }),
    .b({\biu/cache_ctrl_logic/n185 [2],addr_ex[0]}),
    .c({_al_u6339_o,addr_ex[1]}),
    .d({_al_u6340_o,addr_ex[2]}),
    .f({_al_u6341_o,_al_u6340_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6342|_al_u6431  (
    .b({\biu/cache_ctrl_logic/n55_lutinv ,\biu/cache_ctrl_logic/n55_lutinv }),
    .c({_al_u6341_o,_al_u6341_o}),
    .d({_al_u6323_o,\biu/l1i_write_lutinv }),
    .f({\biu/cache/n9 ,\biu/cache/n25 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(~C*B*~D)"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"))
    \_al_u6343|_al_u6338  (
    .b({\exu/lsu/n8_lutinv ,\exu/lsu/n8_lutinv }),
    .c({addr_ex[2],addr_ex[2]}),
    .d({_al_u6339_o,_al_u6326_o}),
    .f({\biu/cache_ctrl_logic/n182 [2],\biu/cache_ctrl_logic/n185 [2]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(B*A*(D@C))"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(B*A*(D@C))"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000100010000000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b0000100010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6345|_al_u6329  (
    .a({\biu/cache_ctrl_logic/n172_lutinv ,\biu/cache_ctrl_logic/n172_lutinv }),
    .b({_al_u3415_o,_al_u3415_o}),
    .c({ex_size[2],ex_size[2]}),
    .d({ex_size[3],ex_size[3]}),
    .f({\biu/cache_ctrl_logic/n189 [5],\biu/cache_ctrl_logic/n189 [6]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(~B*~D))"),
    //.LUTF1("(~D*~A*~(C*~B))"),
    //.LUTG0("(~C*~(~B*~D))"),
    //.LUTG1("(~D*~A*~(C*~B))"),
    .INIT_LUTF0(16'b0000111100001100),
    .INIT_LUTF1(16'b0000000001000101),
    .INIT_LUTG0(16'b0000111100001100),
    .INIT_LUTG1(16'b0000000001000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6346|_al_u6344  (
    .a({\biu/cache_ctrl_logic/n182 [2],open_n41326}),
    .b({_al_u6326_o,addr_ex[1]}),
    .c({_al_u6344_o,addr_ex[2]}),
    .d({\biu/cache_ctrl_logic/n189 [5],\biu/cache_ctrl_logic/n176_lutinv }),
    .f({_al_u6346_o,_al_u6344_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6347|_al_u6432  (
    .b({\biu/cache_ctrl_logic/n55_lutinv ,\biu/cache_ctrl_logic/n55_lutinv }),
    .c({_al_u6346_o,_al_u6346_o}),
    .d({_al_u6323_o,\biu/l1i_write_lutinv }),
    .f({\biu/cache/n7 ,\biu/cache/n23 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~D*C*~A))"),
    //.LUT1("(A*~(~D*C*~B))"),
    .INIT_LUT0(16'b0011001100100011),
    .INIT_LUT1(16'b1010101010001010),
    .MODE("LOGIC"))
    \_al_u6349|_al_u6348  (
    .a({_al_u6348_o,_al_u6326_o}),
    .b({_al_u6339_o,\biu/cache_ctrl_logic/n189 [5]}),
    .c({\exu/lsu/n5_lutinv ,\exu/lsu/n2_lutinv }),
    .d({addr_ex[2],addr_ex[2]}),
    .f({_al_u6349_o,_al_u6348_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u6350|_al_u6433  (
    .b({\biu/cache_ctrl_logic/n55_lutinv ,\biu/cache_ctrl_logic/n55_lutinv }),
    .c({_al_u6349_o,_al_u6349_o}),
    .d({_al_u6323_o,\biu/l1i_write_lutinv }),
    .f({\biu/cache/n5 ,\biu/cache/n21 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6351|_al_u6328  (
    .b({\biu/cache_ctrl_logic/n189 [6],open_n41421}),
    .c({\biu/cache_ctrl_logic/n172_lutinv ,addr_ex[2]}),
    .d({_al_u6326_o,\exu/lsu/n0_lutinv }),
    .f({_al_u6351_o,\biu/cache_ctrl_logic/n172_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*C*~B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(A*~(~D*C*~B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b1010101010001010),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1010101010001010),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6353|_al_u6352  (
    .a({open_n41446,_al_u6351_o}),
    .b({\biu/cache_ctrl_logic/n55_lutinv ,_al_u6339_o}),
    .c({_al_u6352_o,\exu/lsu/n2_lutinv }),
    .d({_al_u6323_o,addr_ex[2]}),
    .f({\biu/cache/n3 ,_al_u6352_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111111011101001),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111011101001),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6355|_al_u6354  (
    .a({open_n41471,ex_size[0]}),
    .b({open_n41472,ex_size[1]}),
    .c({_al_u6354_o,ex_size[2]}),
    .d({\biu/cache_ctrl_logic/n172_lutinv ,ex_size[3]}),
    .f({\biu/cache_ctrl_logic/ex_bsel [0],_al_u6354_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(~D*~(~C*B))"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(~D*~(~C*B))"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0000000011110011),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0000000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6356|_al_u6435  (
    .b({\biu/cache_ctrl_logic/n55_lutinv ,\biu/cache_ctrl_logic/n55_lutinv }),
    .c({\biu/cache_ctrl_logic/ex_bsel [0],\biu/cache_ctrl_logic/ex_bsel [0]}),
    .d({_al_u6323_o,\biu/l1i_write_lutinv }),
    .f({\biu/cache/n1 ,\biu/cache/n17 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*B))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001010101010101),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6358|_al_u6359  (
    .a({open_n41523,\biu/cache_ctrl_logic/n185 [5]}),
    .b({\biu/cache_ctrl_logic/n174_lutinv ,\exu/lsu/n8_lutinv }),
    .c({addr_ex[2],\biu/cache_ctrl_logic/n173_lutinv }),
    .d({\exu/lsu/n5_lutinv ,addr_ex[2]}),
    .f({\biu/cache_ctrl_logic/n185 [5],_al_u6359_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~A*~(D*C*B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001010101010101),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6360|_al_u6357  (
    .a({open_n41544,\biu/cache_ctrl_logic/n189 [6]}),
    .b({open_n41545,\biu/cache_ctrl_logic/n176_lutinv }),
    .c({_al_u6359_o,\exu/lsu/n0_lutinv }),
    .d({_al_u6357_o,addr_ex[2]}),
    .f({_al_u6360_o,_al_u6357_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*B*~(C)+~(A)*~(B)*C+A*~(B)*C))"),
    //.LUT1("(~B*A*~(D*~C))"),
    .INIT_LUT0(16'b0011100000000000),
    .INIT_LUT1(16'b0010000000100010),
    .MODE("LOGIC"))
    \_al_u6363|_al_u6362  (
    .a({_al_u6357_o,\biu/cache_ctrl_logic/n174_lutinv }),
    .b({\biu/cache_ctrl_logic/n189 [2],addr_ex[0]}),
    .c({_al_u6334_o,addr_ex[1]}),
    .d({_al_u6362_o,addr_ex[2]}),
    .f({_al_u6363_o,_al_u6362_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u6364|_al_u6429  (
    .b({\biu/cache_ctrl_logic/n55_lutinv ,\biu/cache_ctrl_logic/n55_lutinv }),
    .c({_al_u6363_o,_al_u6363_o}),
    .d({_al_u6323_o,\biu/l1i_write_lutinv }),
    .f({\biu/cache/n13 ,\biu/cache/n29 }));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6369|biu/cache_ctrl_logic/reg3_b38  (
    .a({_al_u6365_o,\biu/cache_ctrl_logic/l1i_va [38]}),
    .b({_al_u6366_o,\biu/cache_ctrl_logic/l1i_va [63]}),
    .c({_al_u6367_o,addr_ex[38]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6368_o,addr_ex[63]}),
    .mi({open_n41615,addr_ex[38]}),
    .sr(rst_pad),
    .f({_al_u6369_o,_al_u6366_o}),
    .q({open_n41630,\biu/cache_ctrl_logic/l1d_va [38]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6378|biu/cache_ctrl_logic/reg3_b27  (
    .a({_al_u6373_o,\biu/cache_ctrl_logic/l1i_va [27]}),
    .b({_al_u6375_o,\biu/cache_ctrl_logic/l1i_va [35]}),
    .c({_al_u6376_o,addr_ex[27]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6377_o,addr_ex[35]}),
    .mi({open_n41634,addr_ex[27]}),
    .sr(rst_pad),
    .f({_al_u6378_o,_al_u6377_o}),
    .q({open_n41649,\biu/cache_ctrl_logic/l1d_va [27]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6387|biu/cache_ctrl_logic/reg3_b50  (
    .a({_al_u6383_o,\biu/cache_ctrl_logic/l1i_va [50]}),
    .b({_al_u6384_o,\biu/cache_ctrl_logic/l1i_va [54]}),
    .c({_al_u6385_o,addr_ex[50]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6386_o,addr_ex[54]}),
    .mi({open_n41660,addr_ex[50]}),
    .sr(rst_pad),
    .f({_al_u6387_o,_al_u6384_o}),
    .q({open_n41664,\biu/cache_ctrl_logic/l1d_va [50]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*~C))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000010001000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6388|biu/cache_ctrl_logic/reg3_b58  (
    .a({_al_u6371_o,_al_u6369_o}),
    .b({_al_u6378_o,_al_u6370_o}),
    .c({_al_u6382_o,\biu/cache_ctrl_logic/l1i_va [58]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6387_o,addr_ex[58]}),
    .mi({open_n41675,addr_ex[58]}),
    .sr(rst_pad),
    .f({_al_u6388_o,_al_u6371_o}),
    .q({open_n41679,\biu/cache_ctrl_logic/l1d_va [58]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6395|biu/cache_ctrl_logic/reg3_b12  (
    .a({_al_u6391_o,\biu/cache_ctrl_logic/l1i_va [12]}),
    .b({_al_u6392_o,\biu/cache_ctrl_logic/l1i_va [20]}),
    .c({_al_u6393_o,addr_ex[12]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6394_o,addr_ex[20]}),
    .mi({open_n41690,addr_ex[12]}),
    .sr(rst_pad),
    .f({_al_u6395_o,_al_u6393_o}),
    .q({open_n41694,\biu/cache_ctrl_logic/l1d_va [12]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6400|biu/cache_ctrl_logic/reg3_b19  (
    .a({_al_u6395_o,\biu/cache_ctrl_logic/l1i_va [19]}),
    .b({_al_u6397_o,\biu/cache_ctrl_logic/l1i_va [41]}),
    .c({_al_u6398_o,addr_ex[19]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6399_o,addr_ex[41]}),
    .mi({open_n41705,addr_ex[19]}),
    .sr(rst_pad),
    .f({_al_u6400_o,_al_u6399_o}),
    .q({open_n41709,\biu/cache_ctrl_logic/l1d_va [19]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6409|biu/cache_ctrl_logic/reg3_b46  (
    .a({_al_u6405_o,\biu/cache_ctrl_logic/l1i_va [46]}),
    .b({_al_u6406_o,\biu/cache_ctrl_logic/l1i_va [62]}),
    .c({_al_u6407_o,addr_ex[46]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6408_o,addr_ex[62]}),
    .mi({open_n41713,addr_ex[46]}),
    .sr(rst_pad),
    .f({_al_u6409_o,_al_u6408_o}),
    .q({open_n41728,\biu/cache_ctrl_logic/l1d_va [46]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6414|biu/cache_ctrl_logic/reg3_b30  (
    .a({_al_u6409_o,\biu/cache_ctrl_logic/l1i_va [30]}),
    .b({_al_u6411_o,\biu/cache_ctrl_logic/l1i_va [42]}),
    .c({_al_u6412_o,addr_ex[30]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6413_o,addr_ex[42]}),
    .mi({open_n41732,addr_ex[30]}),
    .sr(rst_pad),
    .f({_al_u6414_o,_al_u6412_o}),
    .q({open_n41747,\biu/cache_ctrl_logic/l1d_va [30]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6419|biu/cache_ctrl_logic/reg3_b34  (
    .a({_al_u6415_o,\biu/cache_ctrl_logic/l1i_va [17]}),
    .b({_al_u6416_o,\biu/cache_ctrl_logic/l1i_va [34]}),
    .c({_al_u6417_o,addr_ex[17]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6418_o,addr_ex[34]}),
    .mi({open_n41758,addr_ex[34]}),
    .sr(rst_pad),
    .f({_al_u6419_o,_al_u6415_o}),
    .q({open_n41762,\biu/cache_ctrl_logic/l1d_va [34]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D@C))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(B*A*~(D@C))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000001000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1000000000001000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6420|biu/cache_ctrl_logic/reg3_b49  (
    .a({open_n41763,_al_u6402_o}),
    .b({_al_u6414_o,_al_u6403_o}),
    .c({_al_u6419_o,\biu/cache_ctrl_logic/l1i_va [49]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6404_o,addr_ex[49]}),
    .mi({open_n41767,addr_ex[49]}),
    .sr(rst_pad),
    .f({_al_u6420_o,_al_u6404_o}),
    .q({open_n41782,\biu/cache_ctrl_logic/l1d_va [49]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(A*~(~B*~(D*C)))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1010100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6422|cu_ru/m_s_status/mxr_reg  (
    .a({read,open_n41783}),
    .b({\biu/cache_ctrl_logic/l1i_pte [1],open_n41784}),
    .c({\biu/cache_ctrl_logic/l1i_pte [3],_al_u3427_o}),
    .ce(\cu_ru/m_s_status/u34_sel_is_0_o ),
    .clk(clk_pad),
    .d({mxr,\cu_ru/m_s_status/n0 }),
    .mi({open_n41795,data_csr[19]}),
    .sr(rst_pad),
    .f({\biu/cache_ctrl_logic/n17 ,\cu_ru/m_s_status/u34_sel_is_0_o }),
    .q({open_n41799,mxr}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6423|cu_ru/m_s_status/sum_reg  (
    .a({\biu/bus_unit/mmu/n7_lutinv ,\cu_ru/read_sscratch_sel_lutinv }),
    .b({\biu/bus_unit/mmu/n8_lutinv ,\cu_ru/n90 [32]}),
    .c({\biu/cache_ctrl_logic/l1i_pte [4],\cu_ru/sscratch [18]}),
    .ce(\cu_ru/m_s_status/u34_sel_is_0_o ),
    .clk(clk_pad),
    .d({sum,sum}),
    .mi({open_n41810,data_csr[18]}),
    .sr(rst_pad),
    .f({_al_u6423_o,_al_u7634_o}),
    .q({open_n41814,sum}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~A*~(D*C)))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0011001000100010),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6425|_al_u6424  (
    .a({open_n41815,\biu/cache_ctrl_logic/n17 }),
    .b({open_n41816,_al_u6423_o}),
    .c({_al_u6319_o,write}),
    .d({\biu/cache_ctrl_logic/n26_lutinv ,\biu/cache_ctrl_logic/l1i_pte [2]}),
    .f({_al_u6425_o,\biu/cache_ctrl_logic/n26_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001111000000),
    .MODE("LOGIC"))
    \_al_u6427|_al_u2888  (
    .b({_al_u2886_o,open_n41839}),
    .c({\biu/cache_write_lutinv ,\biu/cache_ctrl_logic/l1d_wr_sel_lutinv }),
    .d({_al_u6426_o,_al_u2886_o}),
    .f({\biu/l1i_write_lutinv ,\biu/bus_unit/mux1_b1_sel_is_0_o }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u6428|_al_u6434  (
    .b({\biu/cache_ctrl_logic/n55_lutinv ,\biu/cache_ctrl_logic/n55_lutinv }),
    .c({_al_u6360_o,_al_u6352_o}),
    .d({\biu/l1i_write_lutinv ,\biu/l1i_write_lutinv }),
    .f({\biu/cache/n31 ,\biu/cache/n19 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~A*~(~D*~(~C*B)))"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0101010100000100),
    .MODE("LOGIC"))
    \_al_u6438|_al_u6437  (
    .a({_al_u4138_o,\cu_ru/mideleg_int_ctrl/sei_ack_m }),
    .b({\cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ,\cu_ru/m_s_status/n5 [1]}),
    .c({\cu_ru/mideleg_int_ctrl/n33_neg_lutinv ,_al_u3244_o}),
    .d({_al_u4139_o,\cu_ru/mstatus [1]}),
    .f({_al_u6438_o,\cu_ru/mideleg_int_ctrl/n33_neg_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUT1("~(~C*~(B*~(~D*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001111),
    .INIT_LUT1(16'b1111110011111000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6439|cu_ru/m_s_cause/reg1_b3  (
    .a({_al_u6436_o,open_n41902}),
    .b({_al_u4142_o,\cu_ru/trap_cause [3]}),
    .c({_al_u6438_o,\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u4143_o,_al_u6727_o}),
    .sr(rst_pad),
    .f({\cu_ru/trap_cause [3],open_n41916}),
    .q({open_n41920,\cu_ru/mcause [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6440|_al_u6057  (
    .c({_al_u3204_o,rst_pad}),
    .d({_al_u5992_o,\cu_ru/trap_target_m }),
    .f({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_cause/mux7_b10_sel_is_0_o }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6567|cu_ru/m_s_tval/reg1_b0  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,open_n41945}),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [0],\cu_ru/m_s_tval/n3 [0]}),
    .clk(clk_pad),
    .d({data_csr[0],_al_u6567_o}),
    .sr(rst_pad),
    .f({_al_u6567_o,open_n41963}),
    .q({open_n41967,\cu_ru/mtval [0]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6704|_al_u9268  (
    .b({open_n41970,_al_u9265_o}),
    .c({_al_u6425_o,\biu/cache_ctrl_logic/n55_lutinv }),
    .d({\biu/cache_ctrl_logic/ex_l1i_hit ,_al_u6704_o}),
    .f({_al_u6704_o,_al_u9268_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u6705|_al_u7193  (
    .b({open_n41997,\biu/cache_ctrl_logic/n55_lutinv }),
    .c({_al_u6704_o,write}),
    .d({_al_u6321_o,_al_u6321_o}),
    .f({\biu/ex_data_sel [0],_al_u7193_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("~(~D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6707|exu/reg3_b11  (
    .a({open_n42018,\biu/ex_data_sel [0]}),
    .b({\biu/bus_unit/mux1_b1_sel_is_0_o ,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .c({_al_u2891_o,addr_ex[11]}),
    .clk(clk_pad),
    .d({_al_u6706_o,addr_if[11]}),
    .mi({open_n42030,addr_ex[11]}),
    .sr(rst_pad),
    .f({\biu/l1i_addr [8],_al_u6706_o}),
    .q({open_n42034,new_pc[11]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("~(~D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6709|exu/reg3_b10  (
    .a({open_n42035,\biu/ex_data_sel [0]}),
    .b({\biu/bus_unit/mux1_b1_sel_is_0_o ,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .c({_al_u2893_o,addr_ex[10]}),
    .clk(clk_pad),
    .d({_al_u6708_o,addr_if[10]}),
    .mi({open_n42047,addr_ex[10]}),
    .sr(rst_pad),
    .f({\biu/l1i_addr [7],_al_u6708_o}),
    .q({open_n42051,new_pc[10]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6711|exu/reg3_b9  (
    .a({open_n42052,\biu/ex_data_sel [0]}),
    .b({\biu/bus_unit/mux1_b1_sel_is_0_o ,\biu/bus_unit/mux1_b1_sel_is_0_o }),
    .c({_al_u2895_o,addr_ex[9]}),
    .clk(clk_pad),
    .d({_al_u6710_o,addr_if[9]}),
    .mi({open_n42057,addr_ex[9]}),
    .sr(rst_pad),
    .f({\biu/l1i_addr [6],_al_u6710_o}),
    .q({open_n42072,new_pc[9]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b0011001100001111),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6713|exu/reg3_b8  (
    .b({\biu/bus_unit/mux1_b1_sel_is_0_o ,addr_ex[8]}),
    .c({_al_u2897_o,addr_if[8]}),
    .clk(clk_pad),
    .d({_al_u6712_o,\biu/ex_data_sel [0]}),
    .mi({open_n42079,addr_ex[8]}),
    .sr(rst_pad),
    .f({\biu/l1i_addr [5],_al_u6712_o}),
    .q({open_n42094,new_pc[8]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b0011001100001111),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6715|exu/reg3_b7  (
    .b({\biu/bus_unit/mux1_b1_sel_is_0_o ,addr_ex[7]}),
    .c({_al_u2899_o,addr_if[7]}),
    .clk(clk_pad),
    .d({_al_u6714_o,\biu/ex_data_sel [0]}),
    .mi({open_n42101,addr_ex[7]}),
    .sr(rst_pad),
    .f({\biu/l1i_addr [4],_al_u6714_o}),
    .q({open_n42116,new_pc[7]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001100001111),
    .INIT_LUT1(16'b0011000011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6717|exu/reg3_b6  (
    .b({\biu/bus_unit/mux1_b1_sel_is_0_o ,addr_ex[6]}),
    .c({_al_u2901_o,addr_if[6]}),
    .clk(clk_pad),
    .d({_al_u6716_o,\biu/ex_data_sel [0]}),
    .mi({open_n42130,addr_ex[6]}),
    .sr(rst_pad),
    .f({\biu/l1i_addr [3],_al_u6716_o}),
    .q({open_n42134,new_pc[6]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001100001111),
    .INIT_LUT1(16'b0011000011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6719|exu/reg3_b5  (
    .b({\biu/bus_unit/mux1_b1_sel_is_0_o ,addr_ex[5]}),
    .c({_al_u2903_o,addr_if[5]}),
    .clk(clk_pad),
    .d({_al_u6718_o,\biu/ex_data_sel [0]}),
    .mi({open_n42148,addr_ex[5]}),
    .sr(rst_pad),
    .f({\biu/l1i_addr [2],_al_u6718_o}),
    .q({open_n42152,new_pc[5]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b0011001100001111),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6721|exu/reg3_b4  (
    .b({\biu/bus_unit/mux1_b1_sel_is_0_o ,addr_ex[4]}),
    .c({_al_u2905_o,addr_if[4]}),
    .clk(clk_pad),
    .d({_al_u6720_o,\biu/ex_data_sel [0]}),
    .mi({open_n42159,addr_ex[4]}),
    .sr(rst_pad),
    .f({\biu/l1i_addr [1],_al_u6720_o}),
    .q({open_n42174,new_pc[4]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b0011001100001111),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6723|exu/reg3_b3  (
    .b({\biu/bus_unit/mux1_b1_sel_is_0_o ,addr_ex[3]}),
    .c({_al_u2907_o,addr_if[3]}),
    .clk(clk_pad),
    .d({_al_u6722_o,\biu/ex_data_sel [0]}),
    .mi({open_n42181,addr_ex[3]}),
    .sr(rst_pad),
    .f({\biu/l1i_addr [0],_al_u6722_o}),
    .q({open_n42196,new_pc[3]}));  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(~(D*C)*~(B*A))"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(~(D*C)*~(B*A))"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0000011101110111),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b0000011101110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6724|_al_u6426  (
    .a({_al_u6309_o,open_n42197}),
    .b({_al_u6320_o,_al_u6425_o}),
    .c({\biu/cache_ctrl_logic/ex_l1i_hit ,write}),
    .d({_al_u6425_o,\biu/cache_ctrl_logic/ex_l1i_hit }),
    .f({_al_u6724_o,_al_u6426_o}));
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6733|exu/reg3_b1  (
    .b({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6731_o}),
    .c({\cu_ru/stvec [3],new_pc[1]}),
    .clk(clk_pad),
    .d({_al_u6732_o,_al_u6055_o}),
    .mi({open_n42235,addr_ex[1]}),
    .sr(rst_pad),
    .f({_al_u6733_o,_al_u6732_o}),
    .q({open_n42239,new_pc[1]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6734|cu_ru/m_s_epc/reg0_b1  (
    .b({open_n42242,_al_u5157_o}),
    .c({\cu_ru/sepc [1],_al_u5604_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u2844_o,\cu_ru/m_s_epc/n2 [1]}),
    .sr(rst_pad),
    .f({_al_u6734_o,open_n42259}),
    .q({open_n42263,\cu_ru/sepc [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(B*~(C*D))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000110011001100),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6738|exu/reg3_b0  (
    .b({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6736_o}),
    .c({\cu_ru/stvec [2],new_pc[0]}),
    .clk(clk_pad),
    .d({_al_u6737_o,_al_u6055_o}),
    .mi({open_n42270,addr_ex[0]}),
    .sr(rst_pad),
    .f({_al_u6738_o,_al_u6737_o}),
    .q({open_n42285,new_pc[0]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000100000001),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6739|ins_fetch/reg2_b0  (
    .a({open_n42286,_al_u6738_o}),
    .b({open_n42287,_al_u6739_o}),
    .c({\cu_ru/sepc [0],\cu_ru/m_s_status/n2 }),
    .ce(pip_flush),
    .clk(clk_pad),
    .d({_al_u2844_o,\cu_ru/mepc [0]}),
    .sr(rst_pad),
    .f({_al_u6739_o,open_n42300}),
    .q({open_n42304,addr_if[0]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u6742|_al_u6741  (
    .b({\cu_ru/m_s_status/n2 ,open_n42307}),
    .c({\cu_ru/mstatus [7],1'b0}),
    .d({_al_u3427_o,\cu_ru/trap_target_m }),
    .f({_al_u6742_o,\cu_ru/m_s_status/mux3_b0_sel_is_2_o }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_LSLICE #(
    //.LUTF0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUTF1("(B*~(D*~C*~A))"),
    //.LUTG0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUTG1("(B*~(D*~C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000100000001),
    .INIT_LUTF1(16'b1100100011001100),
    .INIT_LUTG0(16'b1111000100000001),
    .INIT_LUTG1(16'b1100100011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6743|cu_ru/m_s_status/mie_reg  (
    .a({\cu_ru/m_s_status/mux3_b0_sel_is_2_o ,_al_u6743_o}),
    .b({_al_u6742_o,_al_u6744_o}),
    .c({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n0 }),
    .clk(clk_pad),
    .d({\cu_ru/mie ,data_csr[3]}),
    .sr(rst_pad),
    .f({_al_u6743_o,open_n42345}),
    .q({open_n42349,\cu_ru/mie }));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6744|_al_u6746  (
    .c({\cu_ru/mie ,\cu_ru/m_s_status/n2 }),
    .d({_al_u3427_o,_al_u3427_o}),
    .f({_al_u6744_o,_al_u6746_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b1100010010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6747|cu_ru/m_s_status/mpie_reg  (
    .a({\cu_ru/m_s_status/mux3_b0_sel_is_2_o ,_al_u6747_o}),
    .b({_al_u6746_o,_al_u6748_o}),
    .c({\cu_ru/mie ,\cu_ru/m_s_status/n0 }),
    .clk(clk_pad),
    .d({\cu_ru/mstatus [7],data_csr[7]}),
    .sr(rst_pad),
    .f({_al_u6747_o,open_n42391}),
    .q({open_n42395,\cu_ru/mstatus [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6748|_al_u9533  (
    .c({\cu_ru/mstatus [7],\cu_ru/mepc [31]}),
    .d({_al_u3427_o,\cu_ru/m_s_status/n2 }),
    .f({_al_u6748_o,_al_u9533_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(B*~(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0100110000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6751|cu_ru/m_s_status/reg0_b1  (
    .a({\cu_ru/m_s_status/mux3_b0_sel_is_2_o ,_al_u6751_o}),
    .b({_al_u6746_o,_al_u6752_o}),
    .c({_al_u6750_o,\cu_ru/m_s_status/n0 }),
    .clk(clk_pad),
    .d({\cu_ru/mstatus [12],data_csr[12]}),
    .sr(rst_pad),
    .f({_al_u6751_o,open_n42437}),
    .q({open_n42441,\cu_ru/mstatus [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(B*~(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0100110000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6754|cu_ru/m_s_status/reg0_b0  (
    .a({\cu_ru/m_s_status/mux3_b0_sel_is_2_o ,_al_u6754_o}),
    .b({_al_u6746_o,_al_u6755_o}),
    .c({_al_u6313_o,\cu_ru/m_s_status/n0 }),
    .clk(clk_pad),
    .d({\cu_ru/mstatus [11],data_csr[11]}),
    .sr(rst_pad),
    .f({_al_u6754_o,open_n42455}),
    .q({open_n42459,\cu_ru/mstatus [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6755|_al_u2841  (
    .c({\cu_ru/mstatus [11],\cu_ru/mstatus [11]}),
    .d({_al_u3427_o,\cu_ru/m_s_status/n2 }),
    .f({_al_u6755_o,_al_u2841_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(~D*C*~B*A)"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"))
    \_al_u6758|_al_u7478  (
    .a({_al_u3393_o,_al_u3393_o}),
    .b({id_ins[22],id_ins[22]}),
    .c({id_ins[21],id_ins[21]}),
    .d({id_ins[20],id_ins[20]}),
    .f({_al_u6758_o,_al_u7478_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6759|_al_u6757  (
    .a({open_n42508,_al_u3400_o}),
    .b({open_n42509,id_ins[31]}),
    .c({_al_u6758_o,id_ins[30]}),
    .d({_al_u6757_o,id_ins[29]}),
    .f({\cu_ru/read_minstret_sel_lutinv ,_al_u6757_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6761|_al_u6791  (
    .a({open_n42534,id_ins[29]}),
    .b({_al_u6760_o,id_ins[28]}),
    .c({_al_u3387_o,_al_u3387_o}),
    .d({\ins_dec/n80_lutinv ,_al_u3388_o}),
    .f({_al_u6761_o,_al_u6791_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6762|_al_u6782  (
    .c({_al_u6758_o,_al_u6761_o}),
    .d({_al_u6761_o,_al_u3395_o}),
    .f({\cu_ru/read_instret_sel_lutinv ,\cu_ru/read_time_sel_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*~A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~(C*B)*~(D*~A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0010101000111111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0010101000111111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6763|_al_u7698  (
    .a({open_n42583,_al_u6763_o}),
    .b({open_n42584,\cu_ru/read_time_sel_lutinv }),
    .c({\cu_ru/read_instret_sel_lutinv ,mtime_pad[2]}),
    .d({\cu_ru/read_minstret_sel_lutinv ,\cu_ru/minstret [2]}),
    .f({_al_u6763_o,_al_u7698_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6766|_al_u6765  (
    .b({id_ins[29],id_ins[27]}),
    .c({_al_u3388_o,id_ins[26]}),
    .d({_al_u6765_o,id_ins[28]}),
    .f({_al_u6766_o,_al_u6765_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6767|_al_u7726  (
    .a({open_n42635,\cu_ru/read_mtval_sel_lutinv }),
    .b({open_n42636,\cu_ru/read_time_sel_lutinv }),
    .c({_al_u6766_o,mtime_pad[0]}),
    .d({_al_u6764_o,\cu_ru/mtval [0]}),
    .f({\cu_ru/read_mtval_sel_lutinv ,_al_u7726_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~A*~(D*C*B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001010101010101),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6769|_al_u7873  (
    .a({open_n42661,\cu_ru/n84 [10]}),
    .b({open_n42662,_al_u6769_o}),
    .c({_al_u6765_o,_al_u7478_o}),
    .d({_al_u3399_o,\cu_ru/m_sip [5]}),
    .f({_al_u6769_o,_al_u7873_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6771|_al_u6774  (
    .c({_al_u6766_o,_al_u3397_o}),
    .d({_al_u6758_o,_al_u6766_o}),
    .f({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/read_mscratch_sel_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6772|cu_ru/m_s_scratch/reg1_b59  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n42711}),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/sepc [59]}),
    .c({\cu_ru/mcause [59],data_csr[59]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [59],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n42722,data_csr[59]}),
    .sr(rst_pad),
    .f({_al_u6772_o,_al_u5389_o}),
    .q({open_n42726,\cu_ru/sscratch [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6773|_al_u6770  (
    .c({_al_u6758_o,_al_u3397_o}),
    .d({_al_u6769_o,_al_u6769_o}),
    .f({\cu_ru/read_scause_sel_lutinv ,\cu_ru/read_sscratch_sel_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6775|cu_ru/m_s_cause/reg0_b59  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [59],\cu_ru/scause [59]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [59],data_csr[59]}),
    .sr(rst_pad),
    .f({_al_u6775_o,open_n42771}),
    .q({open_n42775,\cu_ru/scause [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6776|_al_u6783  (
    .c({_al_u6766_o,_al_u6769_o}),
    .d({_al_u3395_o,_al_u3395_o}),
    .f({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/read_sepc_sel_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(D*~C*B*A)"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"))
    \_al_u6778|_al_u6764  (
    .a({_al_u3393_o,_al_u3393_o}),
    .b({id_ins[22],id_ins[22]}),
    .c({id_ins[21],id_ins[21]}),
    .d({id_ins[20],id_ins[20]}),
    .f({_al_u6778_o,_al_u6764_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6779|_al_u6792  (
    .c({_al_u6778_o,_al_u6791_o}),
    .d({_al_u6777_o,_al_u6778_o}),
    .f({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_mtvec_sel_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u6780|cu_ru/m_s_cause/reg1_b59  (
    .a({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [59],\cu_ru/mepc [59]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [59],data_csr[59]}),
    .mi({open_n42851,data_csr[59]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6780_o,_al_u6588_o}),
    .q({open_n42866,\cu_ru/mcause [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6781|_al_u6835  (
    .b({_al_u6775_o,_al_u6833_o}),
    .c({_al_u6780_o,_al_u6834_o}),
    .d({_al_u6772_o,_al_u6832_o}),
    .f({_al_u6781_o,_al_u6835_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6784|cu_ru/m_s_epc/reg0_b59  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n42893}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({mtime_pad[59],_al_u5389_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [59],\cu_ru/m_s_epc/n2 [59]}),
    .sr(rst_pad),
    .f({_al_u6784_o,open_n42910}),
    .q({open_n42914,\cu_ru/sepc [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6785|cu_ru/m_cycle_event/reg0_b59  (
    .a({open_n42915,_al_u6763_o}),
    .b({_al_u6781_o,\cu_ru/read_mtval_sel_lutinv }),
    .c({_al_u6784_o,\cu_ru/minstret [59]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u6768_o,\cu_ru/mtval [59]}),
    .mi({open_n42919,\cu_ru/m_cycle_event/n4 [59]}),
    .sr(rst_pad),
    .f({_al_u6785_o,_al_u6768_o}),
    .q({open_n42934,\cu_ru/minstret [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6787|_al_u7339  (
    .b({open_n42937,\cu_ru/read_cycle_sel_lutinv }),
    .c({_al_u3397_o,\cu_ru/mcycle [6]}),
    .d({_al_u6761_o,\cu_ru/n82 [14]}),
    .f({\cu_ru/read_cycle_sel_lutinv ,_al_u7339_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6788|_al_u7269  (
    .a({open_n42962,\cu_ru/read_cycle_sel_lutinv }),
    .b({open_n42963,\cu_ru/read_sscratch_sel_lutinv }),
    .c({\cu_ru/read_cycle_sel_lutinv ,\cu_ru/mcycle [15]}),
    .d({\cu_ru/read_mcycle_sel_lutinv ,\cu_ru/sscratch [15]}),
    .f({_al_u6788_o,_al_u7269_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"))
    \_al_u6790|_al_u7725  (
    .a({_al_u6788_o,\cu_ru/read_stval_sel_lutinv }),
    .b({\cu_ru/read_stval_sel_lutinv ,\cu_ru/read_sepc_sel_lutinv }),
    .c({\cu_ru/mcycle [59],\cu_ru/sepc [0]}),
    .d({\cu_ru/stval [59],\cu_ru/stval [0]}),
    .f({_al_u6790_o,_al_u7725_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6794|cu_ru/m_s_epc/reg0_b58  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n43008}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [58],_al_u5393_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [58],\cu_ru/m_s_epc/n2 [58]}),
    .sr(rst_pad),
    .f({_al_u6794_o,open_n43025}),
    .q({open_n43029,\cu_ru/sepc [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6796|_al_u7231  (
    .a({_al_u6788_o,_al_u6788_o}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_mepc_sel_lutinv }),
    .c({\cu_ru/mcycle [58],\cu_ru/mcycle [34]}),
    .d({\cu_ru/stvec [58],\cu_ru/mepc [34]}),
    .f({_al_u6796_o,_al_u7231_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6797|cu_ru/m_s_cause/reg0_b58  (
    .a({\cu_ru/read_mcause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [58],\cu_ru/scause [58]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [58],data_csr[58]}),
    .sr(rst_pad),
    .f({_al_u6797_o,open_n43070}),
    .q({open_n43074,\cu_ru/scause [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6798|cu_ru/m_s_scratch/reg0_b58  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mscratch [58],\cu_ru/mtval [58]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [58],data_csr[58]}),
    .mi({open_n43085,data_csr[58]}),
    .sr(rst_pad),
    .f({_al_u6798_o,_al_u6461_o}),
    .q({open_n43089,\cu_ru/mscratch [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6799|cu_ru/m_s_tval/reg1_b58  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n43090}),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [58],\cu_ru/m_s_tval/n3 [58]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [58],_al_u6461_o}),
    .sr(rst_pad),
    .f({_al_u6799_o,open_n43104}),
    .q({open_n43108,\cu_ru/mtval [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6800|_al_u6993  (
    .b({_al_u6798_o,_al_u6991_o}),
    .c({_al_u6799_o,_al_u6992_o}),
    .d({_al_u6797_o,_al_u6990_o}),
    .f({_al_u6800_o,_al_u6993_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6801|cu_ru/m_s_tvec/reg1_b58  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,_al_u6795_o}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u6796_o}),
    .c({mtime_pad[58],_al_u6800_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [58],_al_u6801_o}),
    .sr(rst_pad),
    .f({_al_u6801_o,csr_data[58]}),
    .q({open_n43150,\cu_ru/mtvec [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6803|_al_u7082  (
    .a({_al_u6788_o,_al_u6788_o}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/mcycle [57],\cu_ru/mcycle [29]}),
    .d({\cu_ru/stvec [57],\cu_ru/stvec [29]}),
    .f({_al_u6803_o,_al_u7082_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6804|cu_ru/m_s_scratch/reg1_b57  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n43175}),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/sepc [57]}),
    .c({\cu_ru/mcause [57],data_csr[57]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [57],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n43179,data_csr[57]}),
    .sr(rst_pad),
    .f({_al_u6804_o,_al_u5397_o}),
    .q({open_n43194,\cu_ru/sscratch [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6805|cu_ru/m_s_cause/reg0_b57  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [57],\cu_ru/scause [57]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [57],data_csr[57]}),
    .sr(rst_pad),
    .f({_al_u6805_o,open_n43211}),
    .q({open_n43215,\cu_ru/scause [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6806|cu_ru/m_s_scratch/reg0_b57  (
    .a({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [57],\cu_ru/mtval [57]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [57],data_csr[57]}),
    .mi({open_n43226,data_csr[57]}),
    .sr(rst_pad),
    .f({_al_u6806_o,_al_u6463_o}),
    .q({open_n43230,\cu_ru/mscratch [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6807|_al_u6854  (
    .b({_al_u6805_o,_al_u6852_o}),
    .c({_al_u6806_o,_al_u6853_o}),
    .d({_al_u6804_o,_al_u6851_o}),
    .f({_al_u6807_o,_al_u6854_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6808|_al_u7288  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,\cu_ru/read_mtvec_sel_lutinv }),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/read_time_sel_lutinv }),
    .c({mtime_pad[57],mtime_pad[10]}),
    .d({\cu_ru/mtvec [57],\cu_ru/mtvec [10]}),
    .f({_al_u6808_o,_al_u7288_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6809|cu_ru/m_s_tvec/reg1_b57  (
    .a({open_n43277,_al_u6809_o}),
    .b({_al_u6807_o,_al_u6810_o}),
    .c({_al_u6808_o,\cu_ru/read_sepc_sel_lutinv }),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u6803_o,\cu_ru/sepc [57]}),
    .sr(rst_pad),
    .f({_al_u6809_o,csr_data[57]}),
    .q({open_n43297,\cu_ru/mtvec [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6813|cu_ru/m_s_epc/reg0_b56  (
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [56],_al_u5401_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u6812_o,\cu_ru/m_s_epc/n2 [56]}),
    .sr(rst_pad),
    .f({_al_u6813_o,open_n43316}),
    .q({open_n43320,\cu_ru/sepc [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6814|cu_ru/m_s_cause/reg0_b56  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/mcycle [56],\cu_ru/scause [56]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [56],data_csr[56]}),
    .sr(rst_pad),
    .f({_al_u6814_o,open_n43337}),
    .q({open_n43341,\cu_ru/scause [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6815|cu_ru/m_s_tval/reg1_b56  (
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [56],\cu_ru/m_s_tval/n3 [56]}),
    .clk(clk_pad),
    .d({_al_u6814_o,_al_u6465_o}),
    .sr(rst_pad),
    .f({_al_u6815_o,open_n43361}),
    .q({open_n43365,\cu_ru/mtval [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6816|cu_ru/m_s_scratch/reg0_b56  (
    .a({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcause [56],\cu_ru/mtval [56]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [56],data_csr[56]}),
    .mi({open_n43369,data_csr[56]}),
    .sr(rst_pad),
    .f({_al_u6816_o,_al_u6465_o}),
    .q({open_n43384,\cu_ru/mscratch [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6817|cu_ru/m_s_scratch/reg1_b56  (
    .a({\cu_ru/read_cycle_sel_lutinv ,open_n43385}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/sepc [56]}),
    .c({\cu_ru/mcycle [56],data_csr[56]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [56],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n43389,data_csr[56]}),
    .sr(rst_pad),
    .f({_al_u6817_o,_al_u5401_o}),
    .q({open_n43404,\cu_ru/sscratch [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6819|cu_ru/m_s_tvec/reg1_b56  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,_al_u6813_o}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u6818_o}),
    .c({\cu_ru/stvec [56],_al_u6819_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [56],_al_u6820_o}),
    .sr(rst_pad),
    .f({_al_u6819_o,csr_data[56]}),
    .q({open_n43424,\cu_ru/mtvec [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u6820|cu_ru/m_s_cause/reg1_b56  (
    .a({\cu_ru/read_time_sel_lutinv ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[56],\cu_ru/mepc [56]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [56],data_csr[56]}),
    .mi({open_n43435,data_csr[56]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6820_o,_al_u6594_o}),
    .q({open_n43439,\cu_ru/mcause [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6822|cu_ru/m_s_tval/reg1_b55  (
    .a({_al_u6788_o,open_n43440}),
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [55],\cu_ru/m_s_tval/n3 [55]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [55],_al_u6467_o}),
    .sr(rst_pad),
    .f({_al_u6822_o,open_n43458}),
    .q({open_n43462,\cu_ru/mtval [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6823|cu_ru/m_s_scratch/reg0_b55  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mscratch [55],\cu_ru/mtval [55]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [55],data_csr[55]}),
    .mi({open_n43466,data_csr[55]}),
    .sr(rst_pad),
    .f({_al_u6823_o,_al_u6467_o}),
    .q({open_n43481,\cu_ru/mscratch [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6824|cu_ru/m_s_cause/reg0_b55  (
    .a({\cu_ru/read_mcause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [55],\cu_ru/scause [55]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [55],data_csr[55]}),
    .sr(rst_pad),
    .f({_al_u6824_o,open_n43498}),
    .q({open_n43502,\cu_ru/scause [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u6825|cu_ru/m_s_cause/reg1_b55  (
    .a({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [55],\cu_ru/mepc [55]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [55],data_csr[55]}),
    .mi({open_n43506,data_csr[55]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6825_o,_al_u6596_o}),
    .q({open_n43521,\cu_ru/mcause [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6826|_al_u6828  (
    .b({_al_u6824_o,_al_u6826_o}),
    .c({_al_u6825_o,_al_u6827_o}),
    .d({_al_u6823_o,_al_u6822_o}),
    .f({_al_u6826_o,_al_u6828_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6827|cu_ru/m_s_epc/reg0_b55  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n43548}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({mtime_pad[55],_al_u5405_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [55],\cu_ru/m_s_epc/n2 [55]}),
    .sr(rst_pad),
    .f({_al_u6827_o,open_n43565}),
    .q({open_n43569,\cu_ru/sepc [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6831|cu_ru/m_s_cause/reg0_b54  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/mcycle [54],\cu_ru/scause [54]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [54],data_csr[54]}),
    .sr(rst_pad),
    .f({_al_u6831_o,open_n43586}),
    .q({open_n43590,\cu_ru/scause [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6832|cu_ru/m_s_tval/reg1_b54  (
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [54],\cu_ru/m_s_tval/n3 [54]}),
    .clk(clk_pad),
    .d({_al_u6831_o,_al_u6469_o}),
    .sr(rst_pad),
    .f({_al_u6832_o,open_n43606}),
    .q({open_n43610,\cu_ru/mtval [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6833|cu_ru/m_s_scratch/reg0_b54  (
    .a({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcause [54],\cu_ru/mtval [54]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [54],data_csr[54]}),
    .mi({open_n43621,data_csr[54]}),
    .sr(rst_pad),
    .f({_al_u6833_o,_al_u6469_o}),
    .q({open_n43625,\cu_ru/mscratch [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6834|cu_ru/m_s_scratch/reg1_b54  (
    .a({\cu_ru/read_cycle_sel_lutinv ,open_n43626}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/sepc [54]}),
    .c({\cu_ru/mcycle [54],data_csr[54]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [54],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n43637,data_csr[54]}),
    .sr(rst_pad),
    .f({_al_u6834_o,_al_u5409_o}),
    .q({open_n43641,\cu_ru/sscratch [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6837|cu_ru/m_s_epc/reg0_b54  (
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [54],_al_u5409_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u6836_o,\cu_ru/m_s_epc/n2 [54]}),
    .sr(rst_pad),
    .f({_al_u6837_o,open_n43660}),
    .q({open_n43664,\cu_ru/sepc [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6839|cu_ru/m_s_tvec/reg1_b54  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,_al_u6835_o}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u6837_o}),
    .c({\cu_ru/mepc [54],_al_u6838_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [54],_al_u6839_o}),
    .sr(rst_pad),
    .f({_al_u6839_o,csr_data[54]}),
    .q({open_n43684,\cu_ru/mtvec [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6842|cu_ru/m_cycle_event/reg0_b53  (
    .a({open_n43685,_al_u6763_o}),
    .b({\cu_ru/read_stval_sel_lutinv ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/stval [53],\cu_ru/minstret [53]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u6841_o,\cu_ru/stvec [53]}),
    .mi({open_n43689,\cu_ru/m_cycle_event/n4 [53]}),
    .sr(rst_pad),
    .f({_al_u6842_o,_al_u6841_o}),
    .q({open_n43704,\cu_ru/minstret [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6843|cu_ru/m_s_scratch/reg1_b53  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n43705}),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/sepc [53]}),
    .c({\cu_ru/mcause [53],data_csr[53]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [53],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n43709,data_csr[53]}),
    .sr(rst_pad),
    .f({_al_u6843_o,_al_u5413_o}),
    .q({open_n43724,\cu_ru/sscratch [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6845|cu_ru/m_s_cause/reg0_b53  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [53],\cu_ru/scause [53]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [53],data_csr[53]}),
    .sr(rst_pad),
    .f({_al_u6845_o,open_n43741}),
    .q({open_n43745,\cu_ru/scause [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6846|cu_ru/m_s_tvec/reg1_b53  (
    .a({_al_u6844_o,_al_u6842_o}),
    .b({_al_u6845_o,_al_u6846_o}),
    .c({\cu_ru/read_mtvec_sel_lutinv ,_al_u6847_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [53],_al_u6848_o}),
    .sr(rst_pad),
    .f({_al_u6846_o,csr_data[53]}),
    .q({open_n43761,\cu_ru/mtvec [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6847|cu_ru/m_s_epc/reg0_b53  (
    .a({\cu_ru/read_sepc_sel_lutinv ,open_n43762}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [53],_al_u5413_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [53],\cu_ru/m_s_epc/n2 [53]}),
    .sr(rst_pad),
    .f({_al_u6847_o,open_n43779}),
    .q({open_n43783,\cu_ru/sepc [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6848|cu_ru/m_s_scratch/reg0_b53  (
    .a({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[53],\cu_ru/mtval [53]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [53],data_csr[53]}),
    .mi({open_n43794,data_csr[53]}),
    .sr(rst_pad),
    .f({_al_u6848_o,_al_u6471_o}),
    .q({open_n43798,\cu_ru/mscratch [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6850|cu_ru/m_s_scratch/reg1_b52  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,open_n43799}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/sepc [52]}),
    .c({\cu_ru/mcycle [52],data_csr[52]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [52],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n43803,data_csr[52]}),
    .sr(rst_pad),
    .f({_al_u6850_o,_al_u5417_o}),
    .q({open_n43818,\cu_ru/sscratch [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6851|cu_ru/m_s_scratch/reg0_b52  (
    .a({open_n43819,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [52],\cu_ru/mtval [52]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({_al_u6850_o,data_csr[52]}),
    .mi({open_n43823,data_csr[52]}),
    .sr(rst_pad),
    .f({_al_u6851_o,_al_u6473_o}),
    .q({open_n43838,\cu_ru/mscratch [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6852|cu_ru/m_s_cause/reg0_b52  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [52],\cu_ru/scause [52]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [52],data_csr[52]}),
    .sr(rst_pad),
    .f({_al_u6852_o,open_n43855}),
    .q({open_n43859,\cu_ru/scause [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u6853|cu_ru/m_s_cause/reg1_b52  (
    .a({\cu_ru/read_cycle_sel_lutinv ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [52],\cu_ru/mepc [52]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [52],data_csr[52]}),
    .mi({open_n43870,data_csr[52]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6853_o,_al_u6602_o}),
    .q({open_n43874,\cu_ru/mcause [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6855|cu_ru/m_s_epc/reg0_b52  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n43875}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({mtime_pad[52],_al_u5417_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [52],\cu_ru/m_s_epc/n2 [52]}),
    .sr(rst_pad),
    .f({_al_u6855_o,open_n43892}),
    .q({open_n43896,\cu_ru/sepc [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u6856|_al_u6866  (
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/read_mepc_sel_lutinv }),
    .c(\cu_ru/mepc [52:51]),
    .d({_al_u6855_o,_al_u6865_o}),
    .f({_al_u6856_o,_al_u6866_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6858|cu_ru/m_s_tvec/reg1_b52  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,_al_u6854_o}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u6856_o}),
    .c({\cu_ru/stval [52],_al_u6857_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [52],_al_u6858_o}),
    .sr(rst_pad),
    .f({_al_u6858_o,csr_data[52]}),
    .q({open_n43934,\cu_ru/mtvec [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6860|cu_ru/m_s_scratch/reg1_b51  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,open_n43935}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/sepc [51]}),
    .c({\cu_ru/mcycle [51],data_csr[51]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [51],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n43946,data_csr[51]}),
    .sr(rst_pad),
    .f({_al_u6860_o,_al_u5421_o}),
    .q({open_n43950,\cu_ru/sscratch [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6861|cu_ru/m_s_scratch/reg0_b51  (
    .a({open_n43951,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [51],\cu_ru/mtval [51]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({_al_u6860_o,data_csr[51]}),
    .mi({open_n43955,data_csr[51]}),
    .sr(rst_pad),
    .f({_al_u6861_o,_al_u6475_o}),
    .q({open_n43970,\cu_ru/mscratch [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6862|cu_ru/m_s_cause/reg0_b51  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [51],\cu_ru/scause [51]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [51],data_csr[51]}),
    .sr(rst_pad),
    .f({_al_u6862_o,open_n43987}),
    .q({open_n43991,\cu_ru/scause [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u6863|cu_ru/m_s_cause/reg1_b51  (
    .a({\cu_ru/read_cycle_sel_lutinv ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [51],\cu_ru/mepc [51]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [51],data_csr[51]}),
    .mi({open_n43995,data_csr[51]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6863_o,_al_u6604_o}),
    .q({open_n44010,\cu_ru/mcause [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6864|_al_u6914  (
    .b({_al_u6862_o,_al_u6912_o}),
    .c({_al_u6863_o,_al_u6913_o}),
    .d({_al_u6861_o,_al_u6911_o}),
    .f({_al_u6864_o,_al_u6914_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6865|cu_ru/m_s_epc/reg0_b51  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n44037}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({mtime_pad[51],_al_u5421_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [51],\cu_ru/m_s_epc/n2 [51]}),
    .sr(rst_pad),
    .f({_al_u6865_o,open_n44054}),
    .q({open_n44058,\cu_ru/sepc [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6868|cu_ru/m_s_tvec/reg1_b51  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,_al_u6864_o}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u6866_o}),
    .c({\cu_ru/stval [51],_al_u6867_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [51],_al_u6868_o}),
    .sr(rst_pad),
    .f({_al_u6868_o,csr_data[51]}),
    .q({open_n44078,\cu_ru/mtvec [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6871|cu_ru/m_s_tvec/reg1_b50  (
    .a({open_n44079,_al_u6871_o}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u6876_o}),
    .c({mtime_pad[50],_al_u6877_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u6870_o,_al_u6878_o}),
    .sr(rst_pad),
    .f({_al_u6871_o,csr_data[50]}),
    .q({open_n44099,\cu_ru/mtvec [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6872|cu_ru/m_s_cause/reg0_b50  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [50],\cu_ru/scause [50]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [50],data_csr[50]}),
    .sr(rst_pad),
    .f({_al_u6872_o,open_n44116}),
    .q({open_n44120,\cu_ru/scause [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u6874|cu_ru/m_s_cause/reg1_b50  (
    .a({\cu_ru/read_cycle_sel_lutinv ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [50],\cu_ru/mepc [50]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [50],data_csr[50]}),
    .mi({open_n44124,data_csr[50]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6874_o,_al_u6606_o}),
    .q({open_n44139,\cu_ru/mcause [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6875|cu_ru/m_s_scratch/reg1_b50  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,open_n44140}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/sepc [50]}),
    .c({\cu_ru/mcycle [50],data_csr[50]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [50],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n44151,data_csr[50]}),
    .sr(rst_pad),
    .f({_al_u6875_o,_al_u5425_o}),
    .q({open_n44155,\cu_ru/sscratch [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6876|_al_u6873  (
    .b({_al_u6874_o,\cu_ru/read_mtvec_sel_lutinv }),
    .c({_al_u6875_o,\cu_ru/mtvec [50]}),
    .d({_al_u6873_o,_al_u6872_o}),
    .f({_al_u6876_o,_al_u6873_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6877|cu_ru/m_s_epc/reg0_b50  (
    .a({\cu_ru/read_sepc_sel_lutinv ,open_n44182}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [50],_al_u5425_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [50],\cu_ru/m_s_epc/n2 [50]}),
    .sr(rst_pad),
    .f({_al_u6877_o,open_n44199}),
    .q({open_n44203,\cu_ru/sepc [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6878|cu_ru/m_s_scratch/reg0_b50  (
    .a({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [50],\cu_ru/mtval [50]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [50],data_csr[50]}),
    .mi({open_n44214,data_csr[50]}),
    .sr(rst_pad),
    .f({_al_u6878_o,_al_u6477_o}),
    .q({open_n44218,\cu_ru/mscratch [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6881|cu_ru/m_cycle_event/reg0_b49  (
    .a({open_n44219,_al_u6763_o}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/read_sepc_sel_lutinv }),
    .c({mtime_pad[49],\cu_ru/minstret [49]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u6880_o,\cu_ru/sepc [49]}),
    .mi({open_n44230,\cu_ru/m_cycle_event/n4 [49]}),
    .sr(rst_pad),
    .f({_al_u6881_o,_al_u6880_o}),
    .q({open_n44234,\cu_ru/minstret [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6882|cu_ru/m_s_cause/reg0_b49  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [49],\cu_ru/scause [49]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [49],data_csr[49]}),
    .sr(rst_pad),
    .f({_al_u6882_o,open_n44251}),
    .q({open_n44255,\cu_ru/scause [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6883|_al_u6836  (
    .a({open_n44256,\cu_ru/read_stval_sel_lutinv }),
    .b({\cu_ru/read_stval_sel_lutinv ,\cu_ru/read_time_sel_lutinv }),
    .c({\cu_ru/stval [49],mtime_pad[54]}),
    .d({_al_u6882_o,\cu_ru/stval [54]}),
    .f({_al_u6883_o,_al_u6836_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u6884|cu_ru/m_s_cause/reg1_b49  (
    .a({\cu_ru/read_cycle_sel_lutinv ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [49],\cu_ru/mepc [49]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [49],data_csr[49]}),
    .mi({open_n44291,data_csr[49]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6884_o,_al_u6610_o}),
    .q({open_n44295,\cu_ru/mcause [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6885|cu_ru/m_s_scratch/reg1_b49  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,open_n44296}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/sepc [49]}),
    .c({\cu_ru/mcycle [49],data_csr[49]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [49],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n44300,data_csr[49]}),
    .sr(rst_pad),
    .f({_al_u6885_o,_al_u5433_o}),
    .q({open_n44315,\cu_ru/sscratch [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6886|cu_ru/m_s_tvec/reg1_b49  (
    .a({open_n44316,_al_u6881_o}),
    .b({_al_u6884_o,_al_u6886_o}),
    .c({_al_u6885_o,_al_u6887_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u6883_o,_al_u6888_o}),
    .sr(rst_pad),
    .f({_al_u6886_o,csr_data[49]}),
    .q({open_n44332,\cu_ru/mtvec [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6888|cu_ru/m_s_scratch/reg0_b49  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [49],\cu_ru/mtval [49]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [49],data_csr[49]}),
    .mi({open_n44343,data_csr[49]}),
    .sr(rst_pad),
    .f({_al_u6888_o,_al_u6481_o}),
    .q({open_n44347,\cu_ru/mscratch [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6890|_al_u7072  (
    .a({_al_u6788_o,_al_u6788_o}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_mtvec_sel_lutinv }),
    .c({\cu_ru/mcycle [48],\cu_ru/mcycle [31]}),
    .d({\cu_ru/stvec [48],\cu_ru/mtvec [31]}),
    .f({_al_u6890_o,_al_u7072_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6891|cu_ru/m_s_scratch/reg1_b48  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n44372}),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/sepc [48]}),
    .c({\cu_ru/mcause [48],data_csr[48]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [48],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n44376,data_csr[48]}),
    .sr(rst_pad),
    .f({_al_u6891_o,_al_u5437_o}),
    .q({open_n44391,\cu_ru/sscratch [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6892|cu_ru/m_s_cause/reg0_b48  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [48],\cu_ru/scause [48]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [48],data_csr[48]}),
    .sr(rst_pad),
    .f({_al_u6892_o,open_n44408}),
    .q({open_n44412,\cu_ru/scause [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6893|cu_ru/m_s_scratch/reg0_b48  (
    .a({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [48],\cu_ru/mtval [48]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [48],data_csr[48]}),
    .mi({open_n44416,data_csr[48]}),
    .sr(rst_pad),
    .f({_al_u6893_o,_al_u6483_o}),
    .q({open_n44431,\cu_ru/mscratch [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6894|_al_u6896  (
    .b({_al_u6892_o,_al_u6894_o}),
    .c({_al_u6893_o,_al_u6895_o}),
    .d({_al_u6891_o,_al_u6890_o}),
    .f({_al_u6894_o,_al_u6896_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6895|cu_ru/m_s_epc/reg0_b48  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n44454}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({mtime_pad[48],_al_u5437_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [48],\cu_ru/m_s_epc/n2 [48]}),
    .sr(rst_pad),
    .f({_al_u6895_o,open_n44471}),
    .q({open_n44475,\cu_ru/sepc [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6900|cu_ru/m_s_scratch/reg1_b47  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n44476}),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/sepc [47]}),
    .c({\cu_ru/mcause [47],data_csr[47]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [47],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n44487,data_csr[47]}),
    .sr(rst_pad),
    .f({_al_u6900_o,_al_u5441_o}),
    .q({open_n44491,\cu_ru/sscratch [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6901|cu_ru/m_s_cause/reg0_b47  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [47],\cu_ru/scause [47]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [47],data_csr[47]}),
    .sr(rst_pad),
    .f({_al_u6901_o,open_n44508}),
    .q({open_n44512,\cu_ru/scause [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u6902|cu_ru/m_s_cause/reg1_b47  (
    .a({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [47],\cu_ru/mepc [47]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [47],data_csr[47]}),
    .mi({open_n44516,data_csr[47]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6902_o,_al_u6614_o}),
    .q({open_n44531,\cu_ru/mcause [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6903|_al_u7105  (
    .b({_al_u6901_o,_al_u7103_o}),
    .c({_al_u6902_o,_al_u7104_o}),
    .d({_al_u6900_o,_al_u7102_o}),
    .f({_al_u6903_o,_al_u7105_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u6904|_al_u6971  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,\cu_ru/read_mtvec_sel_lutinv }),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/read_time_sel_lutinv }),
    .c({mtime_pad[47],mtime_pad[61]}),
    .d({\cu_ru/mtvec [47],\cu_ru/mtvec [61]}),
    .f({_al_u6904_o,_al_u6971_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6905|cu_ru/m_cycle_event/reg0_b47  (
    .a({open_n44574,_al_u6763_o}),
    .b({_al_u6903_o,\cu_ru/read_mtval_sel_lutinv }),
    .c({_al_u6904_o,\cu_ru/minstret [47]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u6899_o,\cu_ru/mtval [47]}),
    .mi({open_n44578,\cu_ru/m_cycle_event/n4 [47]}),
    .sr(rst_pad),
    .f({_al_u6905_o,_al_u6899_o}),
    .q({open_n44593,\cu_ru/minstret [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*A*~(D*C))"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("~(B*A*~(D*C))"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111011101110111),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b1111011101110111),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6906|cu_ru/m_s_tvec/reg1_b47  (
    .a({_al_u6788_o,_al_u6905_o}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u6906_o}),
    .c({\cu_ru/mcycle [47],\cu_ru/read_sepc_sel_lutinv }),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/stval [47],\cu_ru/sepc [47]}),
    .sr(rst_pad),
    .f({_al_u6906_o,csr_data[47]}),
    .q({open_n44613,\cu_ru/mtvec [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6908|cu_ru/m_s_epc/reg0_b46  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n44614}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [46],_al_u5445_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [46],\cu_ru/m_s_epc/n2 [46]}),
    .sr(rst_pad),
    .f({_al_u6908_o,open_n44631}),
    .q({open_n44635,\cu_ru/sepc [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6909|_al_u6981  (
    .a({open_n44636,_al_u6788_o}),
    .b({_al_u6908_o,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/mcycle [46],\cu_ru/mcycle [60]}),
    .d({_al_u6788_o,\cu_ru/stvec [60]}),
    .f({_al_u6909_o,_al_u6981_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6911|cu_ru/m_s_cause/reg0_b46  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [46],\cu_ru/scause [46]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [46],data_csr[46]}),
    .sr(rst_pad),
    .f({_al_u6911_o,open_n44677}),
    .q({open_n44681,\cu_ru/scause [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6912|cu_ru/m_s_scratch/reg1_b46  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n44682}),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/sepc [46]}),
    .c({\cu_ru/mcause [46],data_csr[46]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [46],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n44693,data_csr[46]}),
    .sr(rst_pad),
    .f({_al_u6912_o,_al_u5445_o}),
    .q({open_n44697,\cu_ru/sscratch [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6913|cu_ru/m_s_scratch/reg0_b46  (
    .a({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [46],\cu_ru/mtval [46]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [46],data_csr[46]}),
    .mi({open_n44708,data_csr[46]}),
    .sr(rst_pad),
    .f({_al_u6913_o,_al_u6487_o}),
    .q({open_n44712,\cu_ru/mscratch [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6915|cu_ru/m_s_tvec/reg1_b46  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,_al_u6909_o}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u6910_o}),
    .c({mtime_pad[46],_al_u6914_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [46],_al_u6915_o}),
    .sr(rst_pad),
    .f({_al_u6915_o,csr_data[46]}),
    .q({open_n44732,\cu_ru/mtvec [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6917|cu_ru/m_s_epc/reg0_b45  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n44733}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [45],_al_u5449_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [45],\cu_ru/m_s_epc/n2 [45]}),
    .sr(rst_pad),
    .f({_al_u6917_o,open_n44750}),
    .q({open_n44754,\cu_ru/sepc [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u6918|_al_u6948  (
    .b({_al_u6917_o,\cu_ru/read_stval_sel_lutinv }),
    .c({\cu_ru/mcycle [45],\cu_ru/stval [63]}),
    .d({_al_u6788_o,_al_u6947_o}),
    .f({_al_u6918_o,_al_u6948_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6920|cu_ru/m_s_cause/reg0_b45  (
    .a({\cu_ru/read_mcause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [45],\cu_ru/scause [45]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [45],data_csr[45]}),
    .sr(rst_pad),
    .f({_al_u6920_o,open_n44793}),
    .q({open_n44797,\cu_ru/scause [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6921|cu_ru/m_s_scratch/reg0_b45  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mscratch [45],\cu_ru/mtval [45]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [45],data_csr[45]}),
    .mi({open_n44808,data_csr[45]}),
    .sr(rst_pad),
    .f({_al_u6921_o,_al_u6489_o}),
    .q({open_n44812,\cu_ru/mscratch [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6923|_al_u6922  (
    .a({open_n44813,\cu_ru/read_mepc_sel_lutinv }),
    .b({_al_u6921_o,\cu_ru/read_stvec_sel_lutinv }),
    .c({_al_u6922_o,\cu_ru/mepc [45]}),
    .d({_al_u6920_o,\cu_ru/stvec [45]}),
    .f({_al_u6923_o,_al_u6922_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6924|cu_ru/m_s_tvec/reg1_b45  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,_al_u6918_o}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u6919_o}),
    .c({mtime_pad[45],_al_u6923_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [45],_al_u6924_o}),
    .sr(rst_pad),
    .f({_al_u6924_o,csr_data[45]}),
    .q({open_n44853,\cu_ru/mtvec [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6926|cu_ru/m_s_epc/reg0_b44  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n44854}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [44],_al_u5453_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [44],\cu_ru/m_s_epc/n2 [44]}),
    .sr(rst_pad),
    .f({_al_u6926_o,open_n44871}),
    .q({open_n44875,\cu_ru/sepc [44]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"))
    \_al_u6928|_al_u7052  (
    .a({_al_u6788_o,_al_u6788_o}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/mcycle [44],\cu_ru/mcycle [37]}),
    .d({\cu_ru/stvec [44],\cu_ru/stvec [37]}),
    .f({_al_u6928_o,_al_u7052_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6929|cu_ru/m_s_cause/reg0_b44  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [44],\cu_ru/scause [44]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [44],data_csr[44]}),
    .sr(rst_pad),
    .f({_al_u6929_o,open_n44912}),
    .q({open_n44916,\cu_ru/scause [44]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6930|cu_ru/m_s_scratch/reg1_b44  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n44917}),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/sepc [44]}),
    .c({\cu_ru/mcause [44],data_csr[44]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [44],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n44921,data_csr[44]}),
    .sr(rst_pad),
    .f({_al_u6930_o,_al_u5453_o}),
    .q({open_n44936,\cu_ru/sscratch [44]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6931|cu_ru/m_s_tval/reg1_b44  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n44937}),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [44],\cu_ru/m_s_tval/n3 [44]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [44],_al_u6491_o}),
    .sr(rst_pad),
    .f({_al_u6931_o,open_n44955}),
    .q({open_n44959,\cu_ru/mtval [44]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6932|_al_u7230  (
    .b({_al_u6930_o,_al_u7228_o}),
    .c({_al_u6931_o,_al_u7229_o}),
    .d({_al_u6929_o,_al_u7227_o}),
    .f({_al_u6932_o,_al_u7230_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6933|cu_ru/m_s_tvec/reg1_b44  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,_al_u6927_o}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u6928_o}),
    .c({mtime_pad[44],_al_u6932_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [44],_al_u6933_o}),
    .sr(rst_pad),
    .f({_al_u6933_o,csr_data[44]}),
    .q({open_n45001,\cu_ru/mtvec [44]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~((~C*~A))*~(B)+~D*(~C*~A)*~(B)+~(~D)*(~C*~A)*B+~D*(~C*~A)*B)"),
    //.LUTF1("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("~(~D*~((~C*~A))*~(B)+~D*(~C*~A)*~(B)+~(~D)*(~C*~A)*B+~D*(~C*~A)*B)"),
    //.LUTG1("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101111001000),
    .INIT_LUTF1(16'b0011000100100000),
    .INIT_LUTG0(16'b1111101111001000),
    .INIT_LUTG1(16'b0011000100100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6935|cu_ru/m_s_status/spp_reg  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6935_o}),
    .b({_al_u2842_o,\cu_ru/m_s_status/u34_sel_is_0_o }),
    .c({priv[1],_al_u6936_o}),
    .clk(clk_pad),
    .d({\cu_ru/mstatus [8],data_csr[8]}),
    .sr(rst_pad),
    .f({_al_u6935_o,open_n45019}),
    .q({open_n45023,\cu_ru/mstatus [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0001010110111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6938|_al_u9622  (
    .a({open_n45024,\cu_ru/m_s_status/n2 }),
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/mstatus [5],\cu_ru/sepc [19]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/mepc [19]}),
    .f({_al_u6938_o,_al_u9622_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B)"),
    //.LUTF1("(B*~(D*~C*~A))"),
    //.LUTG0("(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B)"),
    //.LUTG1("(B*~(D*~C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011011100000100),
    .INIT_LUTF1(16'b1100100011001100),
    .INIT_LUTG0(16'b0011011100000100),
    .INIT_LUTG1(16'b1100100011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6939|cu_ru/m_s_status/sie_reg  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6939_o}),
    .b({_al_u6938_o,\cu_ru/m_s_status/u34_sel_is_0_o }),
    .c({_al_u2844_o,_al_u6940_o}),
    .clk(clk_pad),
    .d({\cu_ru/mstatus [1],data_csr[1]}),
    .sr(rst_pad),
    .f({_al_u6939_o,open_n45066}),
    .q({open_n45070,\cu_ru/mstatus [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~((~C*~A))*~(B)+~D*(~C*~A)*~(B)+~(~D)*(~C*~A)*B+~D*(~C*~A)*B)"),
    //.LUT1("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111101111001000),
    .INIT_LUT1(16'b0011000100100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6942|cu_ru/m_s_status/spie_reg  (
    .a({\cu_ru/m_s_status/u14_sel_is_2_o ,_al_u6942_o}),
    .b({_al_u2842_o,\cu_ru/m_s_status/u34_sel_is_0_o }),
    .c({\cu_ru/mstatus [1],_al_u6943_o}),
    .clk(clk_pad),
    .d({\cu_ru/mstatus [5],data_csr[5]}),
    .sr(rst_pad),
    .f({_al_u6942_o,open_n45084}),
    .q({open_n45088,\cu_ru/mstatus [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u6943|_al_u6936  (
    .c({\cu_ru/mstatus [5],\cu_ru/mstatus [8]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u6943_o,_al_u6936_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u6945|_al_u6946  (
    .b({id_ins[27],_al_u3399_o}),
    .c({id_ins[26],_al_u6945_o}),
    .d({id_ins[28],_al_u3397_o}),
    .f({_al_u6945_o,\cu_ru/read_satp_sel_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6947|cu_ru/m_s_scratch/reg1_b63  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({satp[63],\cu_ru/mtval [63]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [63],data_csr[63]}),
    .mi({open_n45145,data_csr[63]}),
    .sr(rst_pad),
    .f({_al_u6947_o,_al_u6449_o}),
    .q({open_n45149,\cu_ru/sscratch [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6949|cu_ru/csr_satp/reg1_b3  (
    .a({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/m_s_cause/mux4_b0_sel_is_2_o }),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/scause [63],\cu_ru/mcause [63]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [63],data_csr[63]}),
    .mi({open_n45160,data_csr[63]}),
    .sr(rst_pad),
    .f({_al_u6949_o,_al_u6698_o}),
    .q({open_n45164,satp[63]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6950|cu_ru/m_s_scratch/reg0_b63  (
    .a({_al_u6948_o,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u6949_o,\cu_ru/trap_target_m }),
    .c({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/mepc [63]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [63],data_csr[63]}),
    .mi({open_n45175,data_csr[63]}),
    .sr(rst_pad),
    .f({_al_u6950_o,_al_u6578_o}),
    .q({open_n45179,\cu_ru/mscratch [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6952|cu_ru/m_s_tval/reg1_b63  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n45180}),
    .b({\cu_ru/read_sepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/sepc [63],\cu_ru/m_s_tval/n3 [63]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [63],_al_u6449_o}),
    .sr(rst_pad),
    .f({_al_u6952_o,open_n45198}),
    .q({open_n45202,\cu_ru/mtval [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u6953|_al_u6951  (
    .a({open_n45203,\cu_ru/read_mtvec_sel_lutinv }),
    .b({_al_u6951_o,\cu_ru/read_time_sel_lutinv }),
    .c({_al_u6952_o,mtime_pad[63]}),
    .d({_al_u6950_o,\cu_ru/mtvec [63]}),
    .f({_al_u6953_o,_al_u6951_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6955|cu_ru/m_s_tvec/reg1_b63  (
    .a({\cu_ru/read_mepc_sel_lutinv ,open_n45224}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u6954_o}),
    .c({\cu_ru/mepc [63],_al_u6955_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [63],_al_u6953_o}),
    .sr(rst_pad),
    .f({_al_u6955_o,csr_data[63]}),
    .q({open_n45244,\cu_ru/mtvec [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6957|cu_ru/m_s_scratch/reg1_b62  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n45245}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/stval [62]}),
    .c({satp[62],data_csr[62]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [62],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n45249,data_csr[62]}),
    .sr(rst_pad),
    .f({_al_u6957_o,_al_u5173_o}),
    .q({open_n45264,\cu_ru/sscratch [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6959|cu_ru/m_s_cause/reg0_b62  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [62],\cu_ru/scause [62]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [62],data_csr[62]}),
    .sr(rst_pad),
    .f({_al_u6959_o,open_n45281}),
    .q({open_n45285,\cu_ru/scause [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6960|cu_ru/m_cycle_event/reg0_b62  (
    .a({_al_u6958_o,open_n45286}),
    .b({_al_u6959_o,_al_u6957_o}),
    .c({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/minstret [62]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [62],_al_u6763_o}),
    .mi({open_n45297,\cu_ru/m_cycle_event/n4 [62]}),
    .sr(rst_pad),
    .f({_al_u6960_o,_al_u6958_o}),
    .q({open_n45301,\cu_ru/minstret [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"))
    \_al_u6961|_al_u7022  (
    .a({_al_u6788_o,_al_u6788_o}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/mcycle [62],\cu_ru/mcycle [40]}),
    .d({\cu_ru/stvec [62],\cu_ru/stvec [40]}),
    .f({_al_u6961_o,_al_u7022_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6962|cu_ru/m_s_tval/reg1_b62  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n45322}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[62],\cu_ru/m_s_tval/n3 [62]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [62],_al_u6451_o}),
    .sr(rst_pad),
    .f({_al_u6962_o,open_n45340}),
    .q({open_n45344,\cu_ru/mtval [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6963|cu_ru/m_s_tvec/reg1_b62  (
    .b({_al_u6961_o,_al_u6964_o}),
    .c({_al_u6962_o,_al_u6965_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u6960_o,_al_u6963_o}),
    .sr(rst_pad),
    .f({_al_u6963_o,csr_data[62]}),
    .q({open_n45366,\cu_ru/mtvec [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6964|cu_ru/m_s_tval/reg0_b62  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n45367}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5173_o}),
    .c({\cu_ru/mepc [62],\cu_ru/m_s_tval/n3 [62]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [62],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u6964_o,open_n45384}),
    .q({open_n45388,\cu_ru/stval [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6965|cu_ru/m_s_epc/reg0_b62  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n45389}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [62],_al_u5373_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [62],\cu_ru/m_s_epc/n2 [62]}),
    .sr(rst_pad),
    .f({_al_u6965_o,open_n45406}),
    .q({open_n45410,\cu_ru/sepc [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6967|cu_ru/csr_satp/reg1_b1  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({satp[61],\cu_ru/mepc [61]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [61],data_csr[61]}),
    .mi({open_n45414,data_csr[61]}),
    .sr(rst_pad),
    .f({_al_u6967_o,_al_u6582_o}),
    .q({open_n45429,satp[61]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6968|cu_ru/m_s_tval/reg0_b61  (
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5176_o}),
    .c({\cu_ru/stval [61],\cu_ru/m_s_tval/n3 [61]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u6967_o,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u6968_o,open_n45448}),
    .q({open_n45452,\cu_ru/stval [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6969|cu_ru/m_s_cause/reg0_b61  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [61],\cu_ru/scause [61]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [61],data_csr[61]}),
    .sr(rst_pad),
    .f({_al_u6969_o,open_n45469}),
    .q({open_n45473,\cu_ru/scause [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u6970|cu_ru/m_s_cause/reg1_b61  (
    .a({_al_u6968_o,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({_al_u6969_o,\cu_ru/trap_target_m }),
    .c({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/mtval [61]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [61],data_csr[61]}),
    .mi({open_n45484,data_csr[61]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6970_o,_al_u6453_o}),
    .q({open_n45488,\cu_ru/mcause [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6972|cu_ru/m_s_tval/reg1_b61  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n45489}),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [61],\cu_ru/m_s_tval/n3 [61]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [61],_al_u6453_o}),
    .sr(rst_pad),
    .f({_al_u6972_o,open_n45503}),
    .q({open_n45507,\cu_ru/mtval [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6973|cu_ru/m_s_tvec/reg1_b61  (
    .b({_al_u6971_o,_al_u6974_o}),
    .c({_al_u6972_o,_al_u6975_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u6970_o,_al_u6973_o}),
    .sr(rst_pad),
    .f({_al_u6973_o,csr_data[61]}),
    .q({open_n45525,\cu_ru/mtvec [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6975|cu_ru/m_s_epc/reg0_b61  (
    .a({_al_u6788_o,open_n45526}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/mcycle [61],_al_u5377_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [61],\cu_ru/m_s_epc/n2 [61]}),
    .sr(rst_pad),
    .f({_al_u6975_o,open_n45543}),
    .q({open_n45547,\cu_ru/sepc [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6977|cu_ru/csr_satp/reg1_b0  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({satp[60],\cu_ru/mepc [60]}),
    .ce(\cu_ru/csr_satp/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [60],data_csr[60]}),
    .mi({open_n45558,data_csr[60]}),
    .sr(rst_pad),
    .f({_al_u6977_o,_al_u6584_o}),
    .q({open_n45562,satp[60]}));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6979|cu_ru/m_s_cause/reg0_b60  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [60],\cu_ru/scause [60]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [60],data_csr[60]}),
    .sr(rst_pad),
    .f({_al_u6979_o,open_n45579}),
    .q({open_n45583,\cu_ru/scause [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6980|cu_ru/m_cycle_event/reg0_b60  (
    .a({_al_u6978_o,open_n45584}),
    .b({_al_u6979_o,_al_u6977_o}),
    .c({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/minstret [60]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [60],_al_u6763_o}),
    .mi({open_n45588,\cu_ru/m_cycle_event/n4 [60]}),
    .sr(rst_pad),
    .f({_al_u6980_o,_al_u6978_o}),
    .q({open_n45603,\cu_ru/minstret [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6982|cu_ru/m_s_tval/reg1_b60  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n45604}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[60],\cu_ru/m_s_tval/n3 [60]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [60],_al_u6455_o}),
    .sr(rst_pad),
    .f({_al_u6982_o,open_n45618}),
    .q({open_n45622,\cu_ru/mtval [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6983|cu_ru/m_s_tvec/reg1_b60  (
    .b({_al_u6981_o,_al_u6984_o}),
    .c({_al_u6982_o,_al_u6985_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u6980_o,_al_u6983_o}),
    .sr(rst_pad),
    .f({_al_u6983_o,csr_data[60]}),
    .q({open_n45640,\cu_ru/mtvec [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6984|cu_ru/m_s_tval/reg0_b60  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n45641}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5179_o}),
    .c({\cu_ru/mepc [60],\cu_ru/m_s_tval/n3 [60]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [60],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u6984_o,open_n45654}),
    .q({open_n45658,\cu_ru/stval [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6985|cu_ru/m_s_epc/reg0_b60  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n45659}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [60],_al_u5381_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [60],\cu_ru/m_s_epc/n2 [60]}),
    .sr(rst_pad),
    .f({_al_u6985_o,open_n45676}),
    .q({open_n45680,\cu_ru/sepc [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6987|cu_ru/m_s_cause/reg0_b43  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [43],\cu_ru/scause [43]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [43],data_csr[43]}),
    .sr(rst_pad),
    .f({_al_u6987_o,open_n45697}),
    .q({open_n45701,\cu_ru/scause [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6988|cu_ru/m_s_epc/reg0_b43  (
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [43],_al_u5457_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u6987_o,\cu_ru/m_s_epc/n2 [43]}),
    .sr(rst_pad),
    .f({_al_u6988_o,open_n45720}),
    .q({open_n45724,\cu_ru/sepc [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6989|cu_ru/m_s_scratch/reg1_b43  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n45725}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/stval [43]}),
    .c({satp[43],data_csr[43]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [43],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n45729,data_csr[43]}),
    .sr(rst_pad),
    .f({_al_u6989_o,_al_u5236_o}),
    .q({open_n45744,\cu_ru/sscratch [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u6990|cu_ru/m_s_cause/reg1_b43  (
    .a({_al_u6988_o,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({_al_u6989_o,\cu_ru/trap_target_m }),
    .c({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/mtval [43]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [43],data_csr[43]}),
    .mi({open_n45748,data_csr[43]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6990_o,_al_u6493_o}),
    .q({open_n45763,\cu_ru/mcause [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6991|_al_u6020  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/stvec [43],\cu_ru/stvec [43]}),
    .d({\cu_ru/mtvec [43],\cu_ru/mtvec [43]}),
    .f({_al_u6991_o,\cu_ru/tvec [43]}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6992|cu_ru/m_s_tval/reg0_b43  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n45788}),
    .b({\cu_ru/read_mtval_sel_lutinv ,_al_u5236_o}),
    .c({\cu_ru/stval [43],\cu_ru/m_s_tval/n3 [43]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [43],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u6992_o,open_n45805}),
    .q({open_n45809,\cu_ru/stval [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6995|cu_ru/m_s_tvec/reg1_b43  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n45810}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u6994_o}),
    .c({mtime_pad[43],_al_u6995_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [43],_al_u6993_o}),
    .sr(rst_pad),
    .f({_al_u6995_o,csr_data[43]}),
    .q({open_n45830,\cu_ru/mtvec [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u6997|cu_ru/m_s_cause/reg0_b42  (
    .a({\cu_ru/read_mcause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [42],\cu_ru/scause [42]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [42],data_csr[42]}),
    .sr(rst_pad),
    .f({_al_u6997_o,open_n45847}),
    .q({open_n45851,\cu_ru/scause [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u6998|_al_u7251  (
    .a({open_n45852,\cu_ru/read_cycle_sel_lutinv }),
    .b({\cu_ru/read_instret_sel_lutinv ,\cu_ru/read_instret_sel_lutinv }),
    .c({\cu_ru/minstret [42],\cu_ru/minstret [21]}),
    .d({_al_u6997_o,\cu_ru/mcycle [21]}),
    .f({_al_u6998_o,_al_u7251_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7000|cu_ru/m_s_scratch/reg0_b42  (
    .a({\cu_ru/read_mscratch_sel_lutinv ,open_n45877}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/sepc [42]}),
    .c({satp[42],data_csr[42]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [42],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n45888,data_csr[42]}),
    .sr(rst_pad),
    .f({_al_u7000_o,_al_u5461_o}),
    .q({open_n45892,\cu_ru/mscratch [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7001|cu_ru/m_cycle_event/reg0_b42  (
    .a({open_n45893,\cu_ru/read_minstret_sel_lutinv }),
    .b({_al_u6999_o,\cu_ru/read_sscratch_sel_lutinv }),
    .c({_al_u7000_o,\cu_ru/minstret [42]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u6998_o,\cu_ru/sscratch [42]}),
    .mi({open_n45904,\cu_ru/m_cycle_event/n4 [42]}),
    .sr(rst_pad),
    .f({_al_u7001_o,_al_u6999_o}),
    .q({open_n45908,\cu_ru/minstret [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7002|cu_ru/m_s_epc/reg0_b42  (
    .a({\cu_ru/read_sepc_sel_lutinv ,open_n45909}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [42],_al_u5461_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [42],\cu_ru/m_s_epc/n2 [42]}),
    .sr(rst_pad),
    .f({_al_u7002_o,open_n45926}),
    .q({open_n45930,\cu_ru/sepc [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7003|cu_ru/m_s_tval/reg0_b42  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n45931}),
    .b({\cu_ru/read_mtval_sel_lutinv ,_al_u5239_o}),
    .c({\cu_ru/stval [42],\cu_ru/m_s_tval/n3 [42]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [42],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7003_o,open_n45944}),
    .q({open_n45948,\cu_ru/stval [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7004|_al_u7633  (
    .b({_al_u7002_o,_al_u7631_o}),
    .c({_al_u7003_o,_al_u7632_o}),
    .d({_al_u7001_o,_al_u7630_o}),
    .f({_al_u7004_o,_al_u7633_o}));
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7005|biu/bus_unit/mmu/reg2_b54  (
    .a({_al_u6788_o,open_n45971}),
    .b({\cu_ru/read_mepc_sel_lutinv ,open_n45972}),
    .c({\cu_ru/mcycle [42],_al_u3047_o}),
    .clk(clk_pad),
    .d({\cu_ru/mepc [42],_al_u3046_o}),
    .sr(rst_pad),
    .f({_al_u7005_o,open_n45986}),
    .q({open_n45990,\biu/paddress [118]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7006|cu_ru/m_s_tvec/reg1_b42  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n45991}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u7005_o}),
    .c({mtime_pad[42],_al_u7006_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [42],_al_u7004_o}),
    .sr(rst_pad),
    .f({_al_u7006_o,csr_data[42]}),
    .q({open_n46011,\cu_ru/mtvec [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7008|cu_ru/m_s_scratch/reg1_b41  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n46012}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/stval [41]}),
    .c({satp[41],data_csr[41]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [41],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n46023,data_csr[41]}),
    .sr(rst_pad),
    .f({_al_u7008_o,_al_u5242_o}),
    .q({open_n46027,\cu_ru/sscratch [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7010|cu_ru/m_s_cause/reg0_b41  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [41],\cu_ru/scause [41]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [41],data_csr[41]}),
    .sr(rst_pad),
    .f({_al_u7010_o,open_n46044}),
    .q({open_n46048,\cu_ru/scause [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7011|cu_ru/m_cycle_event/reg0_b41  (
    .a({_al_u7009_o,open_n46049}),
    .b({_al_u7010_o,_al_u7008_o}),
    .c({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/minstret [41]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [41],_al_u6763_o}),
    .mi({open_n46060,\cu_ru/m_cycle_event/n4 [41]}),
    .sr(rst_pad),
    .f({_al_u7011_o,_al_u7009_o}),
    .q({open_n46064,\cu_ru/minstret [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7013|cu_ru/m_s_tval/reg1_b41  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n46065}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[41],\cu_ru/m_s_tval/n3 [41]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [41],_al_u6497_o}),
    .sr(rst_pad),
    .f({_al_u7013_o,open_n46083}),
    .q({open_n46087,\cu_ru/mtval [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7014|_al_u7012  (
    .a({open_n46088,_al_u6788_o}),
    .b({_al_u7012_o,\cu_ru/read_stvec_sel_lutinv }),
    .c({_al_u7013_o,\cu_ru/mcycle [41]}),
    .d({_al_u7011_o,\cu_ru/stvec [41]}),
    .f({_al_u7014_o,_al_u7012_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7015|cu_ru/m_s_epc/reg0_b41  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n46113}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [41],_al_u5465_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [41],\cu_ru/m_s_epc/n2 [41]}),
    .sr(rst_pad),
    .f({_al_u7015_o,open_n46130}),
    .q({open_n46134,\cu_ru/sepc [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7016|cu_ru/m_s_tvec/reg1_b41  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n46135}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u7015_o}),
    .c({\cu_ru/mepc [41],_al_u7016_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [41],_al_u7014_o}),
    .sr(rst_pad),
    .f({_al_u7016_o,csr_data[41]}),
    .q({open_n46151,\cu_ru/mtvec [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7018|cu_ru/m_s_scratch/reg1_b40  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n46152}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/stval [40]}),
    .c({satp[40],data_csr[40]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [40],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n46163,data_csr[40]}),
    .sr(rst_pad),
    .f({_al_u7018_o,_al_u5245_o}),
    .q({open_n46167,\cu_ru/sscratch [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7020|cu_ru/m_s_cause/reg0_b40  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [40],\cu_ru/scause [40]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [40],data_csr[40]}),
    .sr(rst_pad),
    .f({_al_u7020_o,open_n46184}),
    .q({open_n46188,\cu_ru/scause [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7021|cu_ru/m_cycle_event/reg0_b40  (
    .a({_al_u7019_o,open_n46189}),
    .b({_al_u7020_o,_al_u7018_o}),
    .c({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/minstret [40]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [40],_al_u6763_o}),
    .mi({open_n46193,\cu_ru/m_cycle_event/n4 [40]}),
    .sr(rst_pad),
    .f({_al_u7021_o,_al_u7019_o}),
    .q({open_n46208,\cu_ru/minstret [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7023|cu_ru/m_s_tval/reg1_b40  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n46209}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[40],\cu_ru/m_s_tval/n3 [40]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [40],_al_u6499_o}),
    .sr(rst_pad),
    .f({_al_u7023_o,open_n46227}),
    .q({open_n46231,\cu_ru/mtval [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7024|cu_ru/m_s_tvec/reg1_b40  (
    .b({_al_u7022_o,_al_u7025_o}),
    .c({_al_u7023_o,_al_u7026_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7021_o,_al_u7024_o}),
    .sr(rst_pad),
    .f({_al_u7024_o,csr_data[40]}),
    .q({open_n46249,\cu_ru/mtvec [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7025|cu_ru/m_s_tval/reg0_b40  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n46250}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5245_o}),
    .c({\cu_ru/mepc [40],\cu_ru/m_s_tval/n3 [40]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [40],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7025_o,open_n46267}),
    .q({open_n46271,\cu_ru/stval [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7026|cu_ru/m_s_epc/reg0_b40  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n46272}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [40],_al_u5469_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [40],\cu_ru/m_s_epc/n2 [40]}),
    .sr(rst_pad),
    .f({_al_u7026_o,open_n46289}),
    .q({open_n46293,\cu_ru/sepc [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7028|cu_ru/m_s_scratch/reg1_b39  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n46294}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/stval [39]}),
    .c({satp[39],data_csr[39]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [39],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n46298,data_csr[39]}),
    .sr(rst_pad),
    .f({_al_u7028_o,_al_u5251_o}),
    .q({open_n46313,\cu_ru/sscratch [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7030|cu_ru/m_s_cause/reg0_b39  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [39],\cu_ru/scause [39]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [39],data_csr[39]}),
    .sr(rst_pad),
    .f({_al_u7030_o,open_n46330}),
    .q({open_n46334,\cu_ru/scause [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7031|cu_ru/m_cycle_event/reg0_b39  (
    .a({_al_u7029_o,open_n46335}),
    .b({_al_u7030_o,_al_u7028_o}),
    .c({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/minstret [39]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [39],_al_u6763_o}),
    .mi({open_n46339,\cu_ru/m_cycle_event/n4 [39]}),
    .sr(rst_pad),
    .f({_al_u7031_o,_al_u7029_o}),
    .q({open_n46354,\cu_ru/minstret [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*~A))"),
    //.LUT1("(~(C*B)*~(D*~A))"),
    .INIT_LUT0(16'b0010101000111111),
    .INIT_LUT1(16'b0010101000111111),
    .MODE("LOGIC"))
    \_al_u7032|_al_u7214  (
    .a({_al_u6788_o,_al_u6788_o}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/read_time_sel_lutinv }),
    .c({mtime_pad[39],mtime_pad[35]}),
    .d({\cu_ru/mcycle [39],\cu_ru/mcycle [35]}),
    .f({_al_u7032_o,_al_u7214_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b1110110010100000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u7033|_al_u6025  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/stvec [39],\cu_ru/stvec [39]}),
    .d({\cu_ru/mtvec [39],\cu_ru/mtvec [39]}),
    .f({_al_u7033_o,\cu_ru/tvec [39]}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7034|cu_ru/m_s_tvec/reg1_b39  (
    .b({_al_u7032_o,_al_u7035_o}),
    .c({_al_u7033_o,_al_u7036_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7031_o,_al_u7034_o}),
    .sr(rst_pad),
    .f({_al_u7034_o,csr_data[39]}),
    .q({open_n46416,\cu_ru/mtvec [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7035|cu_ru/m_s_tval/reg1_b39  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n46417}),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [39],\cu_ru/m_s_tval/n3 [39]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [39],_al_u6503_o}),
    .sr(rst_pad),
    .f({_al_u7035_o,open_n46431}),
    .q({open_n46435,\cu_ru/mtval [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7036|cu_ru/m_s_epc/reg0_b39  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n46436}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [39],_al_u5477_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [39],\cu_ru/m_s_epc/n2 [39]}),
    .sr(rst_pad),
    .f({_al_u7036_o,open_n46453}),
    .q({open_n46457,\cu_ru/sepc [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7038|cu_ru/m_s_scratch/reg0_b38  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n46458}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [38]}),
    .c({\cu_ru/mscratch [38],data_csr[38]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [38],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n46469,data_csr[38]}),
    .sr(rst_pad),
    .f({_al_u7038_o,_al_u5481_o}),
    .q({open_n46473,\cu_ru/mscratch [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7040|cu_ru/m_s_cause/reg0_b38  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({satp[38],\cu_ru/scause [38]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [38],data_csr[38]}),
    .sr(rst_pad),
    .f({_al_u7040_o,open_n46490}),
    .q({open_n46494,\cu_ru/scause [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7041|cu_ru/m_cycle_event/reg0_b38  (
    .a({_al_u7039_o,open_n46495}),
    .b({_al_u7040_o,_al_u7038_o}),
    .c({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/minstret [38]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [38],_al_u6763_o}),
    .mi({open_n46506,\cu_ru/m_cycle_event/n4 [38]}),
    .sr(rst_pad),
    .f({_al_u7041_o,_al_u7039_o}),
    .q({open_n46510,\cu_ru/minstret [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7042|cu_ru/m_s_tval/reg1_b38  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n46511}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [38],\cu_ru/m_s_tval/n3 [38]}),
    .clk(clk_pad),
    .d({\cu_ru/stvec [38],_al_u6505_o}),
    .sr(rst_pad),
    .f({_al_u7042_o,open_n46529}),
    .q({open_n46533,\cu_ru/mtval [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7043|cu_ru/m_s_tval/reg0_b38  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n46534}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u5254_o}),
    .c({mtime_pad[38],\cu_ru/m_s_tval/n3 [38]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [38],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7043_o,open_n46547}),
    .q({open_n46551,\cu_ru/stval [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7044|_al_u7116  (
    .b({_al_u7042_o,_al_u7114_o}),
    .c({_al_u7043_o,_al_u7115_o}),
    .d({_al_u7041_o,_al_u7113_o}),
    .f({_al_u7044_o,_al_u7116_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7045|cu_ru/m_s_epc/reg0_b38  (
    .a({_al_u6788_o,open_n46574}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/mcycle [38],_al_u5481_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [38],\cu_ru/m_s_epc/n2 [38]}),
    .sr(rst_pad),
    .f({_al_u7045_o,open_n46591}),
    .q({open_n46595,\cu_ru/sepc [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7046|cu_ru/m_s_tvec/reg1_b38  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n46596}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u7045_o}),
    .c({\cu_ru/mepc [38],_al_u7046_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [38],_al_u7044_o}),
    .sr(rst_pad),
    .f({_al_u7046_o,csr_data[38]}),
    .q({open_n46616,\cu_ru/mtvec [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7048|cu_ru/m_s_scratch/reg1_b37  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n46617}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/stval [37]}),
    .c({satp[37],data_csr[37]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [37],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n46628,data_csr[37]}),
    .sr(rst_pad),
    .f({_al_u7048_o,_al_u5257_o}),
    .q({open_n46632,\cu_ru/sscratch [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7050|cu_ru/m_s_cause/reg0_b37  (
    .a({\cu_ru/read_mcause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [37],\cu_ru/scause [37]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [37],data_csr[37]}),
    .sr(rst_pad),
    .f({_al_u7050_o,open_n46649}),
    .q({open_n46653,\cu_ru/scause [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7051|cu_ru/m_s_scratch/reg0_b37  (
    .a({_al_u7049_o,open_n46654}),
    .b({_al_u7050_o,\cu_ru/sepc [37]}),
    .c({\cu_ru/read_mscratch_sel_lutinv ,data_csr[37]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [37],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n46665,data_csr[37]}),
    .sr(rst_pad),
    .f({_al_u7051_o,_al_u5485_o}),
    .q({open_n46669,\cu_ru/mscratch [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7053|cu_ru/m_s_tval/reg1_b37  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n46670}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[37],\cu_ru/m_s_tval/n3 [37]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [37],_al_u6507_o}),
    .sr(rst_pad),
    .f({_al_u7053_o,open_n46688}),
    .q({open_n46692,\cu_ru/mtval [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7054|cu_ru/m_s_tvec/reg1_b37  (
    .b({_al_u7052_o,_al_u7055_o}),
    .c({_al_u7053_o,_al_u7056_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7051_o,_al_u7054_o}),
    .sr(rst_pad),
    .f({_al_u7054_o,csr_data[37]}),
    .q({open_n46710,\cu_ru/mtvec [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7055|cu_ru/m_s_tval/reg0_b37  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n46711}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5257_o}),
    .c({\cu_ru/mepc [37],\cu_ru/m_s_tval/n3 [37]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [37],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7055_o,open_n46728}),
    .q({open_n46732,\cu_ru/stval [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7056|cu_ru/m_s_epc/reg0_b37  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n46733}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [37],_al_u5485_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [37],\cu_ru/m_s_epc/n2 [37]}),
    .sr(rst_pad),
    .f({_al_u7056_o,open_n46750}),
    .q({open_n46754,\cu_ru/sepc [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7058|cu_ru/m_s_cause/reg0_b36  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({satp[36],\cu_ru/scause [36]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [36],data_csr[36]}),
    .sr(rst_pad),
    .f({_al_u7058_o,open_n46771}),
    .q({open_n46775,\cu_ru/scause [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7059|cu_ru/m_s_epc/reg0_b36  (
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [36],_al_u5489_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u7058_o,\cu_ru/m_s_epc/n2 [36]}),
    .sr(rst_pad),
    .f({_al_u7059_o,open_n46794}),
    .q({open_n46798,\cu_ru/sepc [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7060|cu_ru/m_s_scratch/reg1_b36  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n46799}),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/stval [36]}),
    .c({\cu_ru/mcause [36],data_csr[36]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [36],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n46810,data_csr[36]}),
    .sr(rst_pad),
    .f({_al_u7060_o,_al_u5260_o}),
    .q({open_n46814,\cu_ru/sscratch [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7061|cu_ru/m_s_scratch/reg0_b36  (
    .a({_al_u7059_o,open_n46815}),
    .b({_al_u7060_o,\cu_ru/sepc [36]}),
    .c({\cu_ru/read_mscratch_sel_lutinv ,data_csr[36]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [36],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n46819,data_csr[36]}),
    .sr(rst_pad),
    .f({_al_u7061_o,_al_u5489_o}),
    .q({open_n46834,\cu_ru/mscratch [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"))
    \_al_u7062|_al_u7092  (
    .a({_al_u6788_o,_al_u6788_o}),
    .b({\cu_ru/read_mtvec_sel_lutinv ,\cu_ru/read_mtvec_sel_lutinv }),
    .c({\cu_ru/mcycle [36],\cu_ru/mcycle [27]}),
    .d({\cu_ru/mtvec [36],\cu_ru/mtvec [27]}),
    .f({_al_u7062_o,_al_u7092_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7063|cu_ru/m_s_tval/reg0_b36  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n46855}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u5260_o}),
    .c({mtime_pad[36],\cu_ru/m_s_tval/n3 [36]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [36],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7063_o,open_n46872}),
    .q({open_n46876,\cu_ru/stval [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7064|cu_ru/m_s_tvec/reg1_b36  (
    .b({_al_u7062_o,_al_u7065_o}),
    .c({_al_u7063_o,_al_u7066_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7061_o,_al_u7064_o}),
    .sr(rst_pad),
    .f({_al_u7064_o,csr_data[36]}),
    .q({open_n46894,\cu_ru/mtvec [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7066|cu_ru/m_s_tval/reg1_b36  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n46895}),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [36],\cu_ru/m_s_tval/n3 [36]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [36],_al_u6509_o}),
    .sr(rst_pad),
    .f({_al_u7066_o,open_n46909}),
    .q({open_n46913,\cu_ru/mtval [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7068|cu_ru/m_s_scratch/reg1_b31  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n46914}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/stval [31]}),
    .c({satp[31],data_csr[31]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [31],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n46918,data_csr[31]}),
    .sr(rst_pad),
    .f({_al_u7068_o,_al_u5275_o}),
    .q({open_n46933,\cu_ru/sscratch [31]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7070|cu_ru/m_s_cause/reg0_b31  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [31],\cu_ru/scause [31]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [31],data_csr[31]}),
    .sr(rst_pad),
    .f({_al_u7070_o,open_n46950}),
    .q({open_n46954,\cu_ru/scause [31]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D*C))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(B*A*~(D*C))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0000100010001000),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7071|_al_u7091  (
    .a({_al_u7069_o,_al_u7089_o}),
    .b({_al_u7070_o,_al_u7090_o}),
    .c({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/read_mcause_sel_lutinv }),
    .d({\cu_ru/mcause [31],\cu_ru/mcause [27]}),
    .f({_al_u7071_o,_al_u7091_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7073|_al_u7674  (
    .a({\cu_ru/read_time_sel_lutinv ,\cu_ru/read_time_sel_lutinv }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_stvec_sel_lutinv }),
    .c({mtime_pad[31],mtime_pad[8]}),
    .d({\cu_ru/stvec [31],\cu_ru/stvec [8]}),
    .f({_al_u7073_o,_al_u7674_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7074|cu_ru/m_s_tvec/reg1_b31  (
    .b({_al_u7072_o,_al_u7075_o}),
    .c({_al_u7073_o,_al_u7076_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7071_o,_al_u7074_o}),
    .sr(rst_pad),
    .f({_al_u7074_o,csr_data[31]}),
    .q({open_n47024,\cu_ru/mtvec [31]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7075|cu_ru/m_s_tval/reg1_b31  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n47025}),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [31],\cu_ru/m_s_tval/n3 [31]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [31],_al_u6519_o}),
    .sr(rst_pad),
    .f({_al_u7075_o,open_n47039}),
    .q({open_n47043,\cu_ru/mtval [31]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7076|cu_ru/m_s_epc/reg0_b31  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n47044}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [31],_al_u5509_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [31],\cu_ru/m_s_epc/n2 [31]}),
    .sr(rst_pad),
    .f({_al_u7076_o,open_n47061}),
    .q({open_n47065,\cu_ru/sepc [31]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u7078|_al_u7088  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/read_sscratch_sel_lutinv }),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/read_satp_sel_lutinv }),
    .c({satp[29],satp[27]}),
    .d({\cu_ru/sscratch [29],\cu_ru/sscratch [27]}),
    .f({_al_u7078_o,_al_u7088_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7080|cu_ru/m_s_cause/reg0_b29  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [29],\cu_ru/scause [29]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [29],data_csr[29]}),
    .sr(rst_pad),
    .f({_al_u7080_o,open_n47102}),
    .q({open_n47106,\cu_ru/scause [29]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7083|cu_ru/m_s_tval/reg1_b29  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n47107}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[29],\cu_ru/m_s_tval/n3 [29]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [29],_al_u6525_o}),
    .sr(rst_pad),
    .f({_al_u7083_o,open_n47121}),
    .q({open_n47125,\cu_ru/mtval [29]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7084|cu_ru/m_s_tvec/reg1_b29  (
    .b({_al_u7082_o,_al_u7085_o}),
    .c({_al_u7083_o,_al_u7086_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7081_o,_al_u7084_o}),
    .sr(rst_pad),
    .f({_al_u7084_o,csr_data[29]}),
    .q({open_n47147,\cu_ru/mtvec [29]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7085|cu_ru/m_s_tval/reg0_b29  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n47148}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5284_o}),
    .c({\cu_ru/mepc [29],\cu_ru/m_s_tval/n3 [29]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [29],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7085_o,open_n47165}),
    .q({open_n47169,\cu_ru/stval [29]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7086|cu_ru/m_s_epc/reg0_b29  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n47170}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [29],_al_u5521_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [29],\cu_ru/m_s_epc/n2 [29]}),
    .sr(rst_pad),
    .f({_al_u7086_o,open_n47187}),
    .q({open_n47191,\cu_ru/sepc [29]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7090|cu_ru/m_s_cause/reg0_b27  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [27],\cu_ru/scause [27]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [27],data_csr[27]}),
    .sr(rst_pad),
    .f({_al_u7090_o,open_n47208}),
    .q({open_n47212,\cu_ru/scause [27]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u7093|_al_u7616  (
    .a({\cu_ru/read_time_sel_lutinv ,\cu_ru/read_time_sel_lutinv }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_stvec_sel_lutinv }),
    .c({mtime_pad[27],mtime_pad[20]}),
    .d({\cu_ru/stvec [27],\cu_ru/stvec [20]}),
    .f({_al_u7093_o,_al_u7616_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7094|cu_ru/m_s_tvec/reg1_b27  (
    .b({_al_u7092_o,_al_u7095_o}),
    .c({_al_u7093_o,_al_u7096_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7091_o,_al_u7094_o}),
    .sr(rst_pad),
    .f({_al_u7094_o,csr_data[27]}),
    .q({open_n47250,\cu_ru/mtvec [27]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7095|cu_ru/m_s_epc/reg0_b27  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n47251}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [27],_al_u5529_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [27],\cu_ru/m_s_epc/n2 [27]}),
    .sr(rst_pad),
    .f({_al_u7095_o,open_n47268}),
    .q({open_n47272,\cu_ru/sepc [27]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7096|cu_ru/m_s_tval/reg0_b27  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n47273}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5290_o}),
    .c({\cu_ru/mepc [27],\cu_ru/m_s_tval/n3 [27]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [27],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7096_o,open_n47286}),
    .q({open_n47290,\cu_ru/stval [27]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u7098|_al_u7237  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/read_sscratch_sel_lutinv }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/read_mcause_sel_lutinv }),
    .c(\cu_ru/mcause [26:25]),
    .d(\cu_ru/sscratch [26:25]),
    .f({_al_u7098_o,_al_u7237_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7101|cu_ru/m_s_scratch/reg0_b26  (
    .a({\cu_ru/read_mscratch_sel_lutinv ,open_n47311}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/sepc [26]}),
    .c({satp[26],data_csr[26]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [26],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n47322,data_csr[26]}),
    .sr(rst_pad),
    .f({_al_u7101_o,_al_u5533_o}),
    .q({open_n47326,\cu_ru/mscratch [26]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7102|cu_ru/m_cycle_event/reg0_b26  (
    .a({open_n47327,\cu_ru/read_minstret_sel_lutinv }),
    .b({_al_u7100_o,\cu_ru/read_scause_sel_lutinv }),
    .c({_al_u7101_o,\cu_ru/minstret [26]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7099_o,\cu_ru/scause [26]}),
    .mi({open_n47338,\cu_ru/m_cycle_event/n4 [26]}),
    .sr(rst_pad),
    .f({_al_u7102_o,_al_u7100_o}),
    .q({open_n47342,\cu_ru/minstret [26]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7103|cu_ru/m_s_epc/reg0_b26  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n47343}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [26],_al_u5533_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [26],\cu_ru/m_s_epc/n2 [26]}),
    .sr(rst_pad),
    .f({_al_u7103_o,open_n47360}),
    .q({open_n47364,\cu_ru/sepc [26]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7104|cu_ru/m_s_tval/reg0_b26  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n47365}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u5293_o}),
    .c({\cu_ru/stval [26],\cu_ru/m_s_tval/n3 [26]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [26],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7104_o,open_n47382}),
    .q({open_n47386,\cu_ru/stval [26]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7106|cu_ru/m_s_tvec/reg1_b26  (
    .a({_al_u6788_o,open_n47387}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u7106_o}),
    .c({\cu_ru/mcycle [26],_al_u7107_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [26],_al_u7105_o}),
    .sr(rst_pad),
    .f({_al_u7106_o,csr_data[26]}),
    .q({open_n47403,\cu_ru/mtvec [26]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7107|cu_ru/m_s_tval/reg1_b26  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n47404}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[26],\cu_ru/m_s_tval/n3 [26]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [26],_al_u6531_o}),
    .sr(rst_pad),
    .f({_al_u7107_o,open_n47422}),
    .q({open_n47426,\cu_ru/mtval [26]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7110|_al_u7109  (
    .a({open_n47427,\cu_ru/read_sscratch_sel_lutinv }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/read_satp_sel_lutinv }),
    .c({\cu_ru/mcause [24],satp[24]}),
    .d({_al_u7109_o,\cu_ru/sscratch [24]}),
    .f({_al_u7110_o,_al_u7109_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7111|cu_ru/m_s_cause/reg0_b24  (
    .a({\cu_ru/read_minstret_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/minstret [24],\cu_ru/scause [24]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [24],data_csr[24]}),
    .sr(rst_pad),
    .f({_al_u7111_o,open_n47468}),
    .q({open_n47472,\cu_ru/scause [24]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7113|cu_ru/m_cycle_event/reg0_b24  (
    .a({open_n47473,\cu_ru/read_instret_sel_lutinv }),
    .b({_al_u7111_o,\cu_ru/read_mscratch_sel_lutinv }),
    .c({_al_u7112_o,\cu_ru/minstret [24]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7110_o,\cu_ru/mscratch [24]}),
    .mi({open_n47477,\cu_ru/m_cycle_event/n4 [24]}),
    .sr(rst_pad),
    .f({_al_u7113_o,_al_u7112_o}),
    .q({open_n47492,\cu_ru/minstret [24]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7114|cu_ru/m_s_epc/reg0_b24  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n47493}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [24],_al_u5541_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [24],\cu_ru/m_s_epc/n2 [24]}),
    .sr(rst_pad),
    .f({_al_u7114_o,open_n47510}),
    .q({open_n47514,\cu_ru/sepc [24]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7115|cu_ru/m_s_tval/reg0_b24  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n47515}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u5299_o}),
    .c({\cu_ru/stval [24],\cu_ru/m_s_tval/n3 [24]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [24],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7115_o,open_n47528}),
    .q({open_n47532,\cu_ru/stval [24]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(~(C*B)*~(D*~A))"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(~(C*B)*~(D*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b0010101000111111),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b0010101000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7117|cu_ru/m_s_tvec/reg1_b24  (
    .a({_al_u6788_o,open_n47533}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u7117_o}),
    .c({mtime_pad[24],_al_u7118_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mcycle [24],_al_u7116_o}),
    .sr(rst_pad),
    .f({_al_u7117_o,csr_data[24]}),
    .q({open_n47553,\cu_ru/mtvec [24]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7118|cu_ru/m_s_tval/reg1_b24  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n47554}),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [24],\cu_ru/m_s_tval/n3 [24]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [24],_al_u6535_o}),
    .sr(rst_pad),
    .f({_al_u7118_o,open_n47568}),
    .q({open_n47572,\cu_ru/mtval [24]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7120|biu/bus_unit/mmu/reg2_b35  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n47573}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n47574}),
    .c({satp[23],_al_u3104_o}),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [23],_al_u3103_o}),
    .sr(rst_pad),
    .f({_al_u7120_o,open_n47592}),
    .q({open_n47596,\biu/paddress [99]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u7121|_al_u7081  (
    .a({open_n47597,_al_u7079_o}),
    .b({\cu_ru/read_mcause_sel_lutinv ,_al_u7080_o}),
    .c({\cu_ru/mcause [23],\cu_ru/read_mcause_sel_lutinv }),
    .d({_al_u7120_o,\cu_ru/mcause [29]}),
    .f({_al_u7121_o,_al_u7081_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7122|cu_ru/m_s_cause/reg0_b23  (
    .a({\cu_ru/read_minstret_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/minstret [23],\cu_ru/scause [23]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [23],data_csr[23]}),
    .sr(rst_pad),
    .f({_al_u7122_o,open_n47634}),
    .q({open_n47638,\cu_ru/scause [23]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7124|cu_ru/m_cycle_event/reg0_b23  (
    .a({open_n47639,\cu_ru/read_instret_sel_lutinv }),
    .b({_al_u7122_o,\cu_ru/read_mscratch_sel_lutinv }),
    .c({_al_u7123_o,\cu_ru/minstret [23]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7121_o,\cu_ru/mscratch [23]}),
    .mi({open_n47643,\cu_ru/m_cycle_event/n4 [23]}),
    .sr(rst_pad),
    .f({_al_u7124_o,_al_u7123_o}),
    .q({open_n47658,\cu_ru/minstret [23]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7125|cu_ru/m_s_epc/reg0_b23  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n47659}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [23],_al_u5545_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [23],\cu_ru/m_s_epc/n2 [23]}),
    .sr(rst_pad),
    .f({_al_u7125_o,open_n47676}),
    .q({open_n47680,\cu_ru/sepc [23]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7126|cu_ru/m_s_tval/reg0_b23  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n47681}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u5302_o}),
    .c({\cu_ru/stval [23],\cu_ru/m_s_tval/n3 [23]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [23],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7126_o,open_n47694}),
    .q({open_n47698,\cu_ru/stval [23]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7127|_al_u7099  (
    .b({_al_u7125_o,\cu_ru/read_instret_sel_lutinv }),
    .c({_al_u7126_o,\cu_ru/minstret [26]}),
    .d({_al_u7124_o,_al_u7098_o}),
    .f({_al_u7127_o,_al_u7099_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(~(C*B)*~(D*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b0010101000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7128|cu_ru/m_s_tvec/reg1_b23  (
    .a({_al_u6788_o,open_n47721}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u7128_o}),
    .c({mtime_pad[23],_al_u7129_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mcycle [23],_al_u7127_o}),
    .sr(rst_pad),
    .f({_al_u7128_o,csr_data[23]}),
    .q({open_n47737,\cu_ru/mtvec [23]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7129|cu_ru/m_s_tval/reg1_b23  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n47738}),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [23],\cu_ru/m_s_tval/n3 [23]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [23],_al_u6537_o}),
    .sr(rst_pad),
    .f({_al_u7129_o,open_n47756}),
    .q({open_n47760,\cu_ru/mtval [23]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7131|biu/bus_unit/mmu/reg2_b28  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n47761}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n47762}),
    .c({satp[16],_al_u3125_o}),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [16],_al_u3124_o}),
    .sr(rst_pad),
    .f({_al_u7131_o,open_n47780}),
    .q({open_n47784,\biu/paddress [92]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7133|cu_ru/m_s_cause/reg0_b16  (
    .a({\cu_ru/read_mcause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [16],\cu_ru/scause [16]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [16],data_csr[16]}),
    .sr(rst_pad),
    .f({_al_u7133_o,open_n47801}),
    .q({open_n47805,\cu_ru/scause [16]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7134|cu_ru/m_s_scratch/reg0_b16  (
    .a({_al_u7132_o,open_n47806}),
    .b({_al_u7133_o,\cu_ru/sepc [16]}),
    .c({\cu_ru/read_mscratch_sel_lutinv ,data_csr[16]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [16],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n47817,data_csr[16]}),
    .sr(rst_pad),
    .f({_al_u7134_o,_al_u5577_o}),
    .q({open_n47821,\cu_ru/mscratch [16]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7136|cu_ru/m_s_tval/reg1_b16  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n47822}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[16],\cu_ru/m_s_tval/n3 [16]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [16],_al_u6553_o}),
    .sr(rst_pad),
    .f({_al_u7136_o,open_n47840}),
    .q({open_n47844,\cu_ru/mtval [16]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7137|_al_u7135  (
    .a({open_n47845,_al_u6788_o}),
    .b({_al_u7135_o,\cu_ru/read_stvec_sel_lutinv }),
    .c({_al_u7136_o,\cu_ru/mcycle [16]}),
    .d({_al_u7134_o,\cu_ru/stvec [16]}),
    .f({_al_u7137_o,_al_u7135_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7138|cu_ru/m_s_epc/reg0_b16  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n47866}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [16],_al_u5577_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [16],\cu_ru/m_s_epc/n2 [16]}),
    .sr(rst_pad),
    .f({_al_u7138_o,open_n47883}),
    .q({open_n47887,\cu_ru/sepc [16]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7139|cu_ru/m_s_tvec/reg1_b16  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n47888}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u7138_o}),
    .c({\cu_ru/mepc [16],_al_u7139_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [16],_al_u7137_o}),
    .sr(rst_pad),
    .f({_al_u7139_o,csr_data[16]}),
    .q({open_n47904,\cu_ru/mtvec [16]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~A*~(D*C))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("~(B*~A*~(D*C))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101110111011),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111101110111011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7143|ins_dec/ill_ins_reg  (
    .a({_al_u3956_o,\ins_dec/dec_ins_dec_fault_lutinv }),
    .b({_al_u4161_o,_al_u7147_o}),
    .c({_al_u7141_o,tvm}),
    .ce(\ins_dec/u461_sel_is_0_o ),
    .clk(clk_pad),
    .d({_al_u7142_o,\ins_dec/ins_sfencevma }),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/dec_ins_dec_fault_lutinv ,id_ill_ins}),
    .q({open_n47924,ex_ill_ins}));  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u7144|_al_u7240  (
    .b({_al_u3400_o,id_ins[24]}),
    .c({id_ins[25],id_ins[23]}),
    .d({_al_u3399_o,id_ins[25]}),
    .f({\ins_dec/funct7_8_lutinv ,_al_u7240_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7146|cu_ru/m_s_status/tw_reg  (
    .a({open_n47947,\cu_ru/read_mcycle_sel_lutinv }),
    .b({open_n47948,\cu_ru/n90 [32]}),
    .c({tw,\cu_ru/mcycle [21]}),
    .ce(\cu_ru/m_s_status/n0 ),
    .clk(clk_pad),
    .d({id_system,tw}),
    .mi({open_n47959,data_csr[21]}),
    .sr(rst_pad),
    .f({_al_u7146_o,_al_u7255_o}),
    .q({open_n47963,tw}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(D*B)*~(~C*A))"),
    .INIT_LUT0(16'b1111110011000111),
    .INIT_LUT1(16'b0011000111110101),
    .MODE("LOGIC"))
    \_al_u7147|_al_u7145  (
    .a({\ins_dec/n239 ,\ins_dec/n80_lutinv }),
    .b({\ins_dec/funct7_8_lutinv ,priv[0]}),
    .c({_al_u7145_o,priv[1]}),
    .d({_al_u7146_o,priv[3]}),
    .f({_al_u7147_o,_al_u7145_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("(D*(C@B))"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("(D*(C@B))"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b0011110000000000),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b0011110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7150|_al_u3950  (
    .b({\biu/cache_ctrl_logic/statu [0],\biu/cache_ctrl_logic/statu [0]}),
    .c({\biu/cache_ctrl_logic/statu [1],\biu/cache_ctrl_logic/statu [1]}),
    .d({_al_u3944_o,_al_u3944_o}),
    .f({_al_u7150_o,_al_u3950_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(~A*~(~B*~(D*~C)))"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(~A*~(~B*~(D*~C)))"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b0100010101000100),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b0100010101000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7152|_al_u9274  (
    .a({\biu/cache_ctrl_logic/n97_lutinv ,open_n48010}),
    .b({_al_u7150_o,_al_u7150_o}),
    .c({_al_u7151_o,_al_u7151_o}),
    .d({\biu/cache_ctrl_logic/statu [4],_al_u3945_o}),
    .f({_al_u7152_o,_al_u9274_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~D*C*B))"),
    //.LUT1("(C*~(B*~(D*A)))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b1011000000110000),
    .MODE("LOGIC"))
    \_al_u7154|_al_u7153  (
    .a({_al_u7149_o,_al_u3224_o}),
    .b({_al_u7152_o,_al_u2847_o}),
    .c({\biu/cache_ctrl_logic/mux31_b4_sel_is_2_o ,\biu/cache_ctrl_logic/statu [3]}),
    .d({_al_u7150_o,\biu/cache_ctrl_logic/statu [4]}),
    .f({_al_u7154_o,\biu/cache_ctrl_logic/mux31_b4_sel_is_2_o }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7155|_al_u9677  (
    .c({\biu/cache_ctrl_logic/mux31_b4_sel_is_2_o ,_al_u3950_o}),
    .d({_al_u7149_o,_al_u7149_o}),
    .f({_al_u7155_o,_al_u9677_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*~(B*~(D*A)))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000101100000011),
    .MODE("LOGIC"))
    \_al_u7156|_al_u9129  (
    .a({\biu/cache_ctrl_logic/n100 [4],open_n48083}),
    .b({_al_u7154_o,open_n48084}),
    .c({_al_u7155_o,_al_u3224_o}),
    .d({\biu/cache_ctrl_logic/n97_lutinv ,\biu/cache_ctrl_logic/n100 [4]}),
    .f({_al_u7156_o,_al_u9129_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*C*A))"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0001001100110011),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u7157|_al_u7149  (
    .a({open_n48105,_al_u2705_o}),
    .b({_al_u4195_o,_al_u3407_o}),
    .c({\biu/bus_unit/mmu/statu [0],_al_u4195_o}),
    .d({_al_u2705_o,\biu/bus_unit/mmu/statu [0]}),
    .f({_al_u7157_o,_al_u7149_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(~B*~(C*~A)))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(~B*~(C*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000011011100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000011011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u7161|biu/cache_ctrl_logic/reg8_b4  (
    .a({_al_u7156_o,open_n48126}),
    .b({_al_u7158_o,_al_u7192_o}),
    .c({_al_u7159_o,_al_u7193_o}),
    .clk(clk_pad),
    .d({_al_u7160_o,_al_u7161_o}),
    .sr(\biu/cache_ctrl_logic/mux44_b4_sel_is_2_o ),
    .f({_al_u7161_o,open_n48144}),
    .q({open_n48148,\biu/cache_ctrl_logic/statu [4]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7162|_al_u6361  (
    .b({open_n48151,\biu/cache_ctrl_logic/n55_lutinv }),
    .c({\biu/cache_ctrl_logic/n55_lutinv ,_al_u6360_o}),
    .d({_al_u6426_o,_al_u6323_o}),
    .f({_al_u7162_o,\biu/cache/n15 }));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1000001001000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7164|biu/bus_unit/mmu/reg1_b53  (
    .a({cacheability_block_pad[21],open_n48176}),
    .b({cacheability_block_pad[1],open_n48177}),
    .c({\biu/paddress [33],_al_u5026_o}),
    .clk(clk_pad),
    .d({\biu/paddress [53],_al_u5025_o}),
    .sr(rst_pad),
    .f({_al_u7164_o,open_n48191}),
    .q({open_n48195,\biu/paddress [53]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*~B)*~(D*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1000101011001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7165|biu/bus_unit/mmu/reg1_b54  (
    .a({cacheability_block_pad[22],open_n48196}),
    .b({cacheability_block_pad[12],open_n48197}),
    .c({\biu/paddress [44],_al_u5023_o}),
    .clk(clk_pad),
    .d({\biu/paddress [54],_al_u5022_o}),
    .sr(rst_pad),
    .f({_al_u7165_o,open_n48211}),
    .q({open_n48215,\biu/paddress [54]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7166|biu/bus_unit/mmu/reg1_b42  (
    .a({_al_u7164_o,open_n48216}),
    .b({_al_u7165_o,open_n48217}),
    .c({cacheability_block_pad[10],_al_u5059_o}),
    .clk(clk_pad),
    .d({\biu/paddress [42],_al_u5058_o}),
    .sr(rst_pad),
    .f({_al_u7166_o,open_n48235}),
    .q({open_n48239,\biu/paddress [42]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1000001001000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7167|biu/cache_ctrl_logic/reg6_b58  (
    .a({cacheability_block_pad[26],open_n48240}),
    .b({cacheability_block_pad[18],\biu/paddress [58]}),
    .c({\biu/paddress [50],\biu/cache_ctrl_logic/pa_temp [58]}),
    .clk(clk_pad),
    .d({\biu/paddress [58],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u7167_o,open_n48254}),
    .q({open_n48258,\biu/cache_ctrl_logic/pa_temp [58]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7168|biu/bus_unit/mmu/reg1_b34  (
    .a({cacheability_block_pad[2],open_n48259}),
    .b({cacheability_block_pad[0],open_n48260}),
    .c({\biu/paddress [32],_al_u5083_o}),
    .clk(clk_pad),
    .d({\biu/paddress [34],_al_u5082_o}),
    .sr(rst_pad),
    .f({_al_u7168_o,open_n48278}),
    .q({open_n48282,\biu/paddress [34]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1000001001000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7170|biu/cache_ctrl_logic/reg6_b62  (
    .a({cacheability_block_pad[30],open_n48283}),
    .b({cacheability_block_pad[28],\biu/paddress [62]}),
    .c({\biu/paddress [60],\biu/cache_ctrl_logic/pa_temp [62]}),
    .clk(clk_pad),
    .d({\biu/paddress [62],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u7170_o,open_n48297}),
    .q({open_n48301,\biu/cache_ctrl_logic/pa_temp [62]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(B*A*~(D@C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7171|biu/cache_ctrl_logic/reg6_b61  (
    .a({_al_u3411_o,open_n48302}),
    .b({_al_u7170_o,\biu/paddress [61]}),
    .c({cacheability_block_pad[29],\biu/cache_ctrl_logic/pa_temp [61]}),
    .clk(clk_pad),
    .d({\biu/paddress [61],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u7171_o,open_n48316}),
    .q({open_n48320,\biu/cache_ctrl_logic/pa_temp [61]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7172|biu/cache_ctrl_logic/reg6_b56  (
    .a({cacheability_block_pad[24],open_n48321}),
    .b({cacheability_block_pad[20],\biu/paddress [56]}),
    .c({\biu/paddress [52],\biu/cache_ctrl_logic/pa_temp [56]}),
    .clk(clk_pad),
    .d({\biu/paddress [56],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u7172_o,open_n48339}),
    .q({open_n48343,\biu/cache_ctrl_logic/pa_temp [56]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111001101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7173|biu/bus_unit/mmu/reg1_b44  (
    .a({cacheability_block_pad[22],open_n48344}),
    .b({cacheability_block_pad[12],open_n48345}),
    .c({\biu/paddress [44],_al_u5053_o}),
    .clk(clk_pad),
    .d({\biu/paddress [54],_al_u5052_o}),
    .sr(rst_pad),
    .f({_al_u7173_o,open_n48359}),
    .q({open_n48363,\biu/paddress [44]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7174|biu/bus_unit/mmu/reg1_b45  (
    .a({_al_u7172_o,open_n48364}),
    .b({_al_u7173_o,open_n48365}),
    .c({cacheability_block_pad[13],_al_u5050_o}),
    .clk(clk_pad),
    .d({\biu/paddress [45],_al_u5049_o}),
    .sr(rst_pad),
    .f({_al_u7174_o,open_n48383}),
    .q({open_n48387,\biu/paddress [45]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7175|_al_u4196  (
    .b({_al_u7171_o,open_n48390}),
    .c({_al_u7174_o,_al_u4195_o}),
    .d({_al_u7169_o,_al_u3411_o}),
    .f({_al_u7175_o,\biu/bus_unit/mmu/mux10_b0_sel_is_2_o }));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7176|biu/cache_ctrl_logic/reg6_b59  (
    .a({cacheability_block_pad[27],open_n48411}),
    .b({cacheability_block_pad[23],\biu/paddress [59]}),
    .c({\biu/paddress [55],\biu/cache_ctrl_logic/pa_temp [59]}),
    .clk(clk_pad),
    .d({\biu/paddress [59],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u7176_o,open_n48429}),
    .q({open_n48433,\biu/cache_ctrl_logic/pa_temp [59]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7177|biu/bus_unit/mmu/reg1_b51  (
    .a({cacheability_block_pad[19],open_n48434}),
    .b({cacheability_block_pad[8],open_n48435}),
    .c({\biu/paddress [40],_al_u5032_o}),
    .clk(clk_pad),
    .d({\biu/paddress [51],_al_u5031_o}),
    .sr(rst_pad),
    .f({_al_u7177_o,open_n48453}),
    .q({open_n48457,\biu/paddress [51]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1000001001000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7178|biu/cache_ctrl_logic/reg6_b57  (
    .a({cacheability_block_pad[25],open_n48458}),
    .b({cacheability_block_pad[3],\biu/paddress [57]}),
    .c({\biu/paddress [35],\biu/cache_ctrl_logic/pa_temp [57]}),
    .clk(clk_pad),
    .d({\biu/paddress [57],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u7178_o,open_n48472}),
    .q({open_n48476,\biu/cache_ctrl_logic/pa_temp [57]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7179|biu/bus_unit/mmu/reg1_b39  (
    .a({cacheability_block_pad[7],open_n48477}),
    .b({cacheability_block_pad[4],open_n48478}),
    .c({\biu/paddress [36],_al_u5068_o}),
    .clk(clk_pad),
    .d({\biu/paddress [39],_al_u5067_o}),
    .sr(rst_pad),
    .f({_al_u7179_o,open_n48496}),
    .q({open_n48500,\biu/paddress [39]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7180|biu/bus_unit/mmu/reg1_b55  (
    .a({_al_u7176_o,open_n48501}),
    .b({_al_u7177_o,open_n48502}),
    .c({_al_u7178_o,_al_u5020_o}),
    .clk(clk_pad),
    .d({_al_u7179_o,_al_u5019_o}),
    .sr(rst_pad),
    .f({_al_u7180_o,open_n48520}),
    .q({open_n48524,\biu/paddress [55]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1000001001000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7181|biu/bus_unit/mmu/reg1_b47  (
    .a({cacheability_block_pad[15],open_n48525}),
    .b({cacheability_block_pad[9],open_n48526}),
    .c({\biu/paddress [41],_al_u5044_o}),
    .clk(clk_pad),
    .d({\biu/paddress [47],_al_u5043_o}),
    .sr(rst_pad),
    .f({_al_u7181_o,open_n48540}),
    .q({open_n48544,\biu/paddress [47]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7182|biu/bus_unit/mmu/reg1_b38  (
    .a({_al_u7180_o,open_n48545}),
    .b({_al_u7181_o,open_n48546}),
    .c({cacheability_block_pad[6],_al_u5071_o}),
    .clk(clk_pad),
    .d({\biu/paddress [38],_al_u5070_o}),
    .sr(rst_pad),
    .f({_al_u7182_o,open_n48564}),
    .q({open_n48568,\biu/paddress [38]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(~(C*~B)*~(~D*A))"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(~(C*~B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b1100111101000101),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1100111101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7183|biu/cache_ctrl_logic/reg6_b63  (
    .a({cacheability_block_pad[31],open_n48569}),
    .b({cacheability_block_pad[17],\biu/paddress [63]}),
    .c({\biu/paddress [49],\biu/cache_ctrl_logic/pa_temp [63]}),
    .clk(clk_pad),
    .d({\biu/paddress [63],\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .f({_al_u7183_o,open_n48587}),
    .q({open_n48591,\biu/cache_ctrl_logic/pa_temp [63]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*~B)*~(~D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*~B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1100111101000101),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1100111101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7184|biu/bus_unit/mmu/reg1_b49  (
    .a({cacheability_block_pad[17],open_n48592}),
    .b({cacheability_block_pad[16],open_n48593}),
    .c({\biu/paddress [48],_al_u5038_o}),
    .clk(clk_pad),
    .d({\biu/paddress [49],_al_u5037_o}),
    .sr(rst_pad),
    .f({_al_u7184_o,open_n48611}),
    .q({open_n48615,\biu/paddress [49]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(~C*B)*~(~D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(~C*B)*~(~D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111001101010001),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111001101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7185|biu/bus_unit/mmu/reg1_b48  (
    .a({cacheability_block_pad[16],open_n48616}),
    .b({cacheability_block_pad[11],open_n48617}),
    .c({\biu/paddress [43],_al_u5041_o}),
    .clk(clk_pad),
    .d({\biu/paddress [48],_al_u5040_o}),
    .sr(rst_pad),
    .f({_al_u7185_o,open_n48635}),
    .q({open_n48639,\biu/paddress [48]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*~B)*~(D*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1000101011001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7186|biu/bus_unit/mmu/reg1_b43  (
    .a({cacheability_block_pad[31],open_n48640}),
    .b({cacheability_block_pad[11],open_n48641}),
    .c({\biu/paddress [43],_al_u5056_o}),
    .clk(clk_pad),
    .d({\biu/paddress [63],_al_u5055_o}),
    .sr(rst_pad),
    .f({_al_u7186_o,open_n48655}),
    .q({open_n48659,\biu/paddress [43]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u7187|_al_u7189  (
    .a({_al_u7183_o,_al_u7175_o}),
    .b({_al_u7184_o,_al_u7182_o}),
    .c({_al_u7185_o,_al_u7187_o}),
    .d({_al_u7186_o,_al_u7188_o}),
    .f({_al_u7187_o,\biu/cacheable }));
  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1000001001000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7188|biu/bus_unit/mmu/reg1_b46  (
    .a({cacheability_block_pad[14],open_n48680}),
    .b({cacheability_block_pad[5],open_n48681}),
    .c({\biu/paddress [37],_al_u5047_o}),
    .clk(clk_pad),
    .d({\biu/paddress [46],_al_u5046_o}),
    .sr(rst_pad),
    .f({_al_u7188_o,open_n48695}),
    .q({open_n48699,\biu/paddress [46]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*~A)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u7190|_al_u9280  (
    .a({open_n48700,\biu/cache_ctrl_logic/n100 [4]}),
    .b({open_n48701,_al_u7158_o}),
    .c({\biu/cacheable ,\biu/cacheable }),
    .d({\biu/cache_ctrl_logic/n100 [4],_al_u6257_o}),
    .f({_al_u7190_o,_al_u9280_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u7191|_al_u4812  (
    .a({open_n48722,_al_u4809_o}),
    .b({open_n48723,_al_u4811_o}),
    .c({\biu/bus_unit/mmu/n19_lutinv ,\biu/bus_unit/mmu/n19_lutinv }),
    .d({_al_u7157_o,addr_if[2]}),
    .f({_al_u7191_o,_al_u4812_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~A*~(D*~(~C*~B)))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~A*~(D*~(~C*~B)))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000101010101),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7192|_al_u7163  (
    .a({_al_u7162_o,open_n48744}),
    .b({_al_u7163_o,open_n48745}),
    .c({_al_u7190_o,_al_u7149_o}),
    .d({_al_u7191_o,\biu/cache_ctrl_logic/n100 [4]}),
    .f({_al_u7192_o,_al_u7163_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7195|_al_u3221  (
    .c({_al_u3209_o,_al_u3209_o}),
    .d({_al_u2835_o,_al_u2838_o}),
    .f({_al_u7195_o,\biu/cache_ctrl_logic/n97_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*D))"),
    //.LUTF1("(C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("(~C*~(B*D))"),
    //.LUTG1("(C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b0000001100001111),
    .INIT_LUTF1(16'b0001000010110000),
    .INIT_LUTG0(16'b0000001100001111),
    .INIT_LUTG1(16'b0001000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7200|_al_u7199  (
    .a({\biu/bus_unit/mmu/n12_lutinv ,open_n48798}),
    .b({_al_u7198_o,\biu/bus_unit/mmu_hwdata [3]}),
    .c({_al_u7199_o,priv[3]}),
    .d({\biu/bus_unit/mmu_hwdata [2],\biu/bus_unit/mmu/n19_lutinv }),
    .f({_al_u7200_o,_al_u7199_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~C*B*~D)"),
    .INIT_LUTF0(16'b1111110011000111),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b1111110011000111),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7202|_al_u7201  (
    .a({open_n48823,\biu/bus_unit/mmu_hwdata [4]}),
    .b({_al_u2915_o,priv[0]}),
    .c({_al_u7201_o,priv[1]}),
    .d({_al_u7200_o,priv[3]}),
    .f({_al_u7202_o,_al_u7201_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7203|_al_u7206  (
    .b({open_n48850,_al_u7205_o}),
    .c({\biu/bus_unit/mmu/n37_lutinv ,_al_u2915_o}),
    .d({_al_u7202_o,_al_u7203_o}),
    .f({_al_u7203_o,_al_u7206_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(~(C*B)*~(D*~A))"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(~(C*B)*~(D*~A))"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b0010101000111111),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b0010101000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7205|_al_u4195  (
    .a({_al_u4195_o,open_n48875}),
    .b({\biu/bus_unit/mmu/n45_lutinv ,\biu/bus_unit/mmu/statu [2]}),
    .c({hresp_pad,\biu/bus_unit/mmu/statu [3]}),
    .d({\biu/bus_unit/mmu/statu [3],\biu/bus_unit/mmu/statu [1]}),
    .f({_al_u7205_o,_al_u4195_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7208|_al_u4775  (
    .b({\biu/bus_unit/mmu/n37_lutinv ,_al_u2705_o}),
    .c({\biu/bus_unit/mmu_hwdata [6],\biu/bus_unit/mmu_hwdata [6]}),
    .d({\biu/bus_unit/mmu/n2 ,_al_u4774_o}),
    .f({_al_u7208_o,hwdata_pad[6]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(B*~(A*~(~D*~C)))"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(B*~(A*~(~D*~C)))"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0100010001001100),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0100010001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7210|_al_u4135  (
    .a({\cu_ru/medeleg_exc_ctrl/n85_neg_lutinv ,wb_ill_ins}),
    .b({\cu_ru/medeleg_exc_ctrl/n84_neg_lutinv ,wb_ld_acc_fault}),
    .c({_al_u4106_o,wb_ld_addr_mis}),
    .d({\cu_ru/medeleg_exc_ctrl/n87_neg_lutinv ,wb_ld_page_fault}),
    .f({_al_u7210_o,_al_u4135_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~((~D*~A))*~(B)+C*(~D*~A)*~(B)+~(C)*(~D*~A)*B+C*(~D*~A)*B)"),
    //.LUTF1("(~D*C*~(~B*~A))"),
    //.LUTG0("~(C*~((~D*~A))*~(B)+C*(~D*~A)*~(B)+~(C)*(~D*~A)*B+C*(~D*~A)*B)"),
    //.LUTG1("(~D*C*~(~B*~A))"),
    .INIT_LUTF0(16'b1100111110001011),
    .INIT_LUTF1(16'b0000000011100000),
    .INIT_LUTG0(16'b1100111110001011),
    .INIT_LUTG1(16'b0000000011100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7212|_al_u7213  (
    .a({_al_u7211_o,_al_u7212_o}),
    .b({_al_u4117_o,_al_u4138_o}),
    .c({_al_u5099_o,_al_u4233_o}),
    .d({_al_u5154_o,_al_u4141_o}),
    .f({_al_u7212_o,\cu_ru/trap_cause [1]}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7215|cu_ru/m_s_cause/reg0_b35  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [35],\cu_ru/scause [35]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [35],data_csr[35]}),
    .sr(rst_pad),
    .f({_al_u7215_o,open_n48990}),
    .q({open_n48994,\cu_ru/scause [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7216|cu_ru/m_s_scratch/reg1_b35  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n48995}),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/stval [35]}),
    .c({\cu_ru/mcause [35],data_csr[35]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [35],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n48999,data_csr[35]}),
    .sr(rst_pad),
    .f({_al_u7216_o,_al_u5263_o}),
    .q({open_n49014,\cu_ru/sscratch [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7217|_al_u6786  (
    .c({_al_u6791_o,_al_u3397_o}),
    .d({_al_u3397_o,_al_u6757_o}),
    .f({\cu_ru/n90 [32],\cu_ru/read_mcycle_sel_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~B*~(C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7218|cu_ru/m_cycle_event/reg0_b20  (
    .a({open_n49043,\cu_ru/read_minstret_sel_lutinv }),
    .b({\cu_ru/n90 [32],\cu_ru/n90 [32]}),
    .c({satp[35],\cu_ru/minstret [20]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/read_satp_sel_lutinv ,tvm}),
    .mi({open_n49054,\cu_ru/m_cycle_event/n4 [20]}),
    .sr(rst_pad),
    .f({_al_u7218_o,_al_u7621_o}),
    .q({open_n49058,\cu_ru/minstret [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7219|cu_ru/m_s_tval/reg0_b35  (
    .b({_al_u7218_o,_al_u5263_o}),
    .c({\cu_ru/stval [35],\cu_ru/m_s_tval/n3 [35]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/read_stval_sel_lutinv ,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7219_o,open_n49073}),
    .q({open_n49077,\cu_ru/stval [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7220|_al_u3421  (
    .b({_al_u7216_o,open_n49080}),
    .c({_al_u7219_o,_al_u3420_o}),
    .d({_al_u7215_o,_al_u3191_o}),
    .f({_al_u7220_o,\cu_ru/m_s_ip/u12_sel_is_2_o }));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7222|cu_ru/m_s_tvec/reg1_b35  (
    .b({_al_u7220_o,_al_u7223_o}),
    .c({_al_u7221_o,_al_u7224_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7214_o,_al_u7222_o}),
    .sr(rst_pad),
    .f({_al_u7222_o,csr_data[35]}),
    .q({open_n49122,\cu_ru/mtvec [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7224|cu_ru/m_s_epc/reg0_b35  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n49123}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [35],_al_u5493_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [35],\cu_ru/m_s_epc/n2 [35]}),
    .sr(rst_pad),
    .f({_al_u7224_o,open_n49140}),
    .q({open_n49144,\cu_ru/sepc [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7226|cu_ru/m_s_cause/reg0_b34  (
    .a({open_n49145,_al_u5157_o}),
    .b({\cu_ru/n90 [32],\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [34],\cu_ru/scause [34]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/read_scause_sel_lutinv ,data_csr[34]}),
    .sr(rst_pad),
    .f({_al_u7226_o,open_n49162}),
    .q({open_n49166,\cu_ru/scause [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7227|cu_ru/m_s_tval/reg1_b34  (
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [34],\cu_ru/m_s_tval/n3 [34]}),
    .clk(clk_pad),
    .d({_al_u7226_o,_al_u6513_o}),
    .sr(rst_pad),
    .f({_al_u7227_o,open_n49186}),
    .q({open_n49190,\cu_ru/mtval [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7228|cu_ru/m_s_scratch/reg0_b34  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n49191}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [34]}),
    .c({\cu_ru/mscratch [34],data_csr[34]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [34],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n49202,data_csr[34]}),
    .sr(rst_pad),
    .f({_al_u7228_o,_al_u5497_o}),
    .q({open_n49206,\cu_ru/mscratch [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u7229|cu_ru/m_s_cause/reg1_b34  (
    .a({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({satp[34],\cu_ru/mtval [34]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [34],data_csr[34]}),
    .mi({open_n49217,data_csr[34]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u7229_o,_al_u6513_o}),
    .q({open_n49221,\cu_ru/mcause [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u7232|_al_u7504  (
    .a({\cu_ru/read_time_sel_lutinv ,\cu_ru/read_time_sel_lutinv }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_stvec_sel_lutinv }),
    .c({mtime_pad[34],mtime_pad[7]}),
    .d({\cu_ru/stvec [34],\cu_ru/stvec [7]}),
    .f({_al_u7232_o,_al_u7504_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7233|cu_ru/m_s_tvec/reg1_b34  (
    .b({_al_u7231_o,_al_u7234_o}),
    .c({_al_u7232_o,_al_u7235_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7230_o,_al_u7233_o}),
    .sr(rst_pad),
    .f({_al_u7233_o,csr_data[34]}),
    .q({open_n49263,\cu_ru/mtvec [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7235|cu_ru/m_s_tval/reg0_b34  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n49264}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5266_o}),
    .c({\cu_ru/stval [34],\cu_ru/m_s_tval/n3 [34]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [34],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7235_o,open_n49277}),
    .q({open_n49281,\cu_ru/stval [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u7239|_al_u7238  (
    .a({open_n49282,_al_u3400_o}),
    .b({open_n49283,id_ins[31]}),
    .c({id_ins[20],id_ins[30]}),
    .d({_al_u7238_o,id_ins[29]}),
    .f({_al_u7239_o,_al_u7238_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7241|_al_u2681  (
    .b({_al_u7240_o,open_n49306}),
    .c({_al_u3394_o,\ins_fetch/ins_hold [22]}),
    .d({_al_u7239_o,1'b0}),
    .f({\cu_ru/n82 [14],_al_u2681_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7242|cu_ru/m_s_scratch/reg0_b25  (
    .a({_al_u7237_o,open_n49327}),
    .b({\cu_ru/n82 [14],\cu_ru/sepc [25]}),
    .c({\cu_ru/read_mscratch_sel_lutinv ,data_csr[25]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [25],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n49338,data_csr[25]}),
    .sr(rst_pad),
    .f({_al_u7242_o,_al_u5537_o}),
    .q({open_n49342,\cu_ru/mscratch [25]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7243|cu_ru/m_s_cause/reg0_b25  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({satp[25],\cu_ru/scause [25]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [25],data_csr[25]}),
    .sr(rst_pad),
    .f({_al_u7243_o,open_n49359}),
    .q({open_n49363,\cu_ru/scause [25]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7244|cu_ru/m_s_epc/reg0_b25  (
    .a({_al_u7242_o,open_n49364}),
    .b({_al_u7243_o,_al_u5157_o}),
    .c({\cu_ru/read_sepc_sel_lutinv ,_al_u5537_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [25],\cu_ru/m_s_epc/n2 [25]}),
    .sr(rst_pad),
    .f({_al_u7244_o,open_n49381}),
    .q({open_n49385,\cu_ru/sepc [25]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7246|cu_ru/m_s_tval/reg0_b25  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n49386}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5296_o}),
    .c({\cu_ru/stval [25],\cu_ru/m_s_tval/n3 [25]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [25],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7246_o,open_n49403}),
    .q({open_n49407,\cu_ru/stval [25]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*~A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*~A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010101000111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0010101000111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7247|cu_ru/m_cycle_event/reg0_b25  (
    .a({open_n49408,_al_u6763_o}),
    .b({_al_u7245_o,\cu_ru/read_time_sel_lutinv }),
    .c({_al_u7246_o,mtime_pad[25]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7244_o,\cu_ru/minstret [25]}),
    .mi({open_n49412,\cu_ru/m_cycle_event/n4 [25]}),
    .sr(rst_pad),
    .f({_al_u7247_o,_al_u7245_o}),
    .q({open_n49427,\cu_ru/minstret [25]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7248|cu_ru/m_s_tval/reg1_b25  (
    .a({_al_u6788_o,open_n49428}),
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [25],\cu_ru/m_s_tval/n3 [25]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [25],_al_u6533_o}),
    .sr(rst_pad),
    .f({_al_u7248_o,open_n49442}),
    .q({open_n49446,\cu_ru/mtval [25]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*B*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(C*B*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111111111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0011111111111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7249|cu_ru/m_s_tvec/reg1_b25  (
    .a({\cu_ru/read_mepc_sel_lutinv ,open_n49447}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u7248_o}),
    .c({\cu_ru/mepc [25],_al_u7249_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [25],_al_u7247_o}),
    .sr(rst_pad),
    .f({_al_u7249_o,csr_data[25]}),
    .q({open_n49467,\cu_ru/mtvec [25]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7252|cu_ru/m_s_epc/reg0_b21  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n49468}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [21],_al_u5553_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [21],\cu_ru/m_s_epc/n2 [21]}),
    .sr(rst_pad),
    .f({_al_u7252_o,open_n49485}),
    .q({open_n49489,\cu_ru/sepc [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7253|cu_ru/m_s_tval/reg0_b21  (
    .a({_al_u7251_o,open_n49490}),
    .b({_al_u7252_o,_al_u5308_o}),
    .c({\cu_ru/read_stval_sel_lutinv ,\cu_ru/m_s_tval/n3 [21]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [21],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7253_o,open_n49507}),
    .q({open_n49511,\cu_ru/stval [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7256|cu_ru/m_s_scratch/reg1_b21  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n49512}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/stval [21]}),
    .c({satp[21],data_csr[21]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [21],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n49516,data_csr[21]}),
    .sr(rst_pad),
    .f({_al_u7256_o,_al_u5308_o}),
    .q({open_n49531,\cu_ru/sscratch [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7257|cu_ru/m_s_cause/reg0_b21  (
    .a({\cu_ru/read_mcause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [21],\cu_ru/scause [21]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [21],data_csr[21]}),
    .sr(rst_pad),
    .f({_al_u7257_o,open_n49548}),
    .q({open_n49552,\cu_ru/scause [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7258|cu_ru/m_cycle_event/reg0_b21  (
    .a({_al_u7254_o,\cu_ru/read_minstret_sel_lutinv }),
    .b({_al_u7255_o,\cu_ru/read_mscratch_sel_lutinv }),
    .c({_al_u7256_o,\cu_ru/minstret [21]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7257_o,\cu_ru/mscratch [21]}),
    .mi({open_n49563,\cu_ru/m_cycle_event/n4 [21]}),
    .sr(rst_pad),
    .f({_al_u7258_o,_al_u7254_o}),
    .q({open_n49567,\cu_ru/minstret [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7259|cu_ru/m_s_tvec/reg1_b21  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,_al_u7253_o}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u7258_o}),
    .c({\cu_ru/mepc [21],_al_u7259_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [21],_al_u7260_o}),
    .sr(rst_pad),
    .f({_al_u7259_o,csr_data[21]}),
    .q({open_n49583,\cu_ru/mtvec [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7260|_al_u7456  (
    .a({\cu_ru/read_time_sel_lutinv ,\cu_ru/read_time_sel_lutinv }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_stvec_sel_lutinv }),
    .c({mtime_pad[21],mtime_pad[19]}),
    .d({\cu_ru/stvec [21],\cu_ru/stvec [19]}),
    .f({_al_u7260_o,_al_u7456_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7262|cu_ru/m_s_cause/reg0_b15  (
    .a({\cu_ru/read_mcause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [15],\cu_ru/scause [15]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [15],data_csr[15]}),
    .sr(rst_pad),
    .f({_al_u7262_o,open_n49624}),
    .q({open_n49628,\cu_ru/scause [15]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7263|cu_ru/m_s_tval/reg1_b15  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n49629}),
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({mtime_pad[15],\cu_ru/m_s_tval/n3 [15]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [15],_al_u6555_o}),
    .sr(rst_pad),
    .f({_al_u7263_o,open_n49647}),
    .q({open_n49651,\cu_ru/mtval [15]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7264|cu_ru/m_s_tvec/reg1_b15  (
    .a({_al_u7262_o,_al_u7264_o}),
    .b({_al_u7263_o,_al_u7270_o}),
    .c({\cu_ru/read_mepc_sel_lutinv ,_al_u7271_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [15],_al_u7272_o}),
    .sr(rst_pad),
    .f({_al_u7264_o,csr_data[15]}),
    .q({open_n49667,\cu_ru/mtvec [15]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*~(D*A)))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~(~B*~(D*A)))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1110000011000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1110000011000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7265|_al_u7718  (
    .a({open_n49668,_al_u7478_o}),
    .b({open_n49669,_al_u7717_o}),
    .c({_al_u6791_o,_al_u6791_o}),
    .d({_al_u6758_o,\cu_ru/mie }),
    .f({\cu_ru/read_medeleg_sel_lutinv ,_al_u7718_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7267|cu_ru/m_s_scratch/reg0_b15  (
    .a({\cu_ru/read_instret_sel_lutinv ,open_n49694}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [15]}),
    .c({\cu_ru/minstret [15],data_csr[15]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [15],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n49698,data_csr[15]}),
    .sr(rst_pad),
    .f({_al_u7267_o,_al_u5581_o}),
    .q({open_n49713,\cu_ru/mscratch [15]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7270|cu_ru/m_cycle_event/reg0_b15  (
    .a({_al_u7266_o,\cu_ru/read_minstret_sel_lutinv }),
    .b({_al_u7267_o,\cu_ru/read_satp_sel_lutinv }),
    .c({_al_u7268_o,satp[15]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7269_o,\cu_ru/minstret [15]}),
    .mi({open_n49724,\cu_ru/m_cycle_event/n4 [15]}),
    .sr(rst_pad),
    .f({_al_u7270_o,_al_u7268_o}),
    .q({open_n49728,\cu_ru/minstret [15]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7271|cu_ru/m_s_epc/reg0_b15  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n49729}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [15],_al_u5581_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [15],\cu_ru/m_s_epc/n2 [15]}),
    .sr(rst_pad),
    .f({_al_u7271_o,open_n49746}),
    .q({open_n49750,\cu_ru/sepc [15]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7272|cu_ru/m_s_tval/reg0_b15  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n49751}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u5329_o}),
    .c({\cu_ru/stval [15],\cu_ru/m_s_tval/n3 [15]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [15],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7272_o,open_n49768}),
    .q({open_n49772,\cu_ru/stval [15]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7274|cu_ru/m_s_cause/reg0_b13  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [13],\cu_ru/scause [13]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [13],data_csr[13]}),
    .sr(rst_pad),
    .f({_al_u7274_o,open_n49789}),
    .q({open_n49793,\cu_ru/scause [13]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7276|biu/bus_unit/mmu/reg2_b25  (
    .a({\cu_ru/read_medeleg_sel_lutinv ,open_n49794}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n49795}),
    .c({satp[13],_al_u3134_o}),
    .clk(clk_pad),
    .d({\cu_ru/medeleg [13],_al_u3133_o}),
    .sr(rst_pad),
    .f({_al_u7276_o,open_n49809}),
    .q({open_n49813,\biu/paddress [89]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7277|cu_ru/m_s_scratch/reg0_b13  (
    .a({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcause [13],\cu_ru/mtval [13]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [13],data_csr[13]}),
    .mi({open_n49817,data_csr[13]}),
    .sr(rst_pad),
    .f({_al_u7277_o,_al_u6559_o}),
    .q({open_n49832,\cu_ru/mscratch [13]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7278|_al_u7275  (
    .b({_al_u7276_o,_al_u7274_o}),
    .c({_al_u7277_o,\cu_ru/mcycle [13]}),
    .d({_al_u7275_o,_al_u6788_o}),
    .f({_al_u7278_o,_al_u7275_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7280|cu_ru/m_s_tval/reg1_b13  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n49855}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [13],\cu_ru/m_s_tval/n3 [13]}),
    .clk(clk_pad),
    .d({\cu_ru/stvec [13],_al_u6559_o}),
    .sr(rst_pad),
    .f({_al_u7280_o,open_n49869}),
    .q({open_n49873,\cu_ru/mtval [13]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7281|cu_ru/m_cycle_event/reg0_b13  (
    .a({open_n49874,_al_u6763_o}),
    .b({_al_u7279_o,\cu_ru/read_mepc_sel_lutinv }),
    .c({_al_u7280_o,\cu_ru/minstret [13]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7278_o,\cu_ru/mepc [13]}),
    .mi({open_n49878,\cu_ru/m_cycle_event/n4 [13]}),
    .sr(rst_pad),
    .f({_al_u7281_o,_al_u7279_o}),
    .q({open_n49893,\cu_ru/minstret [13]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7282|cu_ru/m_s_epc/reg0_b13  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n49894}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({mtime_pad[13],_al_u5589_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [13],\cu_ru/m_s_epc/n2 [13]}),
    .sr(rst_pad),
    .f({_al_u7282_o,open_n49911}),
    .q({open_n49915,\cu_ru/sepc [13]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7283|cu_ru/m_s_tval/reg0_b13  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n49916}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5335_o}),
    .c({\cu_ru/stval [13],\cu_ru/m_s_tval/n3 [13]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [13],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7283_o,open_n49929}),
    .q({open_n49933,\cu_ru/stval [13]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~B*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*C*~B*A)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7286|_al_u7285  (
    .a({open_n49934,_al_u7240_o}),
    .b({open_n49935,id_ins[22]}),
    .c({_al_u7285_o,id_ins[21]}),
    .d({_al_u7238_o,id_ins[20]}),
    .f({\cu_ru/n84 [10],_al_u7285_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~B*~(C*D))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7287|cu_ru/m_s_cause/reg0_b10  (
    .a({open_n49960,_al_u5157_o}),
    .b({\cu_ru/n84 [10],\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [10],\cu_ru/scause [10]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/read_scause_sel_lutinv ,data_csr[10]}),
    .sr(rst_pad),
    .f({_al_u7287_o,open_n49977}),
    .q({open_n49981,\cu_ru/scause [10]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7289|cu_ru/m_s_tvec/reg1_b10  (
    .a({_al_u7287_o,_al_u7289_o}),
    .b({_al_u7288_o,_al_u7294_o}),
    .c({\cu_ru/read_stvec_sel_lutinv ,_al_u7295_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [10],_al_u7296_o}),
    .sr(rst_pad),
    .f({_al_u7289_o,csr_data[10]}),
    .q({open_n49997,\cu_ru/mtvec [10]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7290|cu_ru/m_s_scratch/reg0_b10  (
    .a({\cu_ru/read_instret_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/minstret [10],\cu_ru/mtval [10]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [10],data_csr[10]}),
    .mi({open_n50001,data_csr[10]}),
    .sr(rst_pad),
    .f({_al_u7290_o,_al_u6565_o}),
    .q({open_n50016,\cu_ru/mscratch [10]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u7291|_al_u7439  (
    .a({\cu_ru/read_cycle_sel_lutinv ,\cu_ru/read_cycle_sel_lutinv }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/read_mcause_sel_lutinv }),
    .c({\cu_ru/mcycle [10],\cu_ru/mcycle [28]}),
    .d({\cu_ru/mcause [10],\cu_ru/mcause [28]}),
    .f({_al_u7291_o,_al_u7439_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7293|cu_ru/m_s_scratch/reg1_b10  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n50037}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/sepc [10]}),
    .c({satp[10],data_csr[10]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [10],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n50041,data_csr[10]}),
    .sr(rst_pad),
    .f({_al_u7293_o,_al_u5601_o}),
    .q({open_n50056,\cu_ru/sscratch [10]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7294|cu_ru/m_cycle_event/reg0_b10  (
    .a({_al_u7290_o,\cu_ru/read_mcycle_sel_lutinv }),
    .b({_al_u7291_o,\cu_ru/read_minstret_sel_lutinv }),
    .c({_al_u7292_o,\cu_ru/minstret [10]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7293_o,\cu_ru/mcycle [10]}),
    .mi({open_n50067,\cu_ru/m_cycle_event/n4 [10]}),
    .sr(rst_pad),
    .f({_al_u7294_o,_al_u7292_o}),
    .q({open_n50071,\cu_ru/minstret [10]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7295|cu_ru/m_s_epc/reg0_b10  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n50072}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [10],_al_u5601_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [10],\cu_ru/m_s_epc/n2 [10]}),
    .sr(rst_pad),
    .f({_al_u7295_o,open_n50089}),
    .q({open_n50093,\cu_ru/sepc [10]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7296|biu/bus_unit/mmu/reg2_b22  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n50094}),
    .b({\cu_ru/read_mepc_sel_lutinv ,open_n50095}),
    .c({\cu_ru/mepc [10],_al_u3143_o}),
    .clk(clk_pad),
    .d({\cu_ru/stval [10],_al_u3142_o}),
    .sr(rst_pad),
    .f({_al_u7296_o,open_n50109}),
    .q({open_n50113,\biu/paddress [86]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*D))"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b1111110011001100),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u7330|_al_u2708  (
    .b({\biu/bus_unit/mmu/n45_lutinv ,_al_u2706_o}),
    .c({hresp_pad,_al_u2707_o}),
    .d({_al_u2707_o,_al_u2705_o}),
    .f({_al_u7330_o,hwrite_pad}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7331|_al_u5981  (
    .b({\biu/bus_unit/mmu/statu [2],open_n50138}),
    .c({\biu/bus_unit/mmu/statu [3],_al_u5980_o}),
    .d({_al_u7330_o,_al_u2915_o}),
    .f({_al_u7331_o,_al_u5981_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7332|_al_u7487  (
    .b({open_n50165,\biu/bus_unit/mmu/n39 [0]}),
    .c({\biu/bus_unit/mmu_hwdata [6],\biu/bus_unit/mmu_hwdata [6]}),
    .d({\biu/bus_unit/mmu/n39 [0],\biu/bus_unit/mmu/n37_lutinv }),
    .f({\biu/bus_unit/mmu/n40 [2],_al_u7487_o}));
  // ../../RTL/CPU/BIU/mmu.v(154)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*D)"),
    //.LUTF1("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTG0("~(~C*D)"),
    //.LUTG1("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b1010100010101100),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b1010100010101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7333|biu/bus_unit/mmu/reg4_b2  (
    .a({_al_u7203_o,open_n50190}),
    .b({_al_u7331_o,open_n50191}),
    .c({_al_u2915_o,_al_u2963_o}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu/n40 [2],_al_u7333_o}),
    .sr(rst_pad),
    .f({_al_u7333_o,open_n50209}),
    .q({open_n50213,\biu/bus_unit/mmu/statu [2]}));  // ../../RTL/CPU/BIU/mmu.v(154)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7340|cu_ru/m_s_tval/reg0_b6  (
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5182_o}),
    .c({\cu_ru/stval [6],\cu_ru/m_s_tval/n3 [6]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u7339_o,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7340_o,open_n50228}),
    .q({open_n50232,\cu_ru/stval [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7342|cu_ru/m_s_scratch/reg0_b6  (
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [6]}),
    .c({\cu_ru/mscratch [6],data_csr[6]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({_al_u7341_o,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n50238,data_csr[6]}),
    .sr(rst_pad),
    .f({_al_u7342_o,_al_u5385_o}),
    .q({open_n50253,\cu_ru/mscratch [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7343|biu/bus_unit/mmu/reg2_b18  (
    .a({\cu_ru/read_mcause_sel_lutinv ,open_n50254}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n50255}),
    .c({satp[6],_al_u3156_o}),
    .clk(clk_pad),
    .d({\cu_ru/mcause [6],_al_u3155_o}),
    .sr(rst_pad),
    .f({_al_u7343_o,open_n50269}),
    .q({open_n50273,\biu/paddress [82]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7344|cu_ru/m_s_cause/reg0_b6  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/mcycle [6],\cu_ru/scause [6]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [6],data_csr[6]}),
    .sr(rst_pad),
    .f({_al_u7344_o,open_n50290}),
    .q({open_n50294,\cu_ru/scause [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7345|cu_ru/m_s_tvec/reg1_b6  (
    .a({_al_u7340_o,_al_u7345_o}),
    .b({_al_u7342_o,_al_u7347_o}),
    .c({_al_u7343_o,_al_u7348_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7344_o,_al_u7349_o}),
    .sr(rst_pad),
    .f({_al_u7345_o,csr_data[6]}),
    .q({open_n50310,\cu_ru/mtvec [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7346|cu_ru/m_s_tval/reg1_b6  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n50311}),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [6],\cu_ru/m_s_tval/n3 [6]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [6],_al_u6447_o}),
    .sr(rst_pad),
    .f({_al_u7346_o,open_n50329}),
    .q({open_n50333,\cu_ru/mtval [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u7347|_al_u7443  (
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/stvec [6],\cu_ru/stvec [28]}),
    .d({_al_u7346_o,_al_u7442_o}),
    .f({_al_u7347_o,_al_u7443_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7349|cu_ru/m_s_epc/reg0_b6  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n50356}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({mtime_pad[6],_al_u5385_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [6],\cu_ru/m_s_epc/n2 [6]}),
    .sr(rst_pad),
    .f({_al_u7349_o,open_n50373}),
    .q({open_n50377,\cu_ru/sepc [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7352|cu_ru/m_s_tvec/reg0_b59  (
    .a({_al_u7351_o,csr_data[59]}),
    .b({rs1_data[59],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[59]}),
    .mi({open_n50381,csr_data[59]}),
    .sr(rst_pad),
    .f({_al_u7352_o,_al_u7351_o}),
    .q({open_n50396,\cu_ru/stvec [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b0000000010101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7356|cu_ru/m_s_tvec/reg0_b58  (
    .a({_al_u7355_o,csr_data[58]}),
    .b({rs1_data[58],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[58]}),
    .mi({open_n50407,csr_data[58]}),
    .sr(rst_pad),
    .f({_al_u7356_o,_al_u7355_o}),
    .q({open_n50411,\cu_ru/stvec [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b0000000010101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7359|cu_ru/m_s_tvec/reg0_b57  (
    .a({_al_u7358_o,csr_data[57]}),
    .b({rs1_data[57],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[57]}),
    .mi({open_n50422,csr_data[57]}),
    .sr(rst_pad),
    .f({_al_u7359_o,_al_u7358_o}),
    .q({open_n50426,\cu_ru/stvec [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7362|cu_ru/m_s_tvec/reg0_b56  (
    .a({_al_u7361_o,csr_data[56]}),
    .b({rs1_data[56],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[56]}),
    .mi({open_n50430,csr_data[56]}),
    .sr(rst_pad),
    .f({_al_u7362_o,_al_u7361_o}),
    .q({open_n50445,\cu_ru/stvec [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7365|cu_ru/m_s_tvec/reg0_b55  (
    .a({_al_u7364_o,csr_data[55]}),
    .b({rs1_data[55],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[55]}),
    .mi({open_n50449,csr_data[55]}),
    .sr(rst_pad),
    .f({_al_u7365_o,_al_u7364_o}),
    .q({open_n50464,\cu_ru/stvec [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b0000000010101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7368|cu_ru/m_s_tvec/reg0_b54  (
    .a({_al_u7367_o,csr_data[54]}),
    .b({rs1_data[54],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[54]}),
    .mi({open_n50475,csr_data[54]}),
    .sr(rst_pad),
    .f({_al_u7368_o,_al_u7367_o}),
    .q({open_n50479,\cu_ru/stvec [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b0000000010101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7371|cu_ru/m_s_tvec/reg0_b53  (
    .a({_al_u7370_o,csr_data[53]}),
    .b({rs1_data[53],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[53]}),
    .mi({open_n50490,csr_data[53]}),
    .sr(rst_pad),
    .f({_al_u7371_o,_al_u7370_o}),
    .q({open_n50494,\cu_ru/stvec [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7374|cu_ru/m_s_tvec/reg0_b52  (
    .a({_al_u7373_o,csr_data[52]}),
    .b({rs1_data[52],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[52]}),
    .mi({open_n50498,csr_data[52]}),
    .sr(rst_pad),
    .f({_al_u7374_o,_al_u7373_o}),
    .q({open_n50513,\cu_ru/stvec [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7377|cu_ru/m_s_tvec/reg0_b51  (
    .a({_al_u7376_o,csr_data[51]}),
    .b({rs1_data[51],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[51]}),
    .mi({open_n50517,csr_data[51]}),
    .sr(rst_pad),
    .f({_al_u7377_o,_al_u7376_o}),
    .q({open_n50532,\cu_ru/stvec [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b0000000010101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7380|cu_ru/m_s_tvec/reg0_b50  (
    .a({_al_u7379_o,csr_data[50]}),
    .b({rs1_data[50],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[50]}),
    .mi({open_n50543,csr_data[50]}),
    .sr(rst_pad),
    .f({_al_u7380_o,_al_u7379_o}),
    .q({open_n50547,\cu_ru/stvec [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7383|cu_ru/m_s_tvec/reg0_b49  (
    .a({_al_u7382_o,csr_data[49]}),
    .b({rs1_data[49],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[49]}),
    .mi({open_n50551,csr_data[49]}),
    .sr(rst_pad),
    .f({_al_u7383_o,_al_u7382_o}),
    .q({open_n50566,\cu_ru/stvec [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7386|cu_ru/m_s_tvec/reg0_b48  (
    .a({_al_u7385_o,csr_data[48]}),
    .b({rs1_data[48],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[48]}),
    .mi({open_n50570,csr_data[48]}),
    .sr(rst_pad),
    .f({_al_u7386_o,_al_u7385_o}),
    .q({open_n50585,\cu_ru/stvec [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b0000000010101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7389|cu_ru/m_s_tvec/reg0_b47  (
    .a({_al_u7388_o,csr_data[47]}),
    .b({rs1_data[47],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[47]}),
    .mi({open_n50596,csr_data[47]}),
    .sr(rst_pad),
    .f({_al_u7389_o,_al_u7388_o}),
    .q({open_n50600,\cu_ru/stvec [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010000000),
    .INIT_LUT1(16'b0000000010101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7392|cu_ru/m_s_tvec/reg0_b46  (
    .a({_al_u7391_o,csr_data[46]}),
    .b({rs1_data[46],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[46]}),
    .mi({open_n50611,csr_data[46]}),
    .sr(rst_pad),
    .f({_al_u7392_o,_al_u7391_o}),
    .q({open_n50615,\cu_ru/stvec [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7395|cu_ru/m_s_tvec/reg0_b45  (
    .a({_al_u7394_o,csr_data[45]}),
    .b({rs1_data[45],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[45]}),
    .mi({open_n50619,csr_data[45]}),
    .sr(rst_pad),
    .f({_al_u7395_o,_al_u7394_o}),
    .q({open_n50634,\cu_ru/stvec [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7398|cu_ru/m_s_tvec/reg0_b44  (
    .a({_al_u7397_o,csr_data[44]}),
    .b({rs1_data[44],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[44]}),
    .mi({open_n50638,csr_data[44]}),
    .sr(rst_pad),
    .f({_al_u7398_o,_al_u7397_o}),
    .q({open_n50653,\cu_ru/stvec [44]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u7400|_al_u6777  (
    .c({_al_u3397_o,_al_u3400_o}),
    .d({_al_u6777_o,_al_u3399_o}),
    .f({\cu_ru/n64 [32],_al_u6777_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u7401|_al_u7483  (
    .a({open_n50678,\cu_ru/read_mcause_sel_lutinv }),
    .b({open_n50679,\cu_ru/n90 [32]}),
    .c({\cu_ru/n90 [32],\cu_ru/mcause [11]}),
    .d({\cu_ru/n64 [32],\cu_ru/mstatus [11]}),
    .f({_al_u7401_o,_al_u7483_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7402|cu_ru/m_s_scratch/reg1_b33  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n50700}),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/stval [33]}),
    .c({\cu_ru/mcause [33],data_csr[33]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [33],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n50711,data_csr[33]}),
    .sr(rst_pad),
    .f({_al_u7402_o,_al_u5269_o}),
    .q({open_n50715,\cu_ru/sscratch [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7403|cu_ru/m_s_cause/reg0_b33  (
    .a({_al_u7401_o,_al_u5157_o}),
    .b({_al_u7402_o,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/read_scause_sel_lutinv ,\cu_ru/scause [33]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [33],data_csr[33]}),
    .sr(rst_pad),
    .f({_al_u7403_o,open_n50732}),
    .q({open_n50736,\cu_ru/scause [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7405|cu_ru/m_s_scratch/reg0_b33  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,open_n50737}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [33]}),
    .c({\cu_ru/mcycle [33],data_csr[33]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [33],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n50748,data_csr[33]}),
    .sr(rst_pad),
    .f({_al_u7405_o,_al_u5501_o}),
    .q({open_n50752,\cu_ru/mscratch [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7406|_al_u7404  (
    .a({open_n50753,\cu_ru/read_cycle_sel_lutinv }),
    .b({_al_u7404_o,\cu_ru/read_satp_sel_lutinv }),
    .c({_al_u7405_o,satp[33]}),
    .d({_al_u7403_o,\cu_ru/mcycle [33]}),
    .f({_al_u7406_o,_al_u7404_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7408|cu_ru/m_s_epc/reg0_b33  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n50774}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [33],_al_u5501_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [33],\cu_ru/m_s_epc/n2 [33]}),
    .sr(rst_pad),
    .f({_al_u7408_o,open_n50791}),
    .q({open_n50795,\cu_ru/sepc [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*~A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010101000111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7409|cu_ru/m_cycle_event/reg0_b33  (
    .a({open_n50796,_al_u6763_o}),
    .b({_al_u7407_o,\cu_ru/read_time_sel_lutinv }),
    .c({_al_u7408_o,mtime_pad[33]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7406_o,\cu_ru/minstret [33]}),
    .mi({open_n50807,\cu_ru/m_cycle_event/n4 [33]}),
    .sr(rst_pad),
    .f({_al_u7409_o,_al_u7407_o}),
    .q({open_n50811,\cu_ru/minstret [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7410|cu_ru/m_s_tval/reg0_b33  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n50812}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5269_o}),
    .c({\cu_ru/mepc [33],\cu_ru/m_s_tval/n3 [33]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [33],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7410_o,open_n50829}),
    .q({open_n50833,\cu_ru/stval [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7411|cu_ru/m_s_tvec/reg1_b33  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n50834}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u7410_o}),
    .c({\cu_ru/stvec [33],_al_u7411_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [33],_al_u7409_o}),
    .sr(rst_pad),
    .f({_al_u7411_o,csr_data[33]}),
    .q({open_n50850,\cu_ru/mtvec [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7413|cu_ru/m_s_cause/reg0_b32  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [32],\cu_ru/scause [32]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [32],data_csr[32]}),
    .sr(rst_pad),
    .f({_al_u7413_o,open_n50867}),
    .q({open_n50871,\cu_ru/scause [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D*~(~C*~B)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0000001010101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u7414|_al_u6844  (
    .a({_al_u7401_o,_al_u6843_o}),
    .b({_al_u7413_o,\cu_ru/read_mcycle_sel_lutinv }),
    .c({\cu_ru/read_mcycle_sel_lutinv ,\cu_ru/read_cycle_sel_lutinv }),
    .d({\cu_ru/mcycle [32],\cu_ru/mcycle [53]}),
    .f({_al_u7414_o,_al_u6844_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7415|cu_ru/m_s_scratch/reg0_b32  (
    .a({\cu_ru/read_mcause_sel_lutinv ,open_n50892}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [32]}),
    .c({\cu_ru/mcause [32],data_csr[32]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [32],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n50896,data_csr[32]}),
    .sr(rst_pad),
    .f({_al_u7415_o,_al_u5505_o}),
    .q({open_n50911,\cu_ru/mscratch [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7417|_al_u7416  (
    .a({open_n50912,\cu_ru/read_cycle_sel_lutinv }),
    .b({_al_u7415_o,\cu_ru/read_satp_sel_lutinv }),
    .c({_al_u7416_o,satp[32]}),
    .d({_al_u7414_o,\cu_ru/mcycle [32]}),
    .f({_al_u7417_o,_al_u7416_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7420|cu_ru/m_cycle_event/reg0_b32  (
    .a({open_n50937,_al_u6763_o}),
    .b({_al_u7418_o,\cu_ru/read_mtval_sel_lutinv }),
    .c({_al_u7419_o,\cu_ru/minstret [32]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7417_o,\cu_ru/mtval [32]}),
    .mi({open_n50941,\cu_ru/m_cycle_event/n4 [32]}),
    .sr(rst_pad),
    .f({_al_u7420_o,_al_u7418_o}),
    .q({open_n50956,\cu_ru/minstret [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7421|cu_ru/m_s_epc/reg0_b32  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n50957}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [32],_al_u5505_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [32],\cu_ru/m_s_epc/n2 [32]}),
    .sr(rst_pad),
    .f({_al_u7421_o,open_n50974}),
    .q({open_n50978,\cu_ru/sepc [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7422|cu_ru/m_s_tval/reg0_b32  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n50979}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u5272_o}),
    .c({\cu_ru/stval [32],\cu_ru/m_s_tval/n3 [32]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [32],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7422_o,open_n50996}),
    .q({open_n51000,\cu_ru/stval [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7425|cu_ru/m_s_cause/reg0_b30  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [30],\cu_ru/scause [30]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [30],data_csr[30]}),
    .sr(rst_pad),
    .f({_al_u7425_o,open_n51017}),
    .q({open_n51021,\cu_ru/scause [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7426|cu_ru/m_s_tval/reg0_b30  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n51022}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5278_o}),
    .c({\cu_ru/stval [30],\cu_ru/m_s_tval/n3 [30]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [30],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7426_o,open_n51035}),
    .q({open_n51039,\cu_ru/stval [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7427|_al_u7424  (
    .a({open_n51040,\cu_ru/read_mcycle_sel_lutinv }),
    .b({_al_u7425_o,\cu_ru/read_satp_sel_lutinv }),
    .c({_al_u7426_o,satp[30]}),
    .d({_al_u7424_o,\cu_ru/mcycle [30]}),
    .f({_al_u7427_o,_al_u7424_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7428|cu_ru/m_s_scratch/reg0_b30  (
    .a({\cu_ru/read_cycle_sel_lutinv ,open_n51065}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [30]}),
    .c({\cu_ru/mcycle [30],data_csr[30]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [30],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n51076,data_csr[30]}),
    .sr(rst_pad),
    .f({_al_u7428_o,_al_u5513_o}),
    .q({open_n51080,\cu_ru/mscratch [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7429|cu_ru/m_s_tvec/reg1_b30  (
    .a({_al_u7427_o,open_n51081}),
    .b({_al_u7428_o,open_n51082}),
    .c({\cu_ru/read_mcause_sel_lutinv ,_al_u7434_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [30],_al_u7429_o}),
    .sr(rst_pad),
    .f({_al_u7429_o,csr_data[30]}),
    .q({open_n51098,\cu_ru/mtvec [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*A*~(D*B))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000001000001010),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u7430|_al_u7653  (
    .a({open_n51099,_al_u7652_o}),
    .b({open_n51100,\cu_ru/read_mcause_sel_lutinv }),
    .c({\cu_ru/n84 [10],\cu_ru/n84 [10]}),
    .d({\cu_ru/n82 [14],\cu_ru/mcause [12]}),
    .f({_al_u7430_o,_al_u7653_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7432|cu_ru/m_s_epc/reg0_b30  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n51121}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({mtime_pad[30],_al_u5513_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [30],\cu_ru/m_s_epc/n2 [30]}),
    .sr(rst_pad),
    .f({_al_u7432_o,open_n51138}),
    .q({open_n51142,\cu_ru/sepc [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7434|cu_ru/m_cycle_event/reg0_b30  (
    .a({_al_u7430_o,_al_u6763_o}),
    .b({_al_u7431_o,\cu_ru/read_mtval_sel_lutinv }),
    .c({_al_u7432_o,\cu_ru/minstret [30]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7433_o,\cu_ru/mtval [30]}),
    .mi({open_n51153,\cu_ru/m_cycle_event/n4 [30]}),
    .sr(rst_pad),
    .f({_al_u7434_o,_al_u7431_o}),
    .q({open_n51157,\cu_ru/minstret [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7436|cu_ru/m_s_epc/reg0_b28  (
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [28],_al_u5525_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u7430_o,\cu_ru/m_s_epc/n2 [28]}),
    .sr(rst_pad),
    .f({_al_u7436_o,open_n51176}),
    .q({open_n51180,\cu_ru/sepc [28]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7437|cu_ru/m_s_cause/reg0_b28  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [28],\cu_ru/scause [28]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [28],data_csr[28]}),
    .sr(rst_pad),
    .f({_al_u7437_o,open_n51197}),
    .q({open_n51201,\cu_ru/scause [28]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7440|cu_ru/m_s_scratch/reg0_b28  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,open_n51202}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [28]}),
    .c({\cu_ru/mcycle [28],data_csr[28]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [28],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n51206,data_csr[28]}),
    .sr(rst_pad),
    .f({_al_u7440_o,_al_u5525_o}),
    .q({open_n51221,\cu_ru/mscratch [28]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7441|cu_ru/m_s_tvec/reg1_b28  (
    .a({_al_u7436_o,_al_u7441_o}),
    .b({_al_u7438_o,_al_u7443_o}),
    .c({_al_u7439_o,_al_u7444_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7440_o,_al_u7445_o}),
    .sr(rst_pad),
    .f({_al_u7441_o,csr_data[28]}),
    .q({open_n51241,\cu_ru/mtvec [28]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7442|cu_ru/m_s_tval/reg0_b28  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n51242}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5287_o}),
    .c({\cu_ru/stval [28],\cu_ru/m_s_tval/n3 [28]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [28],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7442_o,open_n51255}),
    .q({open_n51259,\cu_ru/stval [28]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(~B*~(D*C)))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*~(~B*~(D*C)))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0101010001000100),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010001000100),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7447|_al_u7198  (
    .a({\cu_ru/read_cycle_sel_lutinv ,\biu/bus_unit/mmu/n19_lutinv }),
    .b({\cu_ru/n90 [32],\biu/bus_unit/mmu_hwdata [1]}),
    .c({\cu_ru/mcycle [19],\biu/bus_unit/mmu_hwdata [3]}),
    .d({mxr,mxr}),
    .f({_al_u7447_o,_al_u7198_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7448|cu_ru/m_s_scratch/reg0_b19  (
    .a({\cu_ru/read_minstret_sel_lutinv ,open_n51284}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [19]}),
    .c({\cu_ru/minstret [19],data_csr[19]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [19],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n51295,data_csr[19]}),
    .sr(rst_pad),
    .f({_al_u7448_o,_al_u5565_o}),
    .q({open_n51299,\cu_ru/mscratch [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7449|biu/bus_unit/mmu/reg2_b31  (
    .a({\cu_ru/read_mcause_sel_lutinv ,open_n51300}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n51301}),
    .c({satp[19],_al_u3116_o}),
    .clk(clk_pad),
    .d({\cu_ru/mcause [19],_al_u3115_o}),
    .sr(rst_pad),
    .f({_al_u7449_o,open_n51319}),
    .q({open_n51323,\biu/paddress [95]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7450|cu_ru/m_s_cause/reg0_b19  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/mcycle [19],\cu_ru/scause [19]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [19],data_csr[19]}),
    .sr(rst_pad),
    .f({_al_u7450_o,open_n51340}),
    .q({open_n51344,\cu_ru/scause [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7451|_al_u6752  (
    .a({_al_u7447_o,open_n51345}),
    .b({_al_u7448_o,open_n51346}),
    .c({_al_u7449_o,\cu_ru/mstatus [12]}),
    .d({_al_u7450_o,_al_u3427_o}),
    .f({_al_u7451_o,_al_u6752_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7453|cu_ru/m_s_scratch/reg1_b19  (
    .a({_al_u7451_o,open_n51371}),
    .b({_al_u7452_o,\cu_ru/stval [19]}),
    .c({\cu_ru/read_sscratch_sel_lutinv ,data_csr[19]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [19],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n51382,data_csr[19]}),
    .sr(rst_pad),
    .f({_al_u7453_o,_al_u5317_o}),
    .q({open_n51386,\cu_ru/sscratch [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7454|cu_ru/m_s_tval/reg0_b19  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n51387}),
    .b({\cu_ru/read_mtval_sel_lutinv ,_al_u5317_o}),
    .c({\cu_ru/stval [19],\cu_ru/m_s_tval/n3 [19]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [19],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7454_o,open_n51404}),
    .q({open_n51408,\cu_ru/stval [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7455|cu_ru/m_s_tvec/reg1_b19  (
    .a({open_n51409,_al_u7453_o}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u7455_o}),
    .c({\cu_ru/mepc [19],_al_u7456_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7454_o,_al_u7457_o}),
    .sr(rst_pad),
    .f({_al_u7455_o,csr_data[19]}),
    .q({open_n51429,\cu_ru/mtvec [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7457|cu_ru/m_s_epc/reg0_b19  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n51430}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [19],_al_u5565_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [19],\cu_ru/m_s_epc/n2 [19]}),
    .sr(rst_pad),
    .f({_al_u7457_o,open_n51447}),
    .q({open_n51451,\cu_ru/sepc [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7459|cu_ru/m_s_tval/reg1_b14  (
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [14],\cu_ru/m_s_tval/n3 [14]}),
    .clk(clk_pad),
    .d({_al_u7430_o,_al_u6557_o}),
    .sr(rst_pad),
    .f({_al_u7459_o,open_n51467}),
    .q({open_n51471,\cu_ru/mtval [14]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7460|biu/bus_unit/mmu/reg2_b26  (
    .a({\cu_ru/read_cycle_sel_lutinv ,open_n51472}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n51473}),
    .c({satp[14],_al_u3131_o}),
    .clk(clk_pad),
    .d({\cu_ru/mcycle [14],_al_u3130_o}),
    .sr(rst_pad),
    .f({_al_u7460_o,open_n51487}),
    .q({open_n51491,\biu/paddress [90]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7462|cu_ru/m_s_scratch/reg0_b14  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n51492}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [14]}),
    .c({\cu_ru/mscratch [14],data_csr[14]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [14],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n51503,data_csr[14]}),
    .sr(rst_pad),
    .f({_al_u7462_o,_al_u5585_o}),
    .q({open_n51507,\cu_ru/mscratch [14]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7463|cu_ru/m_s_cause/reg0_b14  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/mcycle [14],\cu_ru/scause [14]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [14],data_csr[14]}),
    .sr(rst_pad),
    .f({_al_u7463_o,open_n51524}),
    .q({open_n51528,\cu_ru/scause [14]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7464|_al_u7461  (
    .a({_al_u7459_o,open_n51529}),
    .b({_al_u7461_o,\cu_ru/read_mcause_sel_lutinv }),
    .c({_al_u7462_o,\cu_ru/mcause [14]}),
    .d({_al_u7463_o,_al_u7460_o}),
    .f({_al_u7464_o,_al_u7461_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7465|cu_ru/m_s_epc/reg0_b14  (
    .a({\cu_ru/read_sepc_sel_lutinv ,open_n51554}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [14],_al_u5585_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [14],\cu_ru/m_s_epc/n2 [14]}),
    .sr(rst_pad),
    .f({_al_u7465_o,open_n51571}),
    .q({open_n51575,\cu_ru/sepc [14]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7466|cu_ru/m_s_tval/reg0_b14  (
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5332_o}),
    .c({\cu_ru/stval [14],\cu_ru/m_s_tval/n3 [14]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u7465_o,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7466_o,open_n51594}),
    .q({open_n51598,\cu_ru/stval [14]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7468|cu_ru/m_s_tvec/reg1_b14  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,_al_u7464_o}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u7466_o}),
    .c({mtime_pad[14],_al_u7467_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [14],_al_u7468_o}),
    .sr(rst_pad),
    .f({_al_u7468_o,csr_data[14]}),
    .q({open_n51618,\cu_ru/mtvec [14]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7470|cu_ru/m_s_scratch/reg0_b11  (
    .a({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({satp[11],\cu_ru/mtval [11]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [11],data_csr[11]}),
    .mi({open_n51622,data_csr[11]}),
    .sr(rst_pad),
    .f({_al_u7470_o,_al_u6563_o}),
    .q({open_n51637,\cu_ru/mscratch [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7471|cu_ru/m_s_tval/reg0_b11  (
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5341_o}),
    .c({\cu_ru/stval [11],\cu_ru/m_s_tval/n3 [11]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u7470_o,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7471_o,open_n51656}),
    .q({open_n51660,\cu_ru/stval [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7472|cu_ru/m_cycle_event/reg0_b11  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,\cu_ru/read_instret_sel_lutinv }),
    .b({\cu_ru/read_minstret_sel_lutinv ,\cu_ru/read_scause_sel_lutinv }),
    .c({\cu_ru/minstret [11],\cu_ru/minstret [11]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcycle [11],\cu_ru/scause [11]}),
    .mi({open_n51671,\cu_ru/m_cycle_event/n4 [11]}),
    .sr(rst_pad),
    .f({_al_u7472_o,_al_u7482_o}),
    .q({open_n51675,\cu_ru/minstret [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7473|cu_ru/m_s_scratch/reg1_b11  (
    .a({\cu_ru/read_cycle_sel_lutinv ,open_n51676}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/sepc [11]}),
    .c({\cu_ru/mcycle [11],data_csr[11]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [11],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n51680,data_csr[11]}),
    .sr(rst_pad),
    .f({_al_u7473_o,_al_u5597_o}),
    .q({open_n51695,\cu_ru/sscratch [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7474|cu_ru/m_s_tvec/reg1_b11  (
    .a({open_n51696,_al_u7474_o}),
    .b({_al_u7472_o,_al_u7481_o}),
    .c({_al_u7473_o,_al_u7482_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7471_o,_al_u7483_o}),
    .sr(rst_pad),
    .f({_al_u7474_o,csr_data[11]}),
    .q({open_n51712,\cu_ru/mtvec [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7475|biu/bus_unit/mmu/reg2_b23  (
    .a({\cu_ru/read_mepc_sel_lutinv ,open_n51713}),
    .b({\cu_ru/read_stvec_sel_lutinv ,open_n51714}),
    .c({\cu_ru/mepc [11],_al_u3140_o}),
    .clk(clk_pad),
    .d({\cu_ru/stvec [11],_al_u3139_o}),
    .sr(rst_pad),
    .f({_al_u7475_o,open_n51732}),
    .q({open_n51736,\biu/paddress [87]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7476|cu_ru/m_s_tval/reg1_b11  (
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [11],\cu_ru/m_s_tval/n3 [11]}),
    .clk(clk_pad),
    .d({_al_u7475_o,_al_u6563_o}),
    .sr(rst_pad),
    .f({_al_u7476_o,open_n51756}),
    .q({open_n51760,\cu_ru/mtval [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7477|cu_ru/m_s_epc/reg0_b11  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n51761}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [11],_al_u5597_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [11],\cu_ru/m_s_epc/n2 [11]}),
    .sr(rst_pad),
    .f({_al_u7477_o,open_n51778}),
    .q({open_n51782,\cu_ru/sepc [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7479|_al_u7864  (
    .a({open_n51783,\cu_ru/read_medeleg_sel_lutinv }),
    .b({open_n51784,_al_u7863_o}),
    .c({_al_u7478_o,_al_u7478_o}),
    .d({_al_u6766_o,\cu_ru/medeleg [1]}),
    .f({\cu_ru/read_mip_sel_lutinv ,_al_u7864_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7481|_al_u7480  (
    .a({open_n51809,\cu_ru/read_time_sel_lutinv }),
    .b({_al_u7477_o,\cu_ru/read_mip_sel_lutinv }),
    .c({_al_u7480_o,mtime_pad[11]}),
    .d({_al_u7476_o,\cu_ru/m_sip [11]}),
    .f({_al_u7481_o,_al_u7480_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("~(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("~(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000111111001100),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000111111001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7486|_al_u7485  (
    .b({_al_u7485_o,\biu/bus_unit/mmu/statu [1]}),
    .c({\biu/bus_unit/mmu_hwdata [6],\biu/bus_unit/mmu/statu [3]}),
    .d({_al_u7202_o,_al_u7330_o}),
    .f({_al_u7486_o,_al_u7485_o}));
  // ../../RTL/CPU/BIU/mmu.v(154)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(~C*~D))"),
    //.LUTF1("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    //.LUTG0("~(~B*~(~C*~D))"),
    //.LUTG1("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011001111),
    .INIT_LUTF1(16'b0011001000000010),
    .INIT_LUTG0(16'b1100110011001111),
    .INIT_LUTG1(16'b0011001000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7489|biu/bus_unit/mmu/reg4_b1  (
    .a({_al_u7488_o,open_n51860}),
    .b({_al_u2697_o,_al_u2963_o}),
    .c({_al_u2964_o,_al_u2698_o}),
    .clk(clk_pad),
    .d({hresp_pad,_al_u7489_o}),
    .sr(rst_pad),
    .f({_al_u7489_o,open_n51878}),
    .q({open_n51882,\biu/bus_unit/mmu/statu [1]}));  // ../../RTL/CPU/BIU/mmu.v(154)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~C*B)*~(D*A))"),
    //.LUT1("(~D*~(~C*~B))"),
    .INIT_LUT0(16'b0101000111110011),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"))
    \_al_u7492|_al_u7491  (
    .a({open_n51883,\biu/bus_unit/mmu/mux10_b0_sel_is_2_o }),
    .b({\biu/bus_unit/mmu/statu [1],\biu/bus_unit/mmu/n45_lutinv }),
    .c({\biu/bus_unit/mmu/statu [3],hresp_pad}),
    .d({_al_u7491_o,\biu/bus_unit/mmu/statu [0]}),
    .f({_al_u7492_o,_al_u7491_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(~C*~(B*~D))"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(~C*~(B*~D))"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b0000111100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7493|_al_u7207  (
    .a({open_n51904,\biu/bus_unit/mmu/n39 [0]}),
    .b({_al_u7487_o,\biu/bus_unit/mmu/i [0]}),
    .c({_al_u2964_o,\biu/bus_unit/mmu/i [1]}),
    .d({\biu/bus_unit/mmu/n2 ,\biu/bus_unit/mmu_hwdata [2]}),
    .f({_al_u7493_o,\biu/bus_unit/mmu/n2 }));
  // ../../RTL/CPU/BIU/mmu.v(154)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(C*~B)*~(~D*~A))"),
    //.LUTF1("(C*~(~D*~(~B*~A)))"),
    //.LUTG0("~(~(C*~B)*~(~D*~A))"),
    //.LUTG1("(C*~(~D*~(~B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000001110101),
    .INIT_LUTF1(16'b1111000000010000),
    .INIT_LUTG0(16'b0011000001110101),
    .INIT_LUTG1(16'b1111000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7494|biu/bus_unit/mmu/reg4_b0  (
    .a({_al_u7202_o,_al_u7494_o}),
    .b({_al_u7492_o,_al_u2914_o}),
    .c({_al_u7493_o,_al_u2698_o}),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu/n37_lutinv ,_al_u7495_o}),
    .sr(rst_pad),
    .f({_al_u7494_o,open_n51946}),
    .q({open_n51950,\biu/bus_unit/mmu/statu [0]}));  // ../../RTL/CPU/BIU/mmu.v(154)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7499|cu_ru/m_cycle_event/reg0_b7  (
    .a({\cu_ru/read_minstret_sel_lutinv ,_al_u7501_o}),
    .b({\cu_ru/read_mcause_sel_lutinv ,_al_u7502_o}),
    .c({\cu_ru/minstret [7],\cu_ru/read_instret_sel_lutinv }),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [7],\cu_ru/minstret [7]}),
    .mi({open_n51961,\cu_ru/m_cycle_event/n4 [7]}),
    .sr(rst_pad),
    .f({_al_u7499_o,_al_u7503_o}),
    .q({open_n51965,\cu_ru/minstret [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7500|biu/bus_unit/mmu/reg2_b19  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,open_n51966}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n51967}),
    .c({satp[7],_al_u3153_o}),
    .clk(clk_pad),
    .d({\cu_ru/mcycle [7],_al_u3152_o}),
    .sr(rst_pad),
    .f({_al_u7500_o,open_n51985}),
    .q({open_n51989,\biu/paddress [83]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7501|cu_ru/m_s_scratch/reg1_b7  (
    .a({_al_u7497_o,\cu_ru/read_sscratch_sel_lutinv }),
    .b({_al_u7498_o,\cu_ru/read_mscratch_sel_lutinv }),
    .c({_al_u7499_o,\cu_ru/mscratch [7]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7500_o,\cu_ru/sscratch [7]}),
    .mi({open_n52000,data_csr[7]}),
    .sr(rst_pad),
    .f({_al_u7501_o,_al_u7498_o}),
    .q({open_n52004,\cu_ru/sscratch [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7505|cu_ru/m_s_tval/reg1_b7  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n52005}),
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [7],\cu_ru/m_s_tval/n3 [7]}),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [7],_al_u6445_o}),
    .sr(rst_pad),
    .f({_al_u7505_o,open_n52019}),
    .q({open_n52023,\cu_ru/mtval [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7506|cu_ru/m_s_epc/reg0_b7  (
    .a({\cu_ru/read_sepc_sel_lutinv ,open_n52024}),
    .b({\cu_ru/read_mip_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [7],_al_u5365_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_sip [7],\cu_ru/m_s_epc/n2 [7]}),
    .sr(rst_pad),
    .f({_al_u7506_o,open_n52041}),
    .q({open_n52045,\cu_ru/sepc [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7507|cu_ru/m_s_tval/reg0_b7  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n52046}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5167_o}),
    .c({\cu_ru/mepc [7],\cu_ru/m_s_tval/n3 [7]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [7],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7507_o,open_n52059}),
    .q({open_n52063,\cu_ru/stval [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7508|cu_ru/m_s_tvec/reg1_b7  (
    .a({_al_u7504_o,open_n52064}),
    .b({_al_u7505_o,open_n52065}),
    .c({_al_u7506_o,_al_u7508_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7507_o,_al_u7503_o}),
    .sr(rst_pad),
    .f({_al_u7508_o,csr_data[7]}),
    .q({open_n52085,\cu_ru/mtvec [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D*~A)))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~B*~(C*~(D*~A)))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001100000011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001001100000011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7510|cu_ru/m_s_tvec/reg0_b63  (
    .a({open_n52086,csr_data[63]}),
    .b({open_n52087,_al_u7510_o}),
    .c({_al_u7141_o,_al_u7511_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[63],id_system}),
    .mi({open_n52091,csr_data[63]}),
    .sr(rst_pad),
    .f({_al_u7510_o,_al_u7512_o}),
    .q({open_n52106,\cu_ru/stvec [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D*~A)))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001100000011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7514|cu_ru/m_s_tvec/reg0_b62  (
    .a({open_n52107,csr_data[62]}),
    .b({open_n52108,_al_u7514_o}),
    .c({_al_u7141_o,_al_u7515_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[62],id_system}),
    .mi({open_n52119,csr_data[62]}),
    .sr(rst_pad),
    .f({_al_u7514_o,_al_u7516_o}),
    .q({open_n52123,\cu_ru/stvec [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D*~A)))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001100000011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7518|cu_ru/m_s_tvec/reg0_b61  (
    .a({open_n52124,csr_data[61]}),
    .b({open_n52125,_al_u7518_o}),
    .c({_al_u7141_o,_al_u7519_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[61],id_system}),
    .mi({open_n52136,csr_data[61]}),
    .sr(rst_pad),
    .f({_al_u7518_o,_al_u7520_o}),
    .q({open_n52140,\cu_ru/stvec [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D*~A)))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~B*~(C*~(D*~A)))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001100000011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001001100000011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7522|cu_ru/m_s_tvec/reg0_b60  (
    .a({open_n52141,csr_data[60]}),
    .b({open_n52142,_al_u7522_o}),
    .c({_al_u7141_o,_al_u7523_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[60],id_system}),
    .mi({open_n52146,csr_data[60]}),
    .sr(rst_pad),
    .f({_al_u7522_o,_al_u7524_o}),
    .q({open_n52161,\cu_ru/stvec [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D*~A)))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~B*~(C*~(D*~A)))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001100000011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001001100000011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7526|cu_ru/m_s_tvec/reg0_b43  (
    .a({open_n52162,csr_data[43]}),
    .b({open_n52163,_al_u7526_o}),
    .c({_al_u7141_o,_al_u7527_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[43],id_system}),
    .mi({open_n52167,csr_data[43]}),
    .sr(rst_pad),
    .f({_al_u7526_o,_al_u7528_o}),
    .q({open_n52182,\cu_ru/stvec [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7531|ins_dec/reg5_b42  (
    .a({open_n52183,_al_u7530_o}),
    .b({open_n52184,_al_u7531_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[42],id_ins[31]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7531_o,open_n52201}),
    .q({open_n52205,ds1[42]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D*~A)))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001100000011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7533|cu_ru/m_s_tvec/reg0_b41  (
    .a({open_n52206,csr_data[41]}),
    .b({open_n52207,_al_u7533_o}),
    .c({_al_u7141_o,_al_u7534_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[41],id_system}),
    .mi({open_n52218,csr_data[41]}),
    .sr(rst_pad),
    .f({_al_u7533_o,_al_u7535_o}),
    .q({open_n52222,\cu_ru/stvec [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D*~A)))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001100000011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7537|cu_ru/m_s_tvec/reg0_b40  (
    .a({open_n52223,csr_data[40]}),
    .b({open_n52224,_al_u7537_o}),
    .c({_al_u7141_o,_al_u7538_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[40],id_system}),
    .mi({open_n52235,csr_data[40]}),
    .sr(rst_pad),
    .f({_al_u7537_o,_al_u7539_o}),
    .q({open_n52239,\cu_ru/stvec [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7541|cu_ru/m_cycle_event/reg0_b4  (
    .a({\cu_ru/read_instret_sel_lutinv ,\cu_ru/read_minstret_sel_lutinv }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/read_mscratch_sel_lutinv }),
    .c({\cu_ru/minstret [4],\cu_ru/minstret [4]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [4],\cu_ru/mscratch [4]}),
    .mi({open_n52250,\cu_ru/m_cycle_event/n4 [4]}),
    .sr(rst_pad),
    .f({_al_u7541_o,_al_u7550_o}),
    .q({open_n52254,\cu_ru/minstret [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7542|cu_ru/m_s_cause/reg0_b4  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/mcycle [4],\cu_ru/scause [4]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [4],data_csr[4]}),
    .sr(rst_pad),
    .f({_al_u7542_o,open_n52271}),
    .q({open_n52275,\cu_ru/scause [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7543|biu/bus_unit/mmu/reg2_b16  (
    .a({\cu_ru/read_cycle_sel_lutinv ,open_n52276}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n52277}),
    .c({satp[4],_al_u3162_o}),
    .clk(clk_pad),
    .d({\cu_ru/mcycle [4],_al_u3161_o}),
    .sr(rst_pad),
    .f({_al_u7543_o,open_n52295}),
    .q({open_n52299,\biu/paddress [80]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7544|cu_ru/m_s_tvec/reg1_b4  (
    .a({_al_u7430_o,_al_u7544_o}),
    .b({_al_u7541_o,_al_u7549_o}),
    .c({_al_u7542_o,_al_u7550_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7543_o,_al_u7551_o}),
    .sr(rst_pad),
    .f({_al_u7544_o,csr_data[4]}),
    .q({open_n52315,\cu_ru/mtvec [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7545|cu_ru/m_s_tval/reg0_b4  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n52316}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5248_o}),
    .c({\cu_ru/stval [4],\cu_ru/m_s_tval/n3 [4]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [4],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7545_o,open_n52333}),
    .q({open_n52337,\cu_ru/stval [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7547|cu_ru/m_s_epc/reg0_b4  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n52338}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({mtime_pad[4],_al_u5473_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [4],\cu_ru/m_s_epc/n2 [4]}),
    .sr(rst_pad),
    .f({_al_u7547_o,open_n52355}),
    .q({open_n52359,\cu_ru/sepc [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7548|cu_ru/m_s_tval/reg1_b4  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n52360}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [4],\cu_ru/m_s_tval/n3 [4]}),
    .clk(clk_pad),
    .d({\cu_ru/stvec [4],_al_u6479_o}),
    .sr(rst_pad),
    .f({_al_u7548_o,open_n52374}),
    .q({open_n52378,\cu_ru/mtval [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7549|_al_u7546  (
    .b({_al_u7547_o,\cu_ru/read_mepc_sel_lutinv }),
    .c({_al_u7548_o,\cu_ru/mepc [4]}),
    .d({_al_u7546_o,_al_u7545_o}),
    .f({_al_u7549_o,_al_u7546_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D*~A)))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~B*~(C*~(D*~A)))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001100000011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001001100000011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7553|cu_ru/m_s_tvec/reg0_b39  (
    .a({open_n52405,csr_data[39]}),
    .b({open_n52406,_al_u7553_o}),
    .c({_al_u7141_o,_al_u7554_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[39],id_system}),
    .mi({open_n52410,csr_data[39]}),
    .sr(rst_pad),
    .f({_al_u7553_o,_al_u7555_o}),
    .q({open_n52425,\cu_ru/stvec [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D*~A)))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~B*~(C*~(D*~A)))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001100000011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001001100000011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7557|cu_ru/m_s_tvec/reg0_b38  (
    .a({open_n52426,csr_data[38]}),
    .b({open_n52427,_al_u7557_o}),
    .c({_al_u7141_o,_al_u7558_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[38],id_system}),
    .mi({open_n52431,csr_data[38]}),
    .sr(rst_pad),
    .f({_al_u7557_o,_al_u7559_o}),
    .q({open_n52446,\cu_ru/stvec [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D*~A)))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001100000011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7561|cu_ru/m_s_tvec/reg0_b37  (
    .a({open_n52447,csr_data[37]}),
    .b({open_n52448,_al_u7561_o}),
    .c({_al_u7141_o,_al_u7562_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[37],id_system}),
    .mi({open_n52459,csr_data[37]}),
    .sr(rst_pad),
    .f({_al_u7561_o,_al_u7563_o}),
    .q({open_n52463,\cu_ru/stvec [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D*~A)))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001100000011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7565|cu_ru/m_s_tvec/reg0_b36  (
    .a({open_n52464,csr_data[36]}),
    .b({open_n52465,_al_u7565_o}),
    .c({_al_u7141_o,_al_u7566_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[36],id_system}),
    .mi({open_n52476,csr_data[36]}),
    .sr(rst_pad),
    .f({_al_u7565_o,_al_u7567_o}),
    .q({open_n52480,\cu_ru/stvec [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D*~A)))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~B*~(C*~(D*~A)))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001100000011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001001100000011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7569|cu_ru/m_s_tvec/reg0_b31  (
    .a({open_n52481,csr_data[31]}),
    .b({open_n52482,_al_u7569_o}),
    .c({_al_u7141_o,_al_u7570_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[31],id_system}),
    .mi({open_n52486,csr_data[31]}),
    .sr(rst_pad),
    .f({_al_u7569_o,_al_u7571_o}),
    .q({open_n52501,\cu_ru/stvec [31]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7573|cu_ru/m_s_cause/reg0_b3  (
    .a({\cu_ru/read_scause_sel_lutinv ,open_n52502}),
    .b({\cu_ru/n90 [32],_al_u5157_o}),
    .c({\cu_ru/scause [3],_al_u6729_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mie ,\cu_ru/trap_cause [3]}),
    .sr(rst_pad),
    .f({_al_u7573_o,open_n52519}),
    .q({open_n52523,\cu_ru/scause [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7574|cu_ru/m_s_scratch/reg1_b3  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n52524}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/sepc [3]}),
    .c({satp[3],data_csr[3]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [3],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n52528,data_csr[3]}),
    .sr(rst_pad),
    .f({_al_u7574_o,_al_u5517_o}),
    .q({open_n52543,\cu_ru/sscratch [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7575|_al_u9602  (
    .a({\cu_ru/read_sepc_sel_lutinv ,open_n52544}),
    .b({\cu_ru/read_mip_sel_lutinv ,_al_u2844_o}),
    .c({\cu_ru/sepc [3],\cu_ru/sepc [3]}),
    .d({\cu_ru/m_sip [3],\cu_ru/m_s_status/n2 }),
    .f({_al_u7575_o,_al_u9602_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7576|_al_u7608  (
    .b({_al_u7574_o,_al_u7606_o}),
    .c({_al_u7575_o,_al_u7607_o}),
    .d({_al_u7573_o,_al_u7605_o}),
    .f({_al_u7576_o,_al_u7608_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7577|cu_ru/m_s_scratch/reg0_b3  (
    .a({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcause [3],\cu_ru/mtval [3]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [3],data_csr[3]}),
    .mi({open_n52594,data_csr[3]}),
    .sr(rst_pad),
    .f({_al_u7577_o,_al_u6501_o}),
    .q({open_n52609,\cu_ru/mscratch [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*D)"),
    //.LUT1("(B*A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111111111111),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7578|cu_ru/m_s_tvec/reg1_b3  (
    .a({_al_u7576_o,open_n52610}),
    .b({_al_u7577_o,open_n52611}),
    .c({\cu_ru/read_medeleg_sel_lutinv ,_al_u7583_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/medeleg [3],_al_u7578_o}),
    .sr(rst_pad),
    .f({_al_u7578_o,csr_data[3]}),
    .q({open_n52627,\cu_ru/mtvec [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7580|cu_ru/m_s_tval/reg1_b3  (
    .a({_al_u6788_o,open_n52628}),
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [3],\cu_ru/m_s_tval/n3 [3]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [3],_al_u6501_o}),
    .sr(rst_pad),
    .f({_al_u7580_o,open_n52646}),
    .q({open_n52650,\cu_ru/mtval [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7581|cu_ru/m_s_epc/reg1_b3  (
    .a({\cu_ru/read_mepc_sel_lutinv ,open_n52651}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/m_s_epc/n2 [3]}),
    .c({\cu_ru/mepc [3],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({\cu_ru/stvec [3],_al_u6630_o}),
    .sr(rst_pad),
    .f({_al_u7581_o,open_n52669}),
    .q({open_n52673,\cu_ru/mepc [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7582|_al_u6731  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n52674}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u2844_o}),
    .c({\cu_ru/stval [3],\cu_ru/mtvec [3]}),
    .d({\cu_ru/mtvec [3],\cu_ru/trap_target_m }),
    .f({_al_u7582_o,_al_u6731_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*~A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*~A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010101000111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0010101000111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7583|cu_ru/m_cycle_event/reg0_b3  (
    .a({_al_u7579_o,_al_u6763_o}),
    .b({_al_u7580_o,\cu_ru/read_time_sel_lutinv }),
    .c({_al_u7581_o,mtime_pad[3]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7582_o,\cu_ru/minstret [3]}),
    .mi({open_n52702,\cu_ru/m_cycle_event/n4 [3]}),
    .sr(rst_pad),
    .f({_al_u7583_o,_al_u7579_o}),
    .q({open_n52717,\cu_ru/minstret [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7586|ins_dec/reg5_b29  (
    .a({open_n52718,_al_u7585_o}),
    .b({open_n52719,_al_u7586_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[29],id_ins[29]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7586_o,open_n52736}),
    .q({open_n52740,ds1[29]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7589|ins_dec/reg5_b27  (
    .a({open_n52741,_al_u7588_o}),
    .b({open_n52742,_al_u7589_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[27],id_ins[27]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7589_o,open_n52755}),
    .q({open_n52759,ds1[27]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7592|ins_dec/reg5_b26  (
    .a({open_n52760,_al_u7591_o}),
    .b({open_n52761,_al_u7592_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[26],id_ins[26]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7592_o,open_n52774}),
    .q({open_n52778,ds1[26]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7595|ins_dec/reg5_b24  (
    .a({open_n52779,_al_u7594_o}),
    .b({open_n52780,_al_u7595_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[24],id_ins[24]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7595_o,open_n52797}),
    .q({open_n52801,ds1[24]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7598|ins_dec/reg5_b23  (
    .a({open_n52802,_al_u7597_o}),
    .b({open_n52803,_al_u7598_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[23],id_ins[23]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7598_o,open_n52820}),
    .q({open_n52824,ds1[23]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u7600|cu_ru/m_s_cause/reg1_b22  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [22],\cu_ru/mtval [22]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [22],data_csr[22]}),
    .mi({open_n52828,data_csr[22]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u7600_o,_al_u6539_o}),
    .q({open_n52843,\cu_ru/mcause [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7601|cu_ru/m_s_cause/reg0_b22  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({satp[22],\cu_ru/scause [22]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [22],data_csr[22]}),
    .sr(rst_pad),
    .f({_al_u7601_o,open_n52860}),
    .q({open_n52864,\cu_ru/scause [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7603|cu_ru/m_s_tvec/reg1_b22  (
    .a({_al_u7430_o,_al_u7603_o}),
    .b({_al_u7600_o,_al_u7608_o}),
    .c({_al_u7601_o,_al_u7609_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7602_o,_al_u7610_o}),
    .sr(rst_pad),
    .f({_al_u7603_o,csr_data[22]}),
    .q({open_n52884,\cu_ru/mtvec [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7604|biu/bus_unit/mmu/reg2_b34  (
    .a({\cu_ru/read_mepc_sel_lutinv ,open_n52885}),
    .b({\cu_ru/read_stvec_sel_lutinv ,open_n52886}),
    .c({\cu_ru/mepc [22],_al_u3107_o}),
    .clk(clk_pad),
    .d({\cu_ru/stvec [22],_al_u3106_o}),
    .sr(rst_pad),
    .f({_al_u7604_o,open_n52900}),
    .q({open_n52904,\biu/paddress [98]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7605|_al_u7642  (
    .b({\cu_ru/read_time_sel_lutinv ,\cu_ru/read_time_sel_lutinv }),
    .c({mtime_pad[22],mtime_pad[17]}),
    .d({_al_u7604_o,_al_u7641_o}),
    .f({_al_u7605_o,_al_u7642_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7606|cu_ru/m_s_tval/reg0_b22  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n52931}),
    .b({\cu_ru/read_mtval_sel_lutinv ,_al_u5305_o}),
    .c({\cu_ru/stval [22],\cu_ru/m_s_tval/n3 [22]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [22],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7606_o,open_n52948}),
    .q({open_n52952,\cu_ru/stval [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7607|cu_ru/m_s_epc/reg0_b22  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n52953}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [22],_al_u5549_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [22],\cu_ru/m_s_epc/n2 [22]}),
    .sr(rst_pad),
    .f({_al_u7607_o,open_n52970}),
    .q({open_n52974,\cu_ru/sepc [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7610|cu_ru/m_s_scratch/reg1_b22  (
    .a({\cu_ru/read_cycle_sel_lutinv ,open_n52975}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/stval [22]}),
    .c({\cu_ru/mcycle [22],data_csr[22]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [22],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n52986,data_csr[22]}),
    .sr(rst_pad),
    .f({_al_u7610_o,_al_u5305_o}),
    .q({open_n52990,\cu_ru/sscratch [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7612|biu/bus_unit/mmu/reg2_b32  (
    .a({\cu_ru/read_mcause_sel_lutinv ,open_n52991}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n52992}),
    .c({satp[20],_al_u3113_o}),
    .clk(clk_pad),
    .d({\cu_ru/mcause [20],_al_u3112_o}),
    .sr(rst_pad),
    .f({_al_u7612_o,open_n53010}),
    .q({open_n53014,\biu/paddress [96]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7613|cu_ru/m_s_scratch/reg1_b20  (
    .a({\cu_ru/read_instret_sel_lutinv ,open_n53015}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/stval [20]}),
    .c({\cu_ru/minstret [20],data_csr[20]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [20],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n53019,data_csr[20]}),
    .sr(rst_pad),
    .f({_al_u7613_o,_al_u5311_o}),
    .q({open_n53034,\cu_ru/sscratch [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7614|cu_ru/m_s_cause/reg0_b20  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/mcycle [20],\cu_ru/scause [20]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [20],data_csr[20]}),
    .sr(rst_pad),
    .f({_al_u7614_o,open_n53051}),
    .q({open_n53055,\cu_ru/scause [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7615|cu_ru/m_s_tvec/reg1_b20  (
    .a({_al_u7430_o,_al_u7615_o}),
    .b({_al_u7612_o,_al_u7620_o}),
    .c({_al_u7613_o,_al_u7621_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7614_o,_al_u7622_o}),
    .sr(rst_pad),
    .f({_al_u7615_o,csr_data[20]}),
    .q({open_n53071,\cu_ru/mtvec [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7617|cu_ru/m_s_epc/reg0_b20  (
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [20],_al_u5557_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u7616_o,\cu_ru/m_s_epc/n2 [20]}),
    .sr(rst_pad),
    .f({_al_u7617_o,open_n53090}),
    .q({open_n53094,\cu_ru/sepc [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7619|cu_ru/m_s_tval/reg0_b20  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n53095}),
    .b({\cu_ru/read_mtval_sel_lutinv ,_al_u5311_o}),
    .c({\cu_ru/stval [20],\cu_ru/m_s_tval/n3 [20]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [20],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7619_o,open_n53108}),
    .q({open_n53112,\cu_ru/stval [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7620|_al_u7618  (
    .a({open_n53113,\cu_ru/read_mtvec_sel_lutinv }),
    .b({_al_u7618_o,\cu_ru/read_mepc_sel_lutinv }),
    .c({_al_u7619_o,\cu_ru/mepc [20]}),
    .d({_al_u7617_o,\cu_ru/mtvec [20]}),
    .f({_al_u7620_o,_al_u7618_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7622|cu_ru/m_s_scratch/reg0_b20  (
    .a({\cu_ru/read_cycle_sel_lutinv ,open_n53138}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [20]}),
    .c({\cu_ru/mcycle [20],data_csr[20]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [20],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n53142,data_csr[20]}),
    .sr(rst_pad),
    .f({_al_u7622_o,_al_u5557_o}),
    .q({open_n53157,\cu_ru/mscratch [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7624|_al_u7625  (
    .b({\cu_ru/n64 [32],\cu_ru/read_stvec_sel_lutinv }),
    .c({sum,\cu_ru/stvec [18]}),
    .d({\cu_ru/n82 [14],_al_u7624_o}),
    .f({_al_u7624_o,_al_u7625_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u7626|cu_ru/m_s_cause/reg1_b18  (
    .a({\cu_ru/read_cycle_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [18],\cu_ru/mtval [18]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [18],data_csr[18]}),
    .mi({open_n53187,data_csr[18]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u7626_o,_al_u6549_o}),
    .q({open_n53202,\cu_ru/mcause [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7627|cu_ru/m_s_scratch/reg0_b18  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,open_n53203}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [18]}),
    .c({\cu_ru/mcycle [18],data_csr[18]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [18],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n53214,data_csr[18]}),
    .sr(rst_pad),
    .f({_al_u7627_o,_al_u5569_o}),
    .q({open_n53218,\cu_ru/mscratch [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7628|cu_ru/m_s_tvec/reg1_b18  (
    .a({open_n53219,_al_u7628_o}),
    .b({_al_u7626_o,_al_u7633_o}),
    .c({_al_u7627_o,_al_u7634_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7625_o,_al_u7635_o}),
    .sr(rst_pad),
    .f({_al_u7628_o,csr_data[18]}),
    .q({open_n53239,\cu_ru/mtvec [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7629|cu_ru/m_s_tval/reg0_b18  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n53240}),
    .b({\cu_ru/read_time_sel_lutinv ,_al_u5320_o}),
    .c({mtime_pad[18],\cu_ru/m_s_tval/n3 [18]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [18],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7629_o,open_n53257}),
    .q({open_n53261,\cu_ru/stval [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7630|cu_ru/m_s_tval/reg1_b18  (
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [18],\cu_ru/m_s_tval/n3 [18]}),
    .clk(clk_pad),
    .d({_al_u7629_o,_al_u6549_o}),
    .sr(rst_pad),
    .f({_al_u7630_o,open_n53277}),
    .q({open_n53281,\cu_ru/mtval [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7632|biu/bus_unit/mmu/reg2_b30  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n53282}),
    .b({\cu_ru/read_mepc_sel_lutinv ,open_n53283}),
    .c({\cu_ru/mepc [18],_al_u3119_o}),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [18],_al_u3118_o}),
    .sr(rst_pad),
    .f({_al_u7632_o,open_n53297}),
    .q({open_n53301,\biu/paddress [94]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7635|cu_ru/m_s_cause/reg0_b18  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({satp[18],\cu_ru/scause [18]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [18],data_csr[18]}),
    .sr(rst_pad),
    .f({_al_u7635_o,open_n53318}),
    .q({open_n53322,\cu_ru/scause [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"))
    \_al_u7637|_al_u7497  (
    .a({\cu_ru/read_instret_sel_lutinv ,\cu_ru/read_cycle_sel_lutinv }),
    .b({\cu_ru/n90 [32],\cu_ru/n90 [32]}),
    .c({\cu_ru/minstret [17],\cu_ru/mcycle [7]}),
    .d({mprv,\cu_ru/mstatus [7]}),
    .f({_al_u7637_o,_al_u7497_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7638|cu_ru/m_s_scratch/reg0_b17  (
    .a({\cu_ru/read_mcause_sel_lutinv ,open_n53343}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [17]}),
    .c({\cu_ru/mcause [17],data_csr[17]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [17],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n53347,data_csr[17]}),
    .sr(rst_pad),
    .f({_al_u7638_o,_al_u5573_o}),
    .q({open_n53362,\cu_ru/mscratch [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7640|cu_ru/m_cycle_event/reg0_b17  (
    .a({_al_u7430_o,\cu_ru/read_mcycle_sel_lutinv }),
    .b({_al_u7637_o,\cu_ru/read_minstret_sel_lutinv }),
    .c({_al_u7638_o,\cu_ru/minstret [17]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7639_o,\cu_ru/mcycle [17]}),
    .mi({open_n53366,\cu_ru/m_cycle_event/n4 [17]}),
    .sr(rst_pad),
    .f({_al_u7640_o,_al_u7639_o}),
    .q({open_n53381,\cu_ru/minstret [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7641|cu_ru/m_s_tval/reg0_b17  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n53382}),
    .b({\cu_ru/read_mtval_sel_lutinv ,_al_u5323_o}),
    .c({\cu_ru/stval [17],\cu_ru/m_s_tval/n3 [17]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [17],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7641_o,open_n53395}),
    .q({open_n53399,\cu_ru/stval [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7643|biu/bus_unit/mmu/reg2_b29  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n53400}),
    .b({\cu_ru/read_mepc_sel_lutinv ,open_n53401}),
    .c({\cu_ru/mepc [17],_al_u3122_o}),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [17],_al_u3121_o}),
    .sr(rst_pad),
    .f({_al_u7643_o,open_n53415}),
    .q({open_n53419,\biu/paddress [93]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7644|cu_ru/m_s_epc/reg0_b17  (
    .a({\cu_ru/read_sepc_sel_lutinv ,open_n53420}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [17],_al_u5573_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [17],\cu_ru/m_s_epc/n2 [17]}),
    .sr(rst_pad),
    .f({_al_u7644_o,open_n53437}),
    .q({open_n53441,\cu_ru/sepc [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7645|cu_ru/m_s_tvec/reg1_b17  (
    .a({open_n53442,_al_u7640_o}),
    .b({_al_u7643_o,_al_u7645_o}),
    .c({_al_u7644_o,_al_u7646_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7642_o,_al_u7647_o}),
    .sr(rst_pad),
    .f({_al_u7645_o,csr_data[17]}),
    .q({open_n53458,\cu_ru/mtvec [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7646|cu_ru/m_s_scratch/reg1_b17  (
    .a({\cu_ru/read_cycle_sel_lutinv ,open_n53459}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/stval [17]}),
    .c({\cu_ru/mcycle [17],data_csr[17]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [17],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n53463,data_csr[17]}),
    .sr(rst_pad),
    .f({_al_u7646_o,_al_u5323_o}),
    .q({open_n53478,\cu_ru/sscratch [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7647|cu_ru/m_s_cause/reg0_b17  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({satp[17],\cu_ru/scause [17]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [17],data_csr[17]}),
    .sr(rst_pad),
    .f({_al_u7647_o,open_n53495}),
    .q({open_n53499,\cu_ru/scause [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7650|ins_dec/reg5_b16  (
    .a({open_n53500,_al_u7649_o}),
    .b({open_n53501,_al_u7650_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[16],id_ins[16]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7650_o,open_n53518}),
    .q({open_n53522,ds1[16]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7652|cu_ru/m_s_scratch/reg1_b12  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n53523}),
    .b({\cu_ru/n90 [32],\cu_ru/sepc [12]}),
    .c({\cu_ru/sscratch [12],data_csr[12]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mstatus [12],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n53534,data_csr[12]}),
    .sr(rst_pad),
    .f({_al_u7652_o,_al_u5593_o}),
    .q({open_n53538,\cu_ru/sscratch [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7654|biu/bus_unit/mmu/reg2_b24  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,open_n53539}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n53540}),
    .c({satp[12],_al_u3137_o}),
    .clk(clk_pad),
    .d({\cu_ru/mcycle [12],_al_u3136_o}),
    .sr(rst_pad),
    .f({_al_u7654_o,open_n53558}),
    .q({open_n53562,\biu/paddress [88]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7655|cu_ru/m_s_cause/reg0_b12  (
    .a({\cu_ru/read_cycle_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/mcycle [12],\cu_ru/scause [12]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [12],data_csr[12]}),
    .sr(rst_pad),
    .f({_al_u7655_o,open_n53579}),
    .q({open_n53583,\cu_ru/scause [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7656|cu_ru/m_s_tvec/reg1_b12  (
    .a({open_n53584,_al_u7656_o}),
    .b({_al_u7654_o,_al_u7661_o}),
    .c({_al_u7655_o,_al_u7662_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7653_o,_al_u7663_o}),
    .sr(rst_pad),
    .f({_al_u7656_o,csr_data[12]}),
    .q({open_n53604,\cu_ru/mtvec [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7657|cu_ru/m_s_scratch/reg0_b12  (
    .a({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [12],\cu_ru/mtval [12]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [12],data_csr[12]}),
    .mi({open_n53615,data_csr[12]}),
    .sr(rst_pad),
    .f({_al_u7657_o,_al_u6561_o}),
    .q({open_n53619,\cu_ru/mscratch [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7658|cu_ru/m_s_tval/reg0_b12  (
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5338_o}),
    .c({\cu_ru/stval [12],\cu_ru/m_s_tval/n3 [12]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u7657_o,_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7658_o,open_n53634}),
    .q({open_n53638,\cu_ru/stval [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0001010110111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u7659|_al_u9667  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,\cu_ru/m_s_status/n2 }),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u2844_o}),
    .c({\cu_ru/mepc [12],\cu_ru/sepc [12]}),
    .d({\cu_ru/mtvec [12],\cu_ru/mepc [12]}),
    .f({_al_u7659_o,_al_u9667_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7660|cu_ru/m_s_epc/reg0_b12  (
    .a({\cu_ru/read_time_sel_lutinv ,open_n53659}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({mtime_pad[12],_al_u5593_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [12],\cu_ru/m_s_epc/n2 [12]}),
    .sr(rst_pad),
    .f({_al_u7660_o,open_n53676}),
    .q({open_n53680,\cu_ru/sepc [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*B*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7661|_al_u3250  (
    .b({_al_u7659_o,open_n53683}),
    .c({_al_u7660_o,\cu_ru/mideleg_int_ctrl/sti_ack_s }),
    .d({_al_u7658_o,\cu_ru/mideleg_int_ctrl/n29_lutinv }),
    .f({_al_u7661_o,_al_u3250_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7662|cu_ru/m_cycle_event/reg0_b12  (
    .a({\cu_ru/read_instret_sel_lutinv ,\cu_ru/read_minstret_sel_lutinv }),
    .b({\cu_ru/read_medeleg_sel_lutinv ,\cu_ru/read_mscratch_sel_lutinv }),
    .c({\cu_ru/minstret [12],\cu_ru/minstret [12]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/medeleg [12],\cu_ru/mscratch [12]}),
    .mi({open_n53711,\cu_ru/m_cycle_event/n4 [12]}),
    .sr(rst_pad),
    .f({_al_u7662_o,_al_u7663_o}),
    .q({open_n53726,\cu_ru/minstret [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7665|cu_ru/m_s_scratch/reg1_b8  (
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/stval [8]}),
    .c({\cu_ru/sscratch [8],data_csr[8]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/n82 [14],\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({open_n53739,data_csr[8]}),
    .sr(rst_pad),
    .f({_al_u7665_o,_al_u5164_o}),
    .q({open_n53743,\cu_ru/sscratch [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7666|cu_ru/m_s_epc/reg0_b8  (
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [8],_al_u5361_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({_al_u7665_o,\cu_ru/m_s_epc/n2 [8]}),
    .sr(rst_pad),
    .f({_al_u7666_o,open_n53762}),
    .q({open_n53766,\cu_ru/sepc [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7667|cu_ru/m_s_cause/reg0_b8  (
    .a({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/scause [8],\cu_ru/scause [8]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [8],data_csr[8]}),
    .sr(rst_pad),
    .f({_al_u7667_o,open_n53783}),
    .q({open_n53787,\cu_ru/scause [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u7668|_al_u7438  (
    .b({\cu_ru/read_instret_sel_lutinv ,\cu_ru/read_satp_sel_lutinv }),
    .c({\cu_ru/minstret [8],satp[28]}),
    .d({_al_u7667_o,_al_u7437_o}),
    .f({_al_u7668_o,_al_u7438_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7671|cu_ru/m_cycle_event/reg0_b8  (
    .a({_al_u7666_o,\cu_ru/read_minstret_sel_lutinv }),
    .b({_al_u7668_o,\cu_ru/read_satp_sel_lutinv }),
    .c({_al_u7669_o,satp[8]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7670_o,\cu_ru/minstret [8]}),
    .mi({open_n53820,\cu_ru/m_cycle_event/n4 [8]}),
    .sr(rst_pad),
    .f({_al_u7671_o,_al_u7669_o}),
    .q({open_n53824,\cu_ru/minstret [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7672|cu_ru/m_s_tval/reg1_b8  (
    .a({_al_u7401_o,open_n53825}),
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mstatus [8],\cu_ru/m_s_tval/n3 [8]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [8],_al_u6443_o}),
    .sr(rst_pad),
    .f({_al_u7672_o,open_n53839}),
    .q({open_n53843,\cu_ru/mtval [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7673|cu_ru/m_s_tval/reg0_b8  (
    .a({_al_u6788_o,open_n53844}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5164_o}),
    .c({\cu_ru/mcycle [8],\cu_ru/m_s_tval/n3 [8]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [8],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7673_o,open_n53861}),
    .q({open_n53865,\cu_ru/stval [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7675|biu/bus_unit/mmu/reg2_b20  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,open_n53866}),
    .b({\cu_ru/read_mepc_sel_lutinv ,open_n53867}),
    .c({\cu_ru/mepc [8],_al_u3149_o}),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [8],_al_u3148_o}),
    .sr(rst_pad),
    .f({_al_u7675_o,open_n53885}),
    .q({open_n53889,\biu/paddress [84]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7676|cu_ru/m_s_tvec/reg1_b8  (
    .a({_al_u7672_o,open_n53890}),
    .b({_al_u7673_o,open_n53891}),
    .c({_al_u7674_o,_al_u7676_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7675_o,_al_u7671_o}),
    .sr(rst_pad),
    .f({_al_u7676_o,csr_data[8]}),
    .q({open_n53911,\cu_ru/mtvec [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~(~A*~(~C*B)))"),
    //.LUTG0("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~(~A*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010000000),
    .INIT_LUTF1(16'b0000000010101110),
    .INIT_LUTG0(16'b1000110010000000),
    .INIT_LUTG1(16'b0000000010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7679|cu_ru/m_s_tvec/reg0_b35  (
    .a({_al_u7678_o,csr_data[35]}),
    .b({rs1_data[35],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[35]}),
    .mi({open_n53915,csr_data[35]}),
    .sr(rst_pad),
    .f({_al_u7679_o,_al_u7678_o}),
    .q({open_n53930,\cu_ru/stvec [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D*~A)))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~B*~(C*~(D*~A)))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001001100000011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001001100000011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7681|cu_ru/m_s_tvec/reg0_b34  (
    .a({open_n53931,csr_data[34]}),
    .b({open_n53932,_al_u7681_o}),
    .c({_al_u7141_o,_al_u7682_o}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({rs1_data[34],id_system}),
    .mi({open_n53936,csr_data[34]}),
    .sr(rst_pad),
    .f({_al_u7681_o,_al_u7683_o}),
    .q({open_n53951,\cu_ru/stvec [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7686|ins_dec/reg5_b25  (
    .a({open_n53952,_al_u7685_o}),
    .b({open_n53953,_al_u7686_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[25],id_ins[25]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7686_o,open_n53970}),
    .q({open_n53974,ds1[25]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7688|ins_dec/reg5_b21  (
    .a({open_n53975,_al_u7688_o}),
    .b({open_n53976,_al_u7689_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[21],id_ins[21]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7688_o,open_n53993}),
    .q({open_n53997,ds1[21]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7691|cu_ru/m_s_scratch/reg1_b2  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,open_n53998}),
    .b({\cu_ru/read_sscratch_sel_lutinv ,\cu_ru/scause [2]}),
    .c({\cu_ru/mcycle [2],data_csr[2]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [2],\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .mi({open_n54009,data_csr[2]}),
    .sr(rst_pad),
    .f({_al_u7691_o,_al_u5662_o}),
    .q({open_n54013,\cu_ru/sscratch [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7692|biu/bus_unit/mmu/reg2_b14  (
    .b({\cu_ru/read_satp_sel_lutinv ,open_n54016}),
    .c({satp[2],_al_u3168_o}),
    .clk(clk_pad),
    .d({_al_u7691_o,_al_u3167_o}),
    .sr(rst_pad),
    .f({_al_u7692_o,open_n54030}),
    .q({open_n54034,\biu/paddress [78]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7693|cu_ru/m_s_scratch/reg0_b2  (
    .a({\cu_ru/read_cycle_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [2],\cu_ru/mtval [2]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [2],data_csr[2]}),
    .mi({open_n54045,data_csr[2]}),
    .sr(rst_pad),
    .f({_al_u7693_o,_al_u6523_o}),
    .q({open_n54049,\cu_ru/mscratch [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u7694|_al_u4180  (
    .b({_al_u7240_o,open_n54052}),
    .c({id_ins[22],id_ins[22]}),
    .d({_al_u7239_o,_al_u3214_o}),
    .f({_al_u7694_o,_al_u4180_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7696|cu_ru/m_s_cause/reg0_b2  (
    .a({\cu_ru/read_mcause_sel_lutinv ,open_n54073}),
    .b({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/scause [2],_al_u5662_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [2],\cu_ru/trap_cause [2]}),
    .sr(rst_pad),
    .f({_al_u7696_o,open_n54090}),
    .q({open_n54094,\cu_ru/scause [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*A*~(D*C))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000001000100010),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u7697|_al_u7695  (
    .a({_al_u7430_o,_al_u7693_o}),
    .b({_al_u7692_o,_al_u7694_o}),
    .c({_al_u7695_o,\cu_ru/read_medeleg_sel_lutinv }),
    .d({_al_u7696_o,\cu_ru/medeleg [2]}),
    .f({_al_u7697_o,_al_u7695_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7699|cu_ru/m_s_tval/reg1_b2  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n54115}),
    .b({\cu_ru/read_sepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/sepc [2],\cu_ru/m_s_tval/n3 [2]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [2],_al_u6523_o}),
    .sr(rst_pad),
    .f({_al_u7699_o,open_n54133}),
    .q({open_n54137,\cu_ru/mtval [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100000001001100),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7700|cu_ru/m_s_tvec/reg0_b2  (
    .a({\cu_ru/read_mtvec_sel_lutinv ,csr_data[2]}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u7141_o}),
    .c({\cu_ru/stvec [2],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [2],id_ins_pc[2]}),
    .mi({open_n54148,csr_data[2]}),
    .sr(rst_pad),
    .f({_al_u7700_o,_al_u7887_o}),
    .q({open_n54152,\cu_ru/stvec [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7701|cu_ru/m_s_epc/reg1_b2  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n54153}),
    .b({\cu_ru/read_mepc_sel_lutinv ,\cu_ru/m_s_epc/n2 [2]}),
    .c({\cu_ru/mepc [2],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({\cu_ru/stval [2],_al_u6652_o}),
    .sr(rst_pad),
    .f({_al_u7701_o,open_n54171}),
    .q({open_n54175,\cu_ru/mepc [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("~(C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000111111111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7702|cu_ru/m_s_tvec/reg1_b2  (
    .a({_al_u7698_o,open_n54176}),
    .b({_al_u7699_o,open_n54177}),
    .c({_al_u7700_o,_al_u7702_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7701_o,_al_u7697_o}),
    .sr(rst_pad),
    .f({_al_u7702_o,csr_data[2]}),
    .q({open_n54197,\cu_ru/mtvec [2]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7704|ins_dec/reg5_b15  (
    .a({open_n54198,_al_u7704_o}),
    .b({open_n54199,_al_u7705_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[15],id_ins[15]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7704_o,open_n54212}),
    .q({open_n54216,ds1[15]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7708|ins_dec/reg5_b13  (
    .a({open_n54217,_al_u7707_o}),
    .b({open_n54218,_al_u7708_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[13],_al_u3217_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7708_o,open_n54235}),
    .q({open_n54239,ds1[13]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7712|cu_ru/m_cycle_event/reg0_b0  (
    .a({\cu_ru/read_instret_sel_lutinv ,open_n54240}),
    .b({\cu_ru/read_medeleg_sel_lutinv ,\cu_ru/m_cycle_event/mcountinhibit[2] }),
    .c({\cu_ru/minstret [0],wb_valid}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/medeleg [0],_al_u3253_o}),
    .mi({open_n54251,\cu_ru/m_cycle_event/n4 [0]}),
    .sr(rst_pad),
    .f({_al_u7712_o,\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o }),
    .q({open_n54255,\cu_ru/minstret [0]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u7713|_al_u3202  (
    .b({\cu_ru/read_mtvec_sel_lutinv ,open_n54258}),
    .c({\cu_ru/mtvec [0],_al_u3201_o}),
    .d({_al_u7712_o,_al_u3195_o}),
    .f({_al_u7713_o,\cu_ru/m_s_tvec/n0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u7714|_al_u7715  (
    .b({_al_u7478_o,\cu_ru/n66_lutinv }),
    .c({\cu_ru/mstatus [1],\cu_ru/sscratch [0]}),
    .d({_al_u6777_o,\cu_ru/read_sscratch_sel_lutinv }),
    .f({\cu_ru/n66_lutinv ,_al_u7715_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*~B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"))
    \_al_u7717|_al_u7716  (
    .b({id_ins[20],_al_u3392_o}),
    .c({_al_u3394_o,\cu_ru/mcountinhibit }),
    .d({_al_u7716_o,id_ins[25]}),
    .f({_al_u7717_o,_al_u7716_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(~C*A*~(D*B))"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(~C*A*~(D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b0000001000001010),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b0000001000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7719|cu_ru/m_s_cause/reg1_b0  (
    .a({_al_u7715_o,open_n54323}),
    .b({\cu_ru/read_mcause_sel_lutinv ,_al_u6702_o}),
    .c({_al_u7718_o,\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({\cu_ru/mcause [0],\cu_ru/trap_cause [0]}),
    .sr(rst_pad),
    .f({_al_u7719_o,open_n54341}),
    .q({open_n54345,\cu_ru/mcause [0]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7720|cu_ru/m_s_cause/reg0_b0  (
    .a({\cu_ru/read_minstret_sel_lutinv ,open_n54346}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/n41 }),
    .c({\cu_ru/minstret [0],_al_u5674_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [0],_al_u4232_o}),
    .sr(rst_pad),
    .f({_al_u7720_o,open_n54363}),
    .q({open_n54367,\cu_ru/scause [0]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7721|biu/bus_unit/mmu/reg2_b12  (
    .a({\cu_ru/read_mscratch_sel_lutinv ,open_n54368}),
    .b({\cu_ru/read_satp_sel_lutinv ,open_n54369}),
    .c({satp[0],_al_u3174_o}),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [0],_al_u3173_o}),
    .sr(rst_pad),
    .f({_al_u7721_o,open_n54387}),
    .q({open_n54391,\biu/paddress [76]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7722|cu_ru/m_s_tvec/reg1_b0  (
    .a({_al_u7713_o,_al_u7722_o}),
    .b({_al_u7719_o,_al_u7724_o}),
    .c({_al_u7720_o,_al_u7725_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7721_o,_al_u7726_o}),
    .sr(rst_pad),
    .f({_al_u7722_o,csr_data[0]}),
    .q({open_n54411,\cu_ru/mtvec [0]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7724|_al_u7723  (
    .a({open_n54412,_al_u6788_o}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/read_mepc_sel_lutinv }),
    .c({\cu_ru/stvec [0],\cu_ru/mcycle [0]}),
    .d({_al_u7723_o,\cu_ru/mepc [0]}),
    .f({_al_u7724_o,_al_u7723_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111010101011100),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111010101011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7728|_al_u6760  (
    .a({_al_u3399_o,open_n54437}),
    .b({_al_u6760_o,open_n54438}),
    .c({id_ins[28],id_ins[30]}),
    .d({id_ins[27],id_ins[31]}),
    .f({_al_u7728_o,_al_u6760_o}));
  // ../../RTL/CPU/ID/ins_dec.v(674)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~C*~A*~(~D*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000010100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7729|ins_dec/and_clr_reg  (
    .a({\ins_dec/n71 ,open_n54463}),
    .b({_al_u3938_o,_al_u3217_o}),
    .c({\ins_dec/n141_lutinv ,_al_u3384_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u7728_o,id_system}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7729_o,\ins_dec/n71 }),
    .q({open_n54479,and_clr}));  // ../../RTL/CPU/ID/ins_dec.v(674)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*D))"),
    //.LUT1("(~D*~C*~B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110011001100),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7730|ins_dec/mem_csr_data_or_reg  (
    .a({_al_u7729_o,open_n54480}),
    .b({\ins_dec/n149_lutinv ,\ins_dec/n149_lutinv }),
    .c({_al_u6059_o,\ins_dec/funct5_8_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,_al_u3938_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7730_o,open_n54493}),
    .q({open_n54497,mem_csr_data_or}));  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(B*~(~D*~C)))"),
    //.LUT1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111011101010),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7731|ins_dec/shift_l_reg  (
    .a({open_n54498,\ins_dec/ins_slli }),
    .b({open_n54499,_al_u4094_o}),
    .c({_al_u7730_o,\ins_dec/op_32_imm_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/n235 ,_al_u3925_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7731_o,\ins_dec/n235 }),
    .q({open_n54515,shift_l}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(C*~B*~D)"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"))
    \_al_u7734|_al_u7733  (
    .b({\exu/store_addr_mis ,_al_u2838_o}),
    .c({_al_u7733_o,_al_u2847_o}),
    .d({\exu/load_addr_mis ,load_acc_fault}),
    .f({_al_u7734_o,_al_u7733_o}));
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7735|exu/reg5_b35  (
    .a({_al_u6724_o,open_n54538}),
    .b({_al_u7734_o,open_n54539}),
    .c({_al_u6725_o,addr_ex[35]}),
    .clk(clk_pad),
    .d({_al_u7195_o,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({ex_more_exception_neg_lutinv,open_n54557}),
    .q({open_n54561,wb_exc_code[35]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7800|cu_ru/m_s_epc/reg0_b9  (
    .a({_al_u6788_o,open_n54562}),
    .b({\cu_ru/read_sepc_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/mcycle [9],_al_u5357_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [9],\cu_ru/m_s_epc/n2 [9]}),
    .sr(rst_pad),
    .f({_al_u7800_o,open_n54579}),
    .q({open_n54583,\cu_ru/sepc [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7801|cu_ru/m_s_tval/reg0_b9  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n54584}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5160_o}),
    .c({\cu_ru/mepc [9],\cu_ru/m_s_tval/n3 [9]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [9],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7801_o,open_n54601}),
    .q({open_n54605,\cu_ru/stval [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u7802|_al_u6789  (
    .c({_al_u6791_o,_al_u6769_o}),
    .d({_al_u6764_o,_al_u6764_o}),
    .f({\cu_ru/read_mideleg_sel_lutinv ,\cu_ru/read_stval_sel_lutinv }));
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7803|cu_ru/m_cycle_event/reg0_b5  (
    .a({\cu_ru/read_time_sel_lutinv ,_al_u6763_o}),
    .b({\cu_ru/read_mideleg_sel_lutinv ,\cu_ru/read_mideleg_sel_lutinv }),
    .c({mtime_pad[9],\cu_ru/minstret [5]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mideleg [9],\cu_ru/mideleg [5]}),
    .mi({open_n54633,\cu_ru/m_cycle_event/n4 [5]}),
    .sr(rst_pad),
    .f({_al_u7803_o,_al_u7875_o}),
    .q({open_n54648,\cu_ru/minstret [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7804|cu_ru/m_s_tval/reg1_b9  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n54649}),
    .b({\cu_ru/read_stvec_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [9],\cu_ru/m_s_tval/n3 [9]}),
    .clk(clk_pad),
    .d({\cu_ru/stvec [9],_al_u6441_o}),
    .sr(rst_pad),
    .f({_al_u7804_o,open_n54667}),
    .q({open_n54671,\cu_ru/mtval [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7805|cu_ru/m_s_tvec/reg1_b9  (
    .a({_al_u7800_o,_al_u7805_o}),
    .b({_al_u7801_o,_al_u7809_o}),
    .c({_al_u7803_o,_al_u7811_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7804_o,_al_u7812_o}),
    .sr(rst_pad),
    .f({_al_u7805_o,csr_data[9]}),
    .q({open_n54691,\cu_ru/mtvec [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7806|cu_ru/m_s_scratch/reg0_b9  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n54692}),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/sepc [9]}),
    .c({\cu_ru/mscratch [9],data_csr[9]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [9],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n54703,data_csr[9]}),
    .sr(rst_pad),
    .f({_al_u7806_o,_al_u5357_o}),
    .q({open_n54707,\cu_ru/mscratch [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(~D*~C))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1000100010000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u7807|_al_u7808  (
    .a({open_n54708,_al_u7478_o}),
    .b({open_n54709,_al_u7807_o}),
    .c({_al_u3388_o,s_ext_int_pad}),
    .d({_al_u6765_o,\cu_ru/m_s_ip/seip }),
    .f({_al_u7807_o,_al_u7808_o}));
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~B*A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7809|biu/bus_unit/mmu/reg2_b21  (
    .a({_al_u7806_o,open_n54730}),
    .b({_al_u7808_o,open_n54731}),
    .c({\cu_ru/read_satp_sel_lutinv ,_al_u3146_o}),
    .clk(clk_pad),
    .d({satp[9],_al_u3145_o}),
    .sr(rst_pad),
    .f({_al_u7809_o,open_n54745}),
    .q({open_n54749,\biu/paddress [85]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~C*A*~(D*B))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~C*A*~(D*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0000001000001010),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0000001000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7811|cu_ru/m_s_cause/reg0_b9  (
    .a({_al_u7810_o,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/n84 [10],\cu_ru/scause [9]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [9],data_csr[9]}),
    .sr(rst_pad),
    .f({_al_u7811_o,open_n54766}),
    .q({open_n54770,\cu_ru/scause [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7817|ins_dec/reg5_b33  (
    .a({open_n54771,_al_u7816_o}),
    .b({open_n54772,_al_u7817_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[33],id_ins[31]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7817_o,open_n54785}),
    .q({open_n54789,ds1[33]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7820|ins_dec/reg5_b32  (
    .a({open_n54790,_al_u7819_o}),
    .b({open_n54791,_al_u7820_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[32],id_ins[31]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7820_o,open_n54804}),
    .q({open_n54808,ds1[32]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7823|ins_dec/reg5_b30  (
    .a({open_n54809,_al_u7822_o}),
    .b({open_n54810,_al_u7823_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[30],id_ins[30]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7823_o,open_n54827}),
    .q({open_n54831,ds1[30]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7826|ins_dec/reg5_b28  (
    .a({open_n54832,_al_u7825_o}),
    .b({open_n54833,_al_u7826_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[28],id_ins[28]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7826_o,open_n54846}),
    .q({open_n54850,ds1[28]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7829|ins_dec/reg5_b19  (
    .a({open_n54851,_al_u7828_o}),
    .b({open_n54852,_al_u7829_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[19],id_ins[19]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7829_o,open_n54865}),
    .q({open_n54869,ds1[19]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7832|ins_dec/reg5_b14  (
    .a({open_n54870,_al_u7831_o}),
    .b({open_n54871,_al_u7832_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[14],_al_u3216_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7832_o,open_n54884}),
    .q({open_n54888,ds1[14]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7843|ins_dec/reg5_b22  (
    .a({open_n54889,_al_u7842_o}),
    .b({open_n54890,_al_u7843_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[22],id_ins[22]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7843_o,open_n54903}),
    .q({open_n54907,ds1[22]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7846|ins_dec/reg5_b20  (
    .a({open_n54908,_al_u7845_o}),
    .b({open_n54909,_al_u7846_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[20],id_ins[20]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7846_o,open_n54926}),
    .q({open_n54930,ds1[20]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7849|ins_dec/reg5_b18  (
    .a({open_n54931,_al_u7848_o}),
    .b({open_n54932,_al_u7849_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[18],id_ins[18]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7849_o,open_n54945}),
    .q({open_n54949,ds1[18]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111000001110),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111000001110),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7852|ins_dec/reg5_b17  (
    .a({open_n54950,_al_u7851_o}),
    .b({open_n54951,_al_u7852_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[17],id_ins[17]}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7852_o,open_n54968}),
    .q({open_n54972,ds1[17]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111000001110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7855|ins_dec/reg5_b12  (
    .a({open_n54973,_al_u7854_o}),
    .b({open_n54974,_al_u7855_o}),
    .c({_al_u7141_o,\ins_dec/op_lui_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[12],_al_u3384_o}),
    .sr(\ins_dec/n107 ),
    .f({_al_u7855_o,open_n54987}),
    .q({open_n54991,ds1[12]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7857|cu_ru/m_s_scratch/reg1_b1  (
    .a({\cu_ru/read_sscratch_sel_lutinv ,open_n54992}),
    .b({\cu_ru/read_satp_sel_lutinv ,\cu_ru/sepc [1]}),
    .c({satp[1],data_csr[1]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sscratch [1],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n55003,data_csr[1]}),
    .sr(rst_pad),
    .f({_al_u7857_o,_al_u5604_o}),
    .q({open_n55007,\cu_ru/sscratch [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7858|cu_ru/m_s_tval/reg1_b1  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n55008}),
    .b({\cu_ru/read_sepc_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/sepc [1],\cu_ru/m_s_tval/n3 [1]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [1],_al_u6545_o}),
    .sr(rst_pad),
    .f({_al_u7858_o,open_n55022}),
    .q({open_n55026,\cu_ru/mtval [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7860|cu_ru/m_s_cause/reg0_b1  (
    .a({\cu_ru/read_cycle_sel_lutinv ,open_n55027}),
    .b({\cu_ru/read_scause_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/mcycle [1],_al_u7337_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [1],\cu_ru/trap_cause [1]}),
    .sr(rst_pad),
    .f({_al_u7860_o,open_n55044}),
    .q({open_n55048,\cu_ru/scause [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTG1("(D*~(C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1100000011001111),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7861|cu_ru/m_s_cause/reg1_b1  (
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/trap_cause [1]}),
    .c({\cu_ru/mcause [1],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u7860_o,_al_u7335_o}),
    .sr(rst_pad),
    .f({_al_u7861_o,open_n55068}),
    .q({open_n55072,\cu_ru/mcause [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7862|cu_ru/m_s_scratch/reg0_b1  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mscratch_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [1],\cu_ru/mtval [1]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mscratch [1],data_csr[1]}),
    .mi({open_n55076,data_csr[1]}),
    .sr(rst_pad),
    .f({_al_u7862_o,_al_u6545_o}),
    .q({open_n55091,\cu_ru/mscratch [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7863|cu_ru/m_s_ip/ssip_reg  (
    .c({\cu_ru/m_sip [1],\cu_ru/m_s_ip/u12_sel_is_2_o }),
    .ce(\cu_ru/m_s_ip/u11_sel_is_0_o ),
    .clk(clk_pad),
    .d({_al_u7807_o,\cu_ru/m_s_ip/n0 }),
    .mi({open_n55099,data_csr[1]}),
    .sr(rst_pad),
    .f({_al_u7863_o,\cu_ru/m_s_ip/u11_sel_is_0_o }),
    .q({open_n55114,\cu_ru/m_sip [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*C))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u7865|_al_u7859  (
    .a({_al_u7859_o,_al_u7857_o}),
    .b({_al_u7861_o,_al_u7858_o}),
    .c({_al_u7862_o,\cu_ru/read_mepc_sel_lutinv }),
    .d({_al_u7864_o,\cu_ru/mepc [1]}),
    .f({_al_u7865_o,_al_u7859_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000001001100),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0100000001001100),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7866|cu_ru/m_s_tvec/reg0_b1  (
    .a({\cu_ru/read_time_sel_lutinv ,csr_data[1]}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u7141_o}),
    .c({mtime_pad[1],id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [1],id_ins_pc[1]}),
    .mi({open_n55138,csr_data[1]}),
    .sr(rst_pad),
    .f({_al_u7866_o,_al_u7893_o}),
    .q({open_n55153,\cu_ru/stvec [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7867|cu_ru/m_s_tvec/reg1_b1  (
    .a({open_n55154,_al_u7865_o}),
    .b({\cu_ru/read_mtvec_sel_lutinv ,_al_u7867_o}),
    .c({\cu_ru/mtvec [1],_al_u7868_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7866_o,_al_u7869_o}),
    .sr(rst_pad),
    .f({_al_u7867_o,csr_data[1]}),
    .q({open_n55170,\cu_ru/mtvec [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7868|cu_ru/m_s_tval/reg0_b1  (
    .a({_al_u7401_o,open_n55171}),
    .b({\cu_ru/read_stval_sel_lutinv ,_al_u5347_o}),
    .c({\cu_ru/mstatus [1],\cu_ru/m_s_tval/n3 [1]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [1],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7868_o,open_n55184}),
    .q({open_n55188,\cu_ru/stval [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*C*B*A)"),
    //.LUT1("(A*~(D*~(~C*~B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111111111111),
    .INIT_LUT1(16'b0000001010101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7874|cu_ru/m_s_tvec/reg1_b5  (
    .a({_al_u7873_o,_al_u7874_o}),
    .b({\cu_ru/n64 [32],_al_u7875_o}),
    .c({\cu_ru/n90 [32],_al_u7880_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mstatus [5],_al_u7885_o}),
    .sr(rst_pad),
    .f({_al_u7874_o,csr_data[5]}),
    .q({open_n55204,\cu_ru/mtvec [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u7876|cu_ru/m_s_cause/reg1_b5  (
    .a({\cu_ru/read_mcycle_sel_lutinv ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/read_mcause_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcycle [5],\cu_ru/mtval [5]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mcause [5],data_csr[5]}),
    .mi({open_n55208,data_csr[5]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u7876_o,_al_u6457_o}),
    .q({open_n55223,\cu_ru/mcause [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7877|cu_ru/m_s_cause/reg0_b5  (
    .a({\cu_ru/read_cycle_sel_lutinv ,_al_u5157_o}),
    .b({\cu_ru/read_scause_sel_lutinv ,\cu_ru/m_s_cause/mux2_b0_sel_is_2_o }),
    .c({\cu_ru/mcycle [5],\cu_ru/scause [5]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/scause [5],data_csr[5]}),
    .sr(rst_pad),
    .f({_al_u7877_o,open_n55240}),
    .q({open_n55244,\cu_ru/scause [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7880|cu_ru/m_s_scratch/reg1_b5  (
    .a({_al_u7876_o,\cu_ru/read_sscratch_sel_lutinv }),
    .b({_al_u7877_o,\cu_ru/read_mscratch_sel_lutinv }),
    .c({_al_u7878_o,\cu_ru/mscratch [5]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u7879_o,\cu_ru/sscratch [5]}),
    .mi({open_n55248,data_csr[5]}),
    .sr(rst_pad),
    .f({_al_u7880_o,_al_u7878_o}),
    .q({open_n55263,\cu_ru/sscratch [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*B))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7881|cu_ru/m_s_tval/reg1_b5  (
    .a({\cu_ru/read_mtval_sel_lutinv ,open_n55264}),
    .b({\cu_ru/read_mip_sel_lutinv ,\cu_ru/trap_target_m }),
    .c({\cu_ru/m_sip [5],\cu_ru/m_s_tval/n3 [5]}),
    .clk(clk_pad),
    .d({\cu_ru/mtval [5],_al_u6457_o}),
    .sr(rst_pad),
    .f({_al_u7881_o,open_n55278}),
    .q({open_n55282,\cu_ru/mtval [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7882|cu_ru/m_s_tval/reg0_b5  (
    .a({\cu_ru/read_stval_sel_lutinv ,open_n55283}),
    .b({\cu_ru/read_mepc_sel_lutinv ,_al_u5215_o}),
    .c({\cu_ru/mepc [5],\cu_ru/m_s_tval/n3 [5]}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stval [5],_al_u5157_o}),
    .sr(rst_pad),
    .f({_al_u7882_o,open_n55296}),
    .q({open_n55300,\cu_ru/stval [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~(D*B)*~(C*A))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~(D*B)*~(C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0001001101011111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0001001101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7884|cu_ru/m_s_epc/reg0_b5  (
    .a({\cu_ru/read_sepc_sel_lutinv ,open_n55301}),
    .b({\cu_ru/read_stvec_sel_lutinv ,_al_u5157_o}),
    .c({\cu_ru/sepc [5],_al_u5429_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/stvec [5],\cu_ru/m_s_epc/n2 [5]}),
    .sr(rst_pad),
    .f({_al_u7884_o,open_n55318}),
    .q({open_n55322,\cu_ru/sepc [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u7885|_al_u7883  (
    .a({_al_u7881_o,\cu_ru/read_mtvec_sel_lutinv }),
    .b({_al_u7882_o,\cu_ru/read_time_sel_lutinv }),
    .c({_al_u7883_o,mtime_pad[5]}),
    .d({_al_u7884_o,\cu_ru/mtvec [5]}),
    .f({_al_u7885_o,_al_u7883_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b1100101000000000),
    .INIT_LUT1(16'b1100101000000000),
    .MODE("LOGIC"))
    \_al_u7897|_al_u7969  (
    .a({\biu/l1d_out [15],\biu/l1d_out [15]}),
    .b({uncache_data[15],uncache_data[15]}),
    .c({_al_u3224_o,_al_u3224_o}),
    .d({\exu/lsu/n2_lutinv ,\exu/lsu/n0_lutinv }),
    .f({_al_u7897_o,_al_u7969_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b1011000010000000),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u7898|_al_u9011  (
    .a({open_n55363,uncache_data[3]}),
    .b({_al_u3224_o,_al_u3224_o}),
    .c({\exu/lsu/n0_lutinv ,\exu/lsu/n0_lutinv }),
    .d({uncache_data[7],\biu/l1d_out [3]}),
    .f({_al_u7898_o,_al_u9011_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b0011000000111111),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u7899|_al_u8739  (
    .b({\biu/l1d_out [7],uncache_data[23]}),
    .c({_al_u3224_o,_al_u3224_o}),
    .d({_al_u7898_o,\biu/l1d_out [23]}),
    .f({_al_u7899_o,_al_u8739_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b1100101000000000),
    .INIT_LUT1(16'b1100101000000000),
    .MODE("LOGIC"))
    \_al_u7901|_al_u7967  (
    .a({\biu/l1d_out [23],\biu/l1d_out [31]}),
    .b({uncache_data[23],uncache_data[31]}),
    .c({_al_u3224_o,_al_u3224_o}),
    .d({\exu/lsu/n5_lutinv ,\exu/lsu/n5_lutinv }),
    .f({_al_u7901_o,_al_u7967_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b1100101000000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100101000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7902|_al_u7900  (
    .a({_al_u7897_o,\biu/l1d_out [31]}),
    .b({_al_u7899_o,uncache_data[31]}),
    .c({_al_u7900_o,_al_u3224_o}),
    .d({_al_u7901_o,\exu/lsu/n8_lutinv }),
    .f({_al_u7902_o,_al_u7900_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u7904|_al_u3430  (
    .b({open_n55452,\exu/alu_au/n5 }),
    .c({unsign,unsign}),
    .d({ex_size[0],\exu/alu_au/n15 }),
    .f({\exu/lsu/n51 ,_al_u3430_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7906|_al_u8552  (
    .b({_al_u3224_o,\exu/lsu/mux27_b56_sel_is_3_o }),
    .c({uncache_data[33],\exu/n60_lutinv }),
    .d({\biu/l1d_out [33],_al_u7906_o}),
    .f({_al_u7906_o,_al_u8552_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7907|_al_u8605  (
    .b({_al_u3224_o,_al_u3224_o}),
    .c({uncache_data[25],\biu/l1d_out [30]}),
    .d({\biu/l1d_out [25],uncache_data[30]}),
    .f({_al_u7907_o,_al_u8605_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT_LUT0(16'b1111001110101111),
    .INIT_LUT1(16'b0101001100000000),
    .MODE("LOGIC"))
    \_al_u7908|_al_u8702  (
    .a({_al_u7906_o,_al_u7906_o}),
    .b({_al_u7907_o,_al_u8383_o}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u7908_o,_al_u8702_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b1111001111000000),
    .MODE("LOGIC"))
    \_al_u7909|_al_u8444  (
    .b({_al_u3224_o,_al_u3224_o}),
    .c({uncache_data[9],\biu/l1d_out [38]}),
    .d({\biu/l1d_out [9],uncache_data[38]}),
    .f({_al_u7909_o,_al_u8444_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u7910|_al_u8859  (
    .a({open_n55567,uncache_data[41]}),
    .b({_al_u3224_o,uncache_data[17]}),
    .c({\biu/l1d_out [17],addr_ex[0]}),
    .d({uncache_data[17],addr_ex[1]}),
    .f({_al_u7910_o,_al_u8859_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUT1("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b0011111111110101),
    .INIT_LUT1(16'b0000000011001010),
    .MODE("LOGIC"))
    \_al_u7911|_al_u8855  (
    .a({_al_u7909_o,_al_u7910_o}),
    .b({_al_u7910_o,_al_u8383_o}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u7911_o,_al_u8855_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7914|_al_u4049  (
    .c({\exu/lsu/n0_lutinv ,\exu/lsu/n0_lutinv }),
    .d({uncache_data[7],\exu/alu_data_mem_csr [2]}),
    .f({\exu/lsu/n22 [7],\exu/lsu/n1 [2]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7916|_al_u7915  (
    .a({\exu/lsu/n22 [7],uncache_data[31]}),
    .b({_al_u7915_o,uncache_data[15]}),
    .c({uncache_data[23],addr_ex[0]}),
    .d({\exu/lsu/n5_lutinv ,addr_ex[1]}),
    .f({_al_u7916_o,_al_u7915_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7917|_al_u7957  (
    .b({open_n55662,_al_u7956_o}),
    .c({\exu/lsu/n51 ,\exu/c_stb_lutinv }),
    .d({_al_u7916_o,_al_u7916_o}),
    .f({\exu/lsu/n52 [10],_al_u7957_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~(~D*C)*~(~B*~A))"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b1110111000001110),
    .MODE("LOGIC"))
    \_al_u7920|_al_u7918  (
    .a({_al_u7918_o,uncache_data[33]}),
    .b({_al_u7919_o,uncache_data[17]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u7920_o,_al_u7918_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(~D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7922|_al_u9073  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[9],data_rd[10]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u7922_o,_al_u9073_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*~A)))"),
    //.LUTF1("(C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*~A)))"),
    //.LUTG1("(C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000000100001111),
    .INIT_LUTF1(16'b0010000011110000),
    .INIT_LUTG0(16'b0000000100001111),
    .INIT_LUTG1(16'b0010000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7923|_al_u7921  (
    .a({_al_u7905_o,\exu/lsu/n52 [10]}),
    .b({_al_u7913_o,_al_u7920_o}),
    .c({_al_u7921_o,\exu/c_stb_lutinv }),
    .d({_al_u7922_o,\exu/n59_lutinv }),
    .f({_al_u7923_o,_al_u7921_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7926|_al_u7924  (
    .a({_al_u7924_o,\exu/c_stb_lutinv }),
    .b({_al_u7925_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [9],ds1[9]}),
    .d({rd_data_add,ds2[9]}),
    .f({_al_u7926_o,_al_u7924_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(C@D))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(C@D))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b0000110011000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b0000110011000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7927|_al_u3437  (
    .a({_al_u7926_o,open_n55781}),
    .b({rd_data_xor,ds1[9]}),
    .c({ds1[9],ds2[9]}),
    .d({ds2[9],and_clr}),
    .f({_al_u7927_o,\exu/alu_au/alu_and [9]}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(B*~D))"),
    //.LUTF1("(~B*~(A*~(D*C)))"),
    //.LUTG0("~(~C*~(B*~D))"),
    //.LUTG1("(~B*~(A*~(D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111100),
    .INIT_LUTF1(16'b0011000100010001),
    .INIT_LUTG0(16'b1111000011111100),
    .INIT_LUTG1(16'b0011000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7928|exu/reg1_b9  (
    .a({_al_u7927_o,open_n55806}),
    .b({_al_u2855_o,_al_u7928_o}),
    .c({\exu/alu_au/alu_and [9],_al_u7930_o}),
    .clk(clk_pad),
    .d({rd_data_and,_al_u7923_o}),
    .sr(rst_pad),
    .f({_al_u7928_o,open_n55824}),
    .q({open_n55828,data_rd[9]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u7929|_al_u7930  (
    .a({open_n55829,_al_u2855_o}),
    .b({data_rd[9],\exu/n57 [9]}),
    .c({shift_r,data_rd[8]}),
    .d({data_rd[10],shift_l}),
    .f({\exu/n57 [9],_al_u7930_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b1111001111000000),
    .INIT_LUT1(16'b1111001111000000),
    .MODE("LOGIC"))
    \_al_u7932|_al_u8383  (
    .b({_al_u3224_o,_al_u3224_o}),
    .c({uncache_data[24],uncache_data[41]}),
    .d({\biu/l1d_out [24],\biu/l1d_out [41]}),
    .f({_al_u7932_o,_al_u8383_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~C*~(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0000001100001010),
    .INIT_LUTF1(16'b1111010100111111),
    .INIT_LUTG0(16'b0000001100001010),
    .INIT_LUTG1(16'b1111010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7934|_al_u8720  (
    .a({_al_u7932_o,_al_u7932_o}),
    .b({_al_u7933_o,_al_u8402_o}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u7934_o,_al_u8720_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b0000001111001111),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b0000001111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7935|_al_u7933  (
    .b({_al_u3224_o,_al_u3224_o}),
    .c({\biu/l1d_out [8],uncache_data[16]}),
    .d({uncache_data[8],\biu/l1d_out [16]}),
    .f({_al_u7935_o,_al_u7933_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUT1("(~(~D*C)*~(B*A))"),
    .INIT_LUT0(16'b0011111111111010),
    .INIT_LUT1(16'b0111011100000111),
    .MODE("LOGIC"))
    \_al_u7938|_al_u7937  (
    .a({_al_u7934_o,_al_u7935_o}),
    .b({_al_u7937_o,_al_u7936_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u7938_o,_al_u7937_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b1010000011000000),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b1010000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7939|_al_u8877  (
    .a({uncache_data[32],uncache_data[32]}),
    .b({uncache_data[16],uncache_data[16]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u7939_o,_al_u8877_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~(~D*C)*~(~B*~A))"),
    //.LUTG0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~(~D*C)*~(~B*~A))"),
    .INIT_LUTF0(16'b0000110000001010),
    .INIT_LUTF1(16'b1110111000001110),
    .INIT_LUTG0(16'b0000110000001010),
    .INIT_LUTG1(16'b1110111000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7941|_al_u7940  (
    .a({_al_u7939_o,uncache_data[8]}),
    .b({_al_u7940_o,uncache_data[24]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u7941_o,_al_u7940_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(~D*~(~C*~B))"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"))
    \_al_u7943|_al_u9036  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[8],data_rd[11]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u7943_o,_al_u9036_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*~A)))"),
    //.LUTF1("(C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*~A)))"),
    //.LUTG1("(C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000000100001111),
    .INIT_LUTF1(16'b0010000011110000),
    .INIT_LUTG0(16'b0000000100001111),
    .INIT_LUTG1(16'b0010000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7944|_al_u7942  (
    .a({_al_u7905_o,\exu/lsu/n52 [10]}),
    .b({_al_u7938_o,_al_u7941_o}),
    .c({_al_u7942_o,\exu/c_stb_lutinv }),
    .d({_al_u7943_o,\exu/n59_lutinv }),
    .f({_al_u7944_o,_al_u7942_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7947|_al_u7945  (
    .a({_al_u7945_o,\exu/c_stb_lutinv }),
    .b({_al_u7946_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [8],ds1[8]}),
    .d({rd_data_add,ds2[8]}),
    .f({_al_u7947_o,_al_u7945_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*(D@C)))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1010001000101010),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u7948|_al_u9114  (
    .a({_al_u7947_o,_al_u9113_o}),
    .b({rd_data_xor,rd_data_xor}),
    .c({ds1[8],ds1[0]}),
    .d({ds2[8],ds2[0]}),
    .f({_al_u7948_o,_al_u9114_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(B*~D))"),
    //.LUTF1("(~B*~(A*~(D*C)))"),
    //.LUTG0("~(~C*~(B*~D))"),
    //.LUTG1("(~B*~(A*~(D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111100),
    .INIT_LUTF1(16'b0011000100010001),
    .INIT_LUTG0(16'b1111000011111100),
    .INIT_LUTG1(16'b0011000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7949|exu/reg1_b8  (
    .a({_al_u7948_o,open_n56080}),
    .b({_al_u2855_o,_al_u7949_o}),
    .c({\exu/alu_au/alu_and [8],_al_u7951_o}),
    .clk(clk_pad),
    .d({rd_data_and,_al_u7944_o}),
    .sr(rst_pad),
    .f({_al_u7949_o,open_n56098}),
    .q({open_n56102,data_rd[8]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7950|_al_u7951  (
    .a({open_n56103,_al_u2855_o}),
    .b({data_rd[9],\exu/n57 [8]}),
    .c({shift_r,data_rd[7]}),
    .d({data_rd[8],shift_l}),
    .f({\exu/n57 [8],_al_u7951_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(B*~(C*D))"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b0000110011001100),
    .MODE("LOGIC"))
    \_al_u7953|_al_u7956  (
    .b({\exu/n60_lutinv ,\exu/n59_lutinv }),
    .c({_al_u7912_o,_al_u7912_o}),
    .d({_al_u3415_o,_al_u3415_o}),
    .f({_al_u7953_o,_al_u7956_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7954|_al_u9088  (
    .c({data_rd[7],data_rd[1]}),
    .d({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .f({_al_u7954_o,_al_u9088_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(~D*~(~C*~(B*~A)))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(~D*~(~C*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b0000000011110100),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b0000000011110100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7955|exu/reg1_b7  (
    .a({_al_u7902_o,_al_u7955_o}),
    .b({_al_u7953_o,_al_u7957_o}),
    .c({_al_u7954_o,_al_u7963_o}),
    .clk(clk_pad),
    .d({\exu/n59_lutinv ,_al_u7965_o}),
    .sr(rst_pad),
    .f({_al_u7955_o,open_n56195}),
    .q({open_n56199,data_rd[7]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7960|_al_u7958  (
    .a({_al_u7958_o,\exu/c_stb_lutinv }),
    .b({_al_u7959_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [7],ds1[7]}),
    .d({rd_data_add,ds2[7]}),
    .f({_al_u7960_o,_al_u7958_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u7961|_al_u3452  (
    .a({_al_u7960_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[7],ds1[7]}),
    .d({ds2[7],ds2[7]}),
    .f({_al_u7961_o,\exu/alu_au/n55 [7]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7963|_al_u7962  (
    .a({open_n56244,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [7],ds1[7]}),
    .d({_al_u7961_o,ds2[7]}),
    .f({_al_u7963_o,\exu/alu_au/n33 [7]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u7964|_al_u7965  (
    .a({open_n56269,_al_u2855_o}),
    .b({data_rd[8],\exu/n57 [7]}),
    .c({shift_r,data_rd[6]}),
    .d({data_rd[7],shift_l}),
    .f({\exu/n57 [7],_al_u7965_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUTF0(16'b1100101000000000),
    .INIT_LUTF1(16'b1100101000000000),
    .INIT_LUTG0(16'b1100101000000000),
    .INIT_LUTG1(16'b1100101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7970|_al_u8423  (
    .a({\biu/l1d_out [39],\biu/l1d_out [39]}),
    .b({uncache_data[39],uncache_data[39]}),
    .c({_al_u3224_o,_al_u3224_o}),
    .d({\exu/lsu/n8_lutinv ,\exu/lsu/n0_lutinv }),
    .f({_al_u7970_o,_al_u8423_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b1100101000000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100101000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7971|_al_u7968  (
    .a({_al_u7967_o,\biu/l1d_out [23]}),
    .b({_al_u7968_o,uncache_data[23]}),
    .c({_al_u7969_o,_al_u3224_o}),
    .d({_al_u7970_o,\exu/lsu/n2_lutinv }),
    .f({_al_u7971_o,_al_u7968_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7973|_al_u7972  (
    .c({\exu/lsu/n53 ,unsign}),
    .d({_al_u7971_o,ex_size[1]}),
    .f({_al_u7973_o,\exu/lsu/n53 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7974|_al_u8747  (
    .a({open_n56366,uncache_data[47]}),
    .b({open_n56367,uncache_data[31]}),
    .c({_al_u3224_o,addr_ex[0]}),
    .d({uncache_data[47],addr_ex[1]}),
    .f({_al_u7974_o,_al_u8747_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~(~B*A)))"),
    //.LUTF1("(D*~(~C*~(~B*A)))"),
    //.LUTG0("(D*~(~C*~(~B*A)))"),
    //.LUTG1("(D*~(~C*~(~B*A)))"),
    .INIT_LUTF0(16'b1111001000000000),
    .INIT_LUTF1(16'b1111001000000000),
    .INIT_LUTG0(16'b1111001000000000),
    .INIT_LUTG1(16'b1111001000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7975|_al_u8420  (
    .a({\biu/l1d_out [47],\biu/l1d_out [47]}),
    .b({_al_u3224_o,_al_u3224_o}),
    .c({_al_u7974_o,_al_u7974_o}),
    .d({\exu/lsu/n5_lutinv ,\exu/lsu/n2_lutinv }),
    .f({_al_u7975_o,_al_u8420_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b1100101000000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100101000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7979|_al_u7976  (
    .a({_al_u7975_o,\biu/l1d_out [31]}),
    .b({_al_u7976_o,uncache_data[31]}),
    .c({_al_u7977_o,_al_u3224_o}),
    .d({_al_u7978_o,\exu/lsu/n0_lutinv }),
    .f({_al_u7979_o,_al_u7976_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~(~B*~A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000111000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u7980|_al_u8421  (
    .a({open_n56440,\biu/l1d_out [63]}),
    .b({open_n56441,_al_u3224_o}),
    .c({_al_u3224_o,_al_u7981_o}),
    .d({\biu/l1d_out [63],\exu/lsu/n8_lutinv }),
    .f({_al_u7980_o,_al_u8421_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u7982|_al_u7981  (
    .c({_al_u7981_o,_al_u3224_o}),
    .d({_al_u7980_o,uncache_data[63]}),
    .f({_al_u7982_o,_al_u7981_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7984|_al_u7912  (
    .c({unsign,unsign}),
    .d({ex_size[2],ex_size[2]}),
    .f({\exu/lsu/n56 ,_al_u7912_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~(C*B)*~(D*~A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~(C*B)*~(D*~A))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0010101000111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0010101000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7985|_al_u9046  (
    .a({_al_u7979_o,open_n56514}),
    .b({_al_u7982_o,open_n56515}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\biu/l1d_out [2]}),
    .d({\exu/lsu/n56 ,_al_u3224_o}),
    .f({_al_u7985_o,_al_u9046_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(~D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7986|_al_u9001  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[63],data_rd[12]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u7986_o,_al_u9001_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D*~(B*~A)))"),
    //.LUT1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111101111110000),
    .INIT_LUT1(16'b1101111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u7987|exu/reg1_b63  (
    .a({_al_u7905_o,_al_u7987_o}),
    .b({_al_u7973_o,_al_u7997_o}),
    .c({_al_u7985_o,_al_u8002_o}),
    .clk(clk_pad),
    .d({_al_u7986_o,_al_u8009_o}),
    .sr(rst_pad),
    .f({_al_u7987_o,open_n56579}),
    .q({open_n56583,data_rd[63]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~B*A*~(D*C))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~B*A*~(D*C))"),
    .INIT_LUTF0(16'b1111010100111111),
    .INIT_LUTF1(16'b0000001000100010),
    .INIT_LUTG0(16'b1111010100111111),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7990|_al_u7988  (
    .a({_al_u7988_o,uncache_data[31]}),
    .b({\exu/lsu/n22 [15],uncache_data[23]}),
    .c({uncache_data[39],addr_ex[0]}),
    .d({\exu/lsu/n8_lutinv ,addr_ex[1]}),
    .f({_al_u7990_o,_al_u7988_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~D*~(C*~B))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~D*~(C*~B))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7991|_al_u8890  (
    .b({_al_u7990_o,open_n56610}),
    .c({\exu/lsu/n53 ,_al_u7912_o}),
    .d({\exu/lsu/n52 [10],_al_u7971_o}),
    .f({_al_u7991_o,_al_u8890_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u7992|_al_u8265  (
    .b({open_n56637,_al_u7981_o}),
    .c({\exu/lsu/n5_lutinv ,\exu/lsu/n5_lutinv }),
    .d({uncache_data[47],_al_u7980_o}),
    .f({\exu/lsu/n25 [31],_al_u8265_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~B*~A*~(D*C))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b0000000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7994|_al_u7993  (
    .a({\exu/lsu/n25 [31],uncache_data[55]}),
    .b({_al_u7993_o,uncache_data[39]}),
    .c({uncache_data[31],addr_ex[0]}),
    .d({\exu/lsu/n0_lutinv ,addr_ex[1]}),
    .f({_al_u7994_o,_al_u7993_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*A)))"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b0000001000001111),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u7995|_al_u8749  (
    .a({open_n56682,_al_u7991_o}),
    .b({_al_u7994_o,_al_u8748_o}),
    .c({\exu/lsu/n56 ,\exu/c_stb_lutinv }),
    .d({_al_u7991_o,\exu/n59_lutinv }),
    .f({_al_u7995_o,_al_u8749_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7996|_al_u8049  (
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/lsu/mux27_b56_sel_is_3_o }),
    .d({uncache_data[63],uncache_data[60]}),
    .f({\exu/lsu/n59 [63],\exu/lsu/n59 [60]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*A)))"),
    //.LUT1("(~C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000001000001111),
    .INIT_LUT1(16'b0000001000001111),
    .MODE("LOGIC"))
    \_al_u7997|_al_u8409  (
    .a({_al_u7995_o,_al_u7995_o}),
    .b({\exu/lsu/n59 [63],\exu/lsu/n59 [40]}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u7997_o,_al_u8409_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(C*D))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(C*D))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u7999|_al_u7998  (
    .b({data_rd[63],open_n56753}),
    .c({unsign,shift_r}),
    .d({\exu/mux27_b32_sel_is_1_o ,ex_size[2]}),
    .f({\exu/n57 [63],\exu/mux27_b32_sel_is_1_o }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u8001|_al_u8013  (
    .b({open_n56780,\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[62]}),
    .d({data_rd[62],\exu/n59_lutinv }),
    .f({_al_u8001_o,_al_u8013_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b0000110010001000),
    .MODE("LOGIC"))
    \_al_u8002|_al_u8000  (
    .a({\exu/n57 [63],open_n56801}),
    .b({_al_u8000_o,data_rd[63]}),
    .c({_al_u8001_o,ex_size[2]}),
    .d({shift_l,_al_u2855_o}),
    .f({_al_u8002_o,_al_u8000_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*(C@B))"),
    .INIT_LUT0(16'b1100100001000000),
    .INIT_LUT1(16'b0011110000000000),
    .MODE("LOGIC"))
    \_al_u8003|_al_u3455  (
    .a({open_n56822,_al_u3430_o}),
    .b({ds1[63],mem_csr_data_max}),
    .c({ds2[63],ds1[63]}),
    .d({rd_data_xor,ds2[63]}),
    .f({\exu/alu_au/n37 [63],\exu/alu_au/n53 [63]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*~B*~(D*~A))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000001000000011),
    .MODE("LOGIC"))
    \_al_u8005|_al_u8004  (
    .a({_al_u3459_o,\exu/alu_au/add_64 [63]}),
    .b({\exu/alu_au/n37 [63],\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [63],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8005_o,\exu/alu_au/n31 [63]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*A*~(D*C))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~B*A*~(D*C))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000001000100010),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8006|_al_u8007  (
    .a({open_n56863,\exu/c_stb_lutinv }),
    .b({ds1[63],\exu/alu_au/n35 [63]}),
    .c({ds2[63],rd_data_ds1}),
    .d({rd_data_or,ds1[63]}),
    .f({\exu/alu_au/n35 [63],_al_u8007_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100000111),
    .MODE("LOGIC"))
    \_al_u8009|_al_u8008  (
    .a({_al_u8005_o,and_clr}),
    .b({_al_u8007_o,rd_data_and}),
    .c({_al_u2855_o,ds1[63]}),
    .d({\exu/alu_au/n33 [63],ds2[63]}),
    .f({_al_u8009_o,\exu/alu_au/n33 [63]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8011|_al_u8449  (
    .a({open_n56908,uncache_data[62]}),
    .b({_al_u3224_o,uncache_data[38]}),
    .c({\biu/l1d_out [62],addr_ex[0]}),
    .d({uncache_data[62],addr_ex[1]}),
    .f({_al_u8011_o,_al_u8449_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1101111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8014|exu/reg1_b62  (
    .a({_al_u7905_o,_al_u8014_o}),
    .b({_al_u7973_o,_al_u8016_o}),
    .c({_al_u8012_o,_al_u8022_o}),
    .clk(clk_pad),
    .d({_al_u8013_o,_al_u8025_o}),
    .sr(rst_pad),
    .f({_al_u8014_o,open_n56946}),
    .q({open_n56950,data_rd[62]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u8015|_al_u8113  (
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/lsu/mux27_b56_sel_is_3_o }),
    .d({uncache_data[62],uncache_data[56]}),
    .f({\exu/lsu/n59 [62],\exu/lsu/n59 [56]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*A)))"),
    //.LUT1("(~C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000001000001111),
    .INIT_LUT1(16'b0000001000001111),
    .MODE("LOGIC"))
    \_al_u8016|_al_u8390  (
    .a({_al_u7995_o,_al_u7995_o}),
    .b({\exu/lsu/n59 [62],\exu/lsu/n59 [41]}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8016_o,_al_u8390_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8018|_al_u8017  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [62]}),
    .b({_al_u3467_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [62],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8018_o,\exu/alu_au/n31 [62]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u8019|_al_u8545  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[62],ds1[34]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8019_o,_al_u8545_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*(D@C)))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(A*~(B*(D@C)))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1010001000101010),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1010001000101010),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8020|_al_u8772  (
    .a({_al_u8019_o,_al_u8771_o}),
    .b({rd_data_xor,rd_data_xor}),
    .c({ds1[62],ds1[22]}),
    .d({ds2[62],ds2[22]}),
    .f({_al_u8020_o,_al_u8772_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8022|_al_u8021  (
    .a({_al_u8018_o,and_clr}),
    .b({_al_u8020_o,rd_data_and}),
    .c({_al_u2855_o,ds1[62]}),
    .d({\exu/alu_au/n33 [62],ds2[62]}),
    .f({_al_u8022_o,\exu/alu_au/n33 [62]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1100000010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1100000010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8023|_al_u8025  (
    .a({open_n57089,\exu/n57 [62]}),
    .b({data_rd[62],_al_u2855_o}),
    .c({data_rd[63],\exu/n54 [30]}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [62],_al_u8025_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8024|_al_u8031  (
    .b({data_rd[62],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[61]}),
    .d({data_rd[61],\exu/n59_lutinv }),
    .f({\exu/n54 [30],_al_u8031_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~(~B*~A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000111000000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u8027|_al_u8463  (
    .a({open_n57140,\biu/l1d_out [61]}),
    .b({open_n57141,_al_u3224_o}),
    .c({_al_u3224_o,_al_u8028_o}),
    .d({\biu/l1d_out [61],\exu/lsu/n8_lutinv }),
    .f({_al_u8027_o,_al_u8463_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u8029|_al_u8028  (
    .c({_al_u8028_o,_al_u3224_o}),
    .d({_al_u8027_o,uncache_data[61]}),
    .f({_al_u8029_o,_al_u8028_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*~A))"),
    //.LUT1("(~(C*B)*~(D*~A))"),
    .INIT_LUT0(16'b0010101000111111),
    .INIT_LUT1(16'b0010101000111111),
    .MODE("LOGIC"))
    \_al_u8030|_al_u8012  (
    .a({_al_u7979_o,_al_u7979_o}),
    .b({_al_u8029_o,_al_u8011_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/lsu/mux27_b56_sel_is_3_o }),
    .d({\exu/lsu/n56 ,\exu/lsu/n56 }),
    .f({_al_u8030_o,_al_u8012_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1101111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8032|exu/reg1_b61  (
    .a({_al_u7905_o,_al_u8032_o}),
    .b({_al_u7973_o,_al_u8034_o}),
    .c({_al_u8030_o,_al_u8040_o}),
    .clk(clk_pad),
    .d({_al_u8031_o,_al_u8043_o}),
    .sr(rst_pad),
    .f({_al_u8032_o,open_n57219}),
    .q({open_n57223,data_rd[61]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8033|_al_u8097  (
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/lsu/mux27_b56_sel_is_3_o }),
    .d({uncache_data[61],uncache_data[57]}),
    .f({\exu/lsu/n59 [61],\exu/lsu/n59 [57]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*A)))"),
    //.LUTF1("(~C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*A)))"),
    //.LUTG1("(~C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000001000001111),
    .INIT_LUTF1(16'b0000001000001111),
    .INIT_LUTG0(16'b0000001000001111),
    .INIT_LUTG1(16'b0000001000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8034|_al_u8371  (
    .a({_al_u7995_o,_al_u7995_o}),
    .b({\exu/lsu/n59 [61],\exu/lsu/n59 [42]}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8034_o,_al_u8371_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8036|_al_u8035  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [61]}),
    .b({_al_u3475_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [61],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8036_o,\exu/alu_au/n31 [61]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u8037|_al_u8524  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[61],ds1[35]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8037_o,_al_u8524_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*(D@C)))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(A*~(B*(D@C)))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1010001000101010),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1010001000101010),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8038|_al_u8598  (
    .a({_al_u8037_o,_al_u8597_o}),
    .b({rd_data_xor,rd_data_xor}),
    .c({ds1[61],ds1[31]}),
    .d({ds2[61],ds2[31]}),
    .f({_al_u8038_o,_al_u8598_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8040|_al_u8039  (
    .a({_al_u8036_o,and_clr}),
    .b({_al_u8038_o,rd_data_and}),
    .c({_al_u2855_o,ds1[61]}),
    .d({\exu/alu_au/n33 [61],ds2[61]}),
    .f({_al_u8040_o,\exu/alu_au/n33 [61]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110001000100),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000110001000100),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8041|_al_u8043  (
    .a({open_n57370,_al_u8041_o}),
    .b({data_rd[61],_al_u2855_o}),
    .c({data_rd[62],_al_u8042_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({_al_u8041_o,_al_u8043_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8042|_al_u8047  (
    .b({data_rd[61],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[60]}),
    .d({data_rd[60],\exu/n59_lutinv }),
    .f({_al_u8042_o,_al_u8047_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b1100101000000000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b1100101000000000),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8046|_al_u8045  (
    .a({open_n57421,\biu/l1d_out [60]}),
    .b({_al_u8045_o,uncache_data[60]}),
    .c({\exu/lsu/n56 ,_al_u3224_o}),
    .d({_al_u7979_o,\exu/lsu/mux27_b56_sel_is_3_o }),
    .f({_al_u8046_o,_al_u8045_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1101111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1101111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8048|exu/reg1_b60  (
    .a({_al_u7905_o,_al_u8048_o}),
    .b({_al_u7973_o,_al_u8050_o}),
    .c({_al_u8046_o,_al_u8056_o}),
    .clk(clk_pad),
    .d({_al_u8047_o,_al_u8059_o}),
    .sr(rst_pad),
    .f({_al_u8048_o,open_n57463}),
    .q({open_n57467,data_rd[60]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*A)))"),
    //.LUTF1("(~C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*A)))"),
    //.LUTG1("(~C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000001000001111),
    .INIT_LUTF1(16'b0000001000001111),
    .INIT_LUTG0(16'b0000001000001111),
    .INIT_LUTG1(16'b0000001000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8050|_al_u8352  (
    .a({_al_u7995_o,_al_u7995_o}),
    .b({\exu/lsu/n59 [60],\exu/lsu/n59 [43]}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8050_o,_al_u8352_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8052|_al_u8051  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [60]}),
    .b({_al_u3483_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [60],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8052_o,\exu/alu_au/n31 [60]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8053|_al_u8500  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[60],ds1[36]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8053_o,_al_u8500_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*(D@C)))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1010001000101010),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8054|_al_u9078  (
    .a({_al_u8053_o,_al_u9077_o}),
    .b({rd_data_xor,rd_data_xor}),
    .c({ds1[60],ds1[10]}),
    .d({ds2[60],ds2[10]}),
    .f({_al_u8054_o,_al_u9078_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8056|_al_u8055  (
    .a({_al_u8052_o,and_clr}),
    .b({_al_u8054_o,rd_data_and}),
    .c({_al_u2855_o,ds1[60]}),
    .d({\exu/alu_au/n33 [60],ds2[60]}),
    .f({_al_u8056_o,\exu/alu_au/n33 [60]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"))
    \_al_u8057|_al_u8059  (
    .a({open_n57578,_al_u8057_o}),
    .b({data_rd[60],_al_u2855_o}),
    .c({data_rd[61],_al_u8058_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({_al_u8057_o,_al_u8059_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8058|_al_u8063  (
    .b({data_rd[60],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[59]}),
    .d({data_rd[59],\exu/n59_lutinv }),
    .f({_al_u8058_o,_al_u8063_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~(C*~B)*~(D*~A))"),
    .INIT_LUT0(16'b0000001111001111),
    .INIT_LUT1(16'b1000101011001111),
    .MODE("LOGIC"))
    \_al_u8062|_al_u8061  (
    .a({_al_u7979_o,open_n57621}),
    .b({_al_u8061_o,_al_u3224_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\biu/l1d_out [59]}),
    .d({\exu/lsu/n56 ,uncache_data[59]}),
    .f({_al_u8062_o,_al_u8061_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1101111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1101111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8064|exu/reg1_b59  (
    .a({_al_u7905_o,_al_u8064_o}),
    .b({_al_u7973_o,_al_u8066_o}),
    .c({_al_u8062_o,_al_u8072_o}),
    .clk(clk_pad),
    .d({_al_u8063_o,_al_u8075_o}),
    .sr(rst_pad),
    .f({_al_u8064_o,open_n57659}),
    .q({open_n57663,data_rd[59]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8065|_al_u8081  (
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/lsu/mux27_b56_sel_is_3_o }),
    .d(uncache_data[59:58]),
    .f(\exu/lsu/n59 [59:58]));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*A)))"),
    //.LUT1("(~C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000001000001111),
    .INIT_LUT1(16'b0000001000001111),
    .MODE("LOGIC"))
    \_al_u8066|_al_u8333  (
    .a({_al_u7995_o,_al_u7995_o}),
    .b({\exu/lsu/n59 [59],\exu/lsu/n59 [44]}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8066_o,_al_u8333_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8068|_al_u8067  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [59]}),
    .b({_al_u3498_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [59],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8068_o,\exu/alu_au/n31 [59]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8069|_al_u8477  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[59],ds1[37]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8069_o,_al_u8477_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*(D@C)))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1010001000101010),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8070|_al_u9041  (
    .a({_al_u8069_o,_al_u9040_o}),
    .b({rd_data_xor,rd_data_xor}),
    .c({ds1[59],ds1[11]}),
    .d({ds2[59],ds2[11]}),
    .f({_al_u8070_o,_al_u9041_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8072|_al_u8071  (
    .a({_al_u8068_o,and_clr}),
    .b({_al_u8070_o,rd_data_and}),
    .c({_al_u2855_o,ds1[59]}),
    .d({\exu/alu_au/n33 [59],ds2[59]}),
    .f({_al_u8072_o,\exu/alu_au/n33 [59]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110010001000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u8073|_al_u8075  (
    .a({open_n57798,\exu/n57 [59]}),
    .b({data_rd[59],_al_u2855_o}),
    .c({data_rd[60],_al_u8074_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [59],_al_u8075_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8074|_al_u8079  (
    .b({data_rd[59],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[58]}),
    .d({data_rd[58],\exu/n59_lutinv }),
    .f({_al_u8074_o,_al_u8079_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~(C*~B)*~(D*~A))"),
    .INIT_LUT0(16'b0000001111001111),
    .INIT_LUT1(16'b1000101011001111),
    .MODE("LOGIC"))
    \_al_u8078|_al_u8077  (
    .a({_al_u7979_o,open_n57841}),
    .b({_al_u8077_o,_al_u3224_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\biu/l1d_out [58]}),
    .d({\exu/lsu/n56 ,uncache_data[58]}),
    .f({_al_u8078_o,_al_u8077_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1101111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8080|exu/reg1_b58  (
    .a({_al_u7905_o,_al_u8080_o}),
    .b({_al_u7973_o,_al_u8082_o}),
    .c({_al_u8078_o,_al_u8088_o}),
    .clk(clk_pad),
    .d({_al_u8079_o,_al_u8091_o}),
    .sr(rst_pad),
    .f({_al_u8080_o,open_n57875}),
    .q({open_n57879,data_rd[58]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*A)))"),
    //.LUT1("(~C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000001000001111),
    .INIT_LUT1(16'b0000001000001111),
    .MODE("LOGIC"))
    \_al_u8082|_al_u8313  (
    .a({_al_u7995_o,_al_u7995_o}),
    .b({\exu/lsu/n59 [58],\exu/lsu/n59 [45]}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8082_o,_al_u8313_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8084|_al_u8083  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [58]}),
    .b({_al_u3506_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [58],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8084_o,\exu/alu_au/n31 [58]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u8085|_al_u8455  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[58],ds1[38]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8085_o,_al_u8455_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*(D@C)))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(A*~(B*(D@C)))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1010001000101010),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1010001000101010),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8086|_al_u9006  (
    .a({_al_u8085_o,_al_u9005_o}),
    .b({rd_data_xor,rd_data_xor}),
    .c({ds1[58],ds1[12]}),
    .d({ds2[58],ds2[12]}),
    .f({_al_u8086_o,_al_u9006_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8088|_al_u8087  (
    .a({_al_u8084_o,and_clr}),
    .b({_al_u8086_o,rd_data_and}),
    .c({_al_u2855_o,ds1[58]}),
    .d({\exu/alu_au/n33 [58],ds2[58]}),
    .f({_al_u8088_o,\exu/alu_au/n33 [58]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000110010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8089|_al_u8091  (
    .a({open_n57994,\exu/n57 [58]}),
    .b({data_rd[58],_al_u2855_o}),
    .c({data_rd[59],_al_u8090_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [58],_al_u8091_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8090|_al_u8095  (
    .b({data_rd[58],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[57]}),
    .d({data_rd[57],\exu/n59_lutinv }),
    .f({_al_u8090_o,_al_u8095_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(~(C*B)*~(D*~A))"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(~(C*B)*~(D*~A))"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b0010101000111111),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b0010101000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8094|_al_u8093  (
    .a({_al_u7979_o,open_n58045}),
    .b({_al_u8093_o,_al_u3224_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,uncache_data[57]}),
    .d({\exu/lsu/n56 ,\biu/l1d_out [57]}),
    .f({_al_u8094_o,_al_u8093_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1101111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8096|exu/reg1_b57  (
    .a({_al_u7905_o,_al_u8096_o}),
    .b({_al_u7973_o,_al_u8098_o}),
    .c({_al_u8094_o,_al_u8104_o}),
    .clk(clk_pad),
    .d({_al_u8095_o,_al_u8107_o}),
    .sr(rst_pad),
    .f({_al_u8096_o,open_n58083}),
    .q({open_n58087,data_rd[57]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*A)))"),
    //.LUTF1("(~C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*A)))"),
    //.LUTG1("(~C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000001000001111),
    .INIT_LUTF1(16'b0000001000001111),
    .INIT_LUTG0(16'b0000001000001111),
    .INIT_LUTG1(16'b0000001000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8098|_al_u8293  (
    .a({_al_u7995_o,_al_u7995_o}),
    .b({\exu/lsu/n59 [57],\exu/lsu/n59 [46]}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8098_o,_al_u8293_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8100|_al_u8099  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [57]}),
    .b({_al_u3514_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [57],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8100_o,\exu/alu_au/n31 [57]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8101|_al_u8437  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[57],ds1[39]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8101_o,_al_u8437_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*(D@C)))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(A*~(B*(D@C)))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1010001000101010),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1010001000101010),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8102|_al_u8971  (
    .a({_al_u8101_o,_al_u8970_o}),
    .b({rd_data_xor,rd_data_xor}),
    .c({ds1[57],ds1[13]}),
    .d({ds2[57],ds2[13]}),
    .f({_al_u8102_o,_al_u8971_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8104|_al_u8103  (
    .a({_al_u8100_o,and_clr}),
    .b({_al_u8102_o,rd_data_and}),
    .c({_al_u2855_o,ds1[57]}),
    .d({\exu/alu_au/n33 [57],ds2[57]}),
    .f({_al_u8104_o,\exu/alu_au/n33 [57]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000110010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8105|_al_u8107  (
    .a({open_n58210,\exu/n57 [57]}),
    .b({data_rd[57],_al_u2855_o}),
    .c({data_rd[58],_al_u8106_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [57],_al_u8107_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8106|_al_u8111  (
    .b({data_rd[57],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[56]}),
    .d({data_rd[56],\exu/n59_lutinv }),
    .f({_al_u8106_o,_al_u8111_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(~(C*~B)*~(D*~A))"),
    //.LUTG0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(~(C*~B)*~(D*~A))"),
    .INIT_LUTF0(16'b0000001111001111),
    .INIT_LUTF1(16'b1000101011001111),
    .INIT_LUTG0(16'b0000001111001111),
    .INIT_LUTG1(16'b1000101011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8110|_al_u8109  (
    .a({_al_u7979_o,open_n58261}),
    .b({_al_u8109_o,_al_u3224_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\biu/l1d_out [56]}),
    .d({\exu/lsu/n56 ,uncache_data[56]}),
    .f({_al_u8110_o,_al_u8109_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1101111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1101111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8112|exu/reg1_b56  (
    .a({_al_u7905_o,_al_u8112_o}),
    .b({_al_u7973_o,_al_u8114_o}),
    .c({_al_u8110_o,_al_u8120_o}),
    .clk(clk_pad),
    .d({_al_u8111_o,_al_u8123_o}),
    .sr(rst_pad),
    .f({_al_u8112_o,open_n58303}),
    .q({open_n58307,data_rd[56]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(B*A)))"),
    //.LUT1("(~C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000100000001111),
    .INIT_LUT1(16'b0000001000001111),
    .MODE("LOGIC"))
    \_al_u8114|_al_u8237  (
    .a({_al_u7995_o,_al_u7995_o}),
    .b({\exu/lsu/n59 [56],_al_u8236_o}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8114_o,_al_u8237_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8116|_al_u8115  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [56]}),
    .b({_al_u3522_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [56],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8116_o,\exu/alu_au/n31 [56]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8117|_al_u8415  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[56],ds1[40]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8117_o,_al_u8415_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*(D@C)))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1010001000101010),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8118|_al_u8934  (
    .a({_al_u8117_o,_al_u8933_o}),
    .b({rd_data_xor,rd_data_xor}),
    .c({ds1[56],ds1[14]}),
    .d({ds2[56],ds2[14]}),
    .f({_al_u8118_o,_al_u8934_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8120|_al_u8119  (
    .a({_al_u8116_o,and_clr}),
    .b({_al_u8118_o,rd_data_and}),
    .c({_al_u2855_o,ds1[56]}),
    .d({\exu/alu_au/n33 [56],ds2[56]}),
    .f({_al_u8120_o,\exu/alu_au/n33 [56]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110010001000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u8121|_al_u8123  (
    .a({open_n58414,\exu/n57 [56]}),
    .b({data_rd[56],_al_u2855_o}),
    .c({data_rd[57],_al_u8122_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [56],_al_u8123_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8122|_al_u8131  (
    .b({data_rd[56],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[55]}),
    .d({data_rd[55],\exu/n59_lutinv }),
    .f({_al_u8122_o,_al_u8131_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8125|_al_u8590  (
    .c({\exu/lsu/n56 ,_al_u7912_o}),
    .d({_al_u7979_o,_al_u7979_o}),
    .f({_al_u8125_o,_al_u8590_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8126|_al_u7905  (
    .a({_al_u7902_o,open_n58485}),
    .b({_al_u7971_o,\exu/n60_lutinv }),
    .c({\exu/lsu/n51 ,\exu/lsu/n51 }),
    .d({\exu/lsu/n53 ,_al_u7902_o}),
    .f({_al_u8126_o,_al_u7905_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~A*~(C*~B))"),
    //.LUT1("(C*~B*~D)"),
    .INIT_LUT0(16'b0100010100000000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"))
    \_al_u8128|_al_u8130  (
    .a({open_n58510,_al_u8128_o}),
    .b({_al_u7981_o,_al_u8129_o}),
    .c({_al_u8127_o,\exu/lsu/mux27_b56_sel_is_3_o }),
    .d({_al_u7980_o,\exu/n60_lutinv }),
    .f({_al_u8128_o,_al_u8130_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1100101000000000),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8129|_al_u7978  (
    .a({open_n58531,\biu/l1d_out [55]}),
    .b({uncache_data[55],uncache_data[55]}),
    .c({_al_u3224_o,_al_u3224_o}),
    .d({\biu/l1d_out [55],\exu/lsu/n8_lutinv }),
    .f({_al_u8129_o,_al_u7978_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*B*~A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1011111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8132|exu/reg1_b55  (
    .a({_al_u8125_o,_al_u8132_o}),
    .b({_al_u8126_o,_al_u8134_o}),
    .c({_al_u8130_o,_al_u8140_o}),
    .clk(clk_pad),
    .d({_al_u8131_o,_al_u8143_o}),
    .sr(rst_pad),
    .f({_al_u8132_o,open_n58569}),
    .q({open_n58573,data_rd[55]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b1100101000000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u8133|_al_u8422  (
    .a({uncache_data[63],\biu/l1d_out [55]}),
    .b({uncache_data[55],uncache_data[55]}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,_al_u3224_o}),
    .d({_al_u8127_o,\exu/lsu/n5_lutinv }),
    .f({_al_u8133_o,_al_u8422_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(B*A)))"),
    //.LUTF1("(~C*~(D*~(B*A)))"),
    //.LUTG0("(~C*~(D*~(B*A)))"),
    //.LUTG1("(~C*~(D*~(B*A)))"),
    .INIT_LUTF0(16'b0000100000001111),
    .INIT_LUTF1(16'b0000100000001111),
    .INIT_LUTG0(16'b0000100000001111),
    .INIT_LUTG1(16'b0000100000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8134|_al_u8203  (
    .a({_al_u7995_o,_al_u7995_o}),
    .b({_al_u8133_o,_al_u8202_o}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8134_o,_al_u8203_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8136|_al_u8135  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [55]}),
    .b({_al_u3530_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [55],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8136_o,\exu/alu_au/n31 [55]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u8137|_al_u8396  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[55],ds1[41]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8137_o,_al_u8396_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8138|_al_u3532  (
    .a({_al_u8137_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[55],ds1[55]}),
    .d({ds2[55],ds2[55]}),
    .f({_al_u8138_o,\exu/alu_au/n55 [55]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8140|_al_u8139  (
    .a({_al_u8136_o,and_clr}),
    .b({_al_u8138_o,rd_data_and}),
    .c({_al_u2855_o,ds1[55]}),
    .d({\exu/alu_au/n33 [55],ds2[55]}),
    .f({_al_u8140_o,\exu/alu_au/n33 [55]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110010001000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u8141|_al_u8143  (
    .a({open_n58704,\exu/n57 [55]}),
    .b({data_rd[55],_al_u2855_o}),
    .c({data_rd[56],_al_u8142_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [55],_al_u8143_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8142|_al_u8148  (
    .b({data_rd[55],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[54]}),
    .d({data_rd[54],\exu/n59_lutinv }),
    .f({_al_u8142_o,_al_u8148_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("(C*~(B*D))"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("(C*~(B*D))"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0011000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8145|_al_u8214  (
    .b({_al_u8127_o,_al_u8127_o}),
    .c({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .d({_al_u8011_o,_al_u8077_o}),
    .f({_al_u8145_o,_al_u8214_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b0000110000111111),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u8147|_al_u8146  (
    .b({_al_u8146_o,_al_u3224_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,uncache_data[54]}),
    .d({_al_u8145_o,\biu/l1d_out [54]}),
    .f({_al_u8147_o,_al_u8146_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8149|exu/reg1_b54  (
    .a({_al_u8125_o,_al_u8149_o}),
    .b({_al_u8126_o,_al_u8151_o}),
    .c({_al_u8147_o,_al_u8157_o}),
    .clk(clk_pad),
    .d({_al_u8148_o,_al_u8160_o}),
    .sr(rst_pad),
    .f({_al_u8149_o,open_n58808}),
    .q({open_n58812,data_rd[54]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(B*A)))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D*~(B*A)))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0000100000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000100000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8150|_al_u8151  (
    .a({uncache_data[62],_al_u7995_o}),
    .b({uncache_data[54],_al_u8150_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/c_stb_lutinv }),
    .d({_al_u8127_o,\exu/n59_lutinv }),
    .f({_al_u8150_o,_al_u8151_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8153|_al_u8152  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [54]}),
    .b({_al_u3538_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [54],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8153_o,\exu/alu_au/n31 [54]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8154|_al_u8336  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[54],ds1[44]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8154_o,_al_u8336_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8155|_al_u3540  (
    .a({_al_u8154_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[54],ds1[54]}),
    .d({ds2[54],ds2[54]}),
    .f({_al_u8155_o,\exu/alu_au/n55 [54]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8157|_al_u8156  (
    .a({_al_u8153_o,and_clr}),
    .b({_al_u8155_o,rd_data_and}),
    .c({_al_u2855_o,ds1[54]}),
    .d({\exu/alu_au/n33 [54],ds2[54]}),
    .f({_al_u8157_o,\exu/alu_au/n33 [54]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000110010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8158|_al_u8160  (
    .a({open_n58935,\exu/n57 [54]}),
    .b({data_rd[54],_al_u2855_o}),
    .c({data_rd[55],_al_u8159_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [54],_al_u8160_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8159|_al_u8166  (
    .b({data_rd[54],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[53]}),
    .d({data_rd[53],\exu/n59_lutinv }),
    .f({_al_u8159_o,_al_u8166_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~B*~D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"))
    \_al_u8162|_al_u8127  (
    .b({_al_u8028_o,open_n58988}),
    .c({_al_u8127_o,unsign}),
    .d({_al_u8027_o,\exu/lsu/n2_lutinv }),
    .f({_al_u8162_o,_al_u8127_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1111010100111111),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111010100111111),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8163|_al_u8471  (
    .a({open_n59009,uncache_data[53]}),
    .b({open_n59010,uncache_data[45]}),
    .c({_al_u3224_o,addr_ex[0]}),
    .d({uncache_data[53],addr_ex[1]}),
    .f({_al_u8163_o,_al_u8471_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~(~B*~A))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b0000111000000000),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8164|_al_u8464  (
    .a({open_n59035,\biu/l1d_out [53]}),
    .b({_al_u3224_o,_al_u3224_o}),
    .c({_al_u8163_o,_al_u8163_o}),
    .d({\biu/l1d_out [53],\exu/lsu/n5_lutinv }),
    .f({_al_u8164_o,_al_u8464_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUT1("(D*~A*~(C*B))"),
    .INIT_LUT0(16'b1010110000000000),
    .INIT_LUT1(16'b0001010100000000),
    .MODE("LOGIC"))
    \_al_u8165|_al_u8627  (
    .a({_al_u8162_o,_al_u8164_o}),
    .b({_al_u8164_o,_al_u8306_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,addr_ex[0]}),
    .d({\exu/n60_lutinv ,addr_ex[1]}),
    .f({_al_u8165_o,_al_u8627_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8167|exu/reg1_b53  (
    .a({_al_u8125_o,_al_u8167_o}),
    .b({_al_u8126_o,_al_u8169_o}),
    .c({_al_u8165_o,_al_u8175_o}),
    .clk(clk_pad),
    .d({_al_u8166_o,_al_u8178_o}),
    .sr(rst_pad),
    .f({_al_u8167_o,open_n59089}),
    .q({open_n59093,data_rd[53]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(B*A)))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0000100000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u8168|_al_u8169  (
    .a({uncache_data[61],_al_u7995_o}),
    .b({uncache_data[53],_al_u8168_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/c_stb_lutinv }),
    .d({_al_u8127_o,\exu/n59_lutinv }),
    .f({_al_u8168_o,_al_u8169_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8171|_al_u8170  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [53]}),
    .b({_al_u3546_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [53],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8171_o,\exu/alu_au/n31 [53]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u8172|_al_u8316  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[53],ds1[45]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8172_o,_al_u8316_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8173|_al_u3548  (
    .a({_al_u8172_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[53],ds1[53]}),
    .d({ds2[53],ds2[53]}),
    .f({_al_u8173_o,\exu/alu_au/n55 [53]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8175|_al_u8174  (
    .a({_al_u8171_o,and_clr}),
    .b({_al_u8173_o,rd_data_and}),
    .c({_al_u2855_o,ds1[53]}),
    .d({\exu/alu_au/n33 [53],ds2[53]}),
    .f({_al_u8175_o,\exu/alu_au/n33 [53]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000110010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8176|_al_u8178  (
    .a({open_n59204,\exu/n57 [53]}),
    .b({data_rd[53],_al_u2855_o}),
    .c({data_rd[54],_al_u8177_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [53],_al_u8178_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8177|_al_u8183  (
    .b({data_rd[53],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[52]}),
    .d({data_rd[52],\exu/n59_lutinv }),
    .f({_al_u8177_o,_al_u8183_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1100101000000000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1100101000000000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8180|_al_u8487  (
    .a({open_n59255,\biu/l1d_out [52]}),
    .b({uncache_data[52],uncache_data[52]}),
    .c({_al_u3224_o,_al_u3224_o}),
    .d({\biu/l1d_out [52],\exu/lsu/n5_lutinv }),
    .f({_al_u8180_o,_al_u8487_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b1100101000000000),
    .INIT_LUT1(16'b1100101000000000),
    .MODE("LOGIC"))
    \_al_u8181|_al_u8486  (
    .a({\biu/l1d_out [60],\biu/l1d_out [60]}),
    .b({uncache_data[60],uncache_data[60]}),
    .c({_al_u3224_o,_al_u3224_o}),
    .d({_al_u8127_o,\exu/lsu/n8_lutinv }),
    .f({_al_u8181_o,_al_u8486_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(D*~B*~(C*A))"),
    //.LUTG0("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(D*~B*~(C*A))"),
    .INIT_LUTF0(16'b1010110000000000),
    .INIT_LUTF1(16'b0001001100000000),
    .INIT_LUTG0(16'b1010110000000000),
    .INIT_LUTG1(16'b0001001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8182|_al_u8647  (
    .a({_al_u8180_o,_al_u8180_o}),
    .b({_al_u8181_o,_al_u8327_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,addr_ex[0]}),
    .d({\exu/n60_lutinv ,addr_ex[1]}),
    .f({_al_u8182_o,_al_u8647_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*B*~A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1011111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8184|exu/reg1_b52  (
    .a({_al_u8125_o,_al_u8184_o}),
    .b({_al_u8126_o,_al_u8186_o}),
    .c({_al_u8182_o,_al_u8192_o}),
    .clk(clk_pad),
    .d({_al_u8183_o,_al_u8195_o}),
    .sr(rst_pad),
    .f({_al_u8184_o,open_n59341}),
    .q({open_n59345,data_rd[52]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(B*A)))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0000100000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u8185|_al_u8186  (
    .a({uncache_data[60],_al_u7995_o}),
    .b({uncache_data[52],_al_u8185_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/c_stb_lutinv }),
    .d({_al_u8127_o,\exu/n59_lutinv }),
    .f({_al_u8185_o,_al_u8186_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8188|_al_u8187  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [52]}),
    .b({_al_u3554_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [52],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8188_o,\exu/alu_au/n31 [52]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u8189|_al_u8296  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[52],ds1[46]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8189_o,_al_u8296_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8190|_al_u3556  (
    .a({_al_u8189_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[52],ds1[52]}),
    .d({ds2[52],ds2[52]}),
    .f({_al_u8190_o,\exu/alu_au/n55 [52]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8192|_al_u8191  (
    .a({_al_u8188_o,and_clr}),
    .b({_al_u8190_o,rd_data_and}),
    .c({_al_u2855_o,ds1[52]}),
    .d({\exu/alu_au/n33 [52],ds2[52]}),
    .f({_al_u8192_o,\exu/alu_au/n33 [52]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110010001000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u8193|_al_u8195  (
    .a({open_n59448,\exu/n57 [52]}),
    .b({data_rd[52],_al_u2855_o}),
    .c({data_rd[53],_al_u8194_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [52],_al_u8195_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8194|_al_u8200  (
    .b({data_rd[52],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[51]}),
    .d({data_rd[51],\exu/n59_lutinv }),
    .f({_al_u8194_o,_al_u8200_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8198|_al_u8670  (
    .a({open_n59491,uncache_data[51]}),
    .b({_al_u3224_o,uncache_data[27]}),
    .c({\biu/l1d_out [51],addr_ex[0]}),
    .d({uncache_data[51],addr_ex[1]}),
    .f({_al_u8198_o,_al_u8670_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("(D*~(C*B))"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("(D*~(C*B))"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8199|_al_u8197  (
    .b({_al_u8198_o,_al_u8127_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/n60_lutinv }),
    .d({_al_u8197_o,_al_u8061_o}),
    .f({_al_u8199_o,_al_u8197_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*B*~A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1011111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8201|exu/reg1_b51  (
    .a({_al_u8125_o,_al_u8201_o}),
    .b({_al_u8126_o,_al_u8203_o}),
    .c({_al_u8199_o,_al_u8209_o}),
    .clk(clk_pad),
    .d({_al_u8200_o,_al_u8212_o}),
    .sr(rst_pad),
    .f({_al_u8201_o,open_n59559}),
    .q({open_n59563,data_rd[51]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u8202|_al_u8515  (
    .a({uncache_data[59],uncache_data[51]}),
    .b({uncache_data[51],uncache_data[43]}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,addr_ex[0]}),
    .d({_al_u8127_o,addr_ex[1]}),
    .f({_al_u8202_o,_al_u8515_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8205|_al_u8204  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [51]}),
    .b({_al_u3562_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [51],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8205_o,\exu/alu_au/n31 [51]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~B*~(C*D))"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~B*~(C*D))"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8206|_al_u8257  (
    .b({rd_data_or,rd_data_or}),
    .c({ds1[51],ds1[48]}),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8206_o,_al_u8257_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8207|_al_u3564  (
    .a({_al_u8206_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[51],ds1[51]}),
    .d({ds2[51],ds2[51]}),
    .f({_al_u8207_o,\exu/alu_au/n55 [51]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8209|_al_u8208  (
    .a({_al_u8205_o,and_clr}),
    .b({_al_u8207_o,rd_data_and}),
    .c({_al_u2855_o,ds1[51]}),
    .d({\exu/alu_au/n33 [51],ds2[51]}),
    .f({_al_u8209_o,\exu/alu_au/n33 [51]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110010001000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u8210|_al_u8212  (
    .a({open_n59674,\exu/n57 [51]}),
    .b({data_rd[51],_al_u2855_o}),
    .c({data_rd[52],_al_u8211_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [51],_al_u8212_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8211|_al_u8217  (
    .b({data_rd[51],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[50]}),
    .d({data_rd[50],\exu/n59_lutinv }),
    .f({_al_u8211_o,_al_u8217_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("(D*~(C*~B))"),
    .INIT_LUT0(16'b0000110000111111),
    .INIT_LUT1(16'b1100111100000000),
    .MODE("LOGIC"))
    \_al_u8216|_al_u8215  (
    .b({_al_u8215_o,_al_u3224_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,uncache_data[50]}),
    .d({_al_u8214_o,\biu/l1d_out [50]}),
    .f({_al_u8216_o,_al_u8215_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8218|exu/reg1_b50  (
    .a({_al_u8125_o,_al_u8218_o}),
    .b({_al_u8126_o,_al_u8220_o}),
    .c({_al_u8216_o,_al_u8226_o}),
    .clk(clk_pad),
    .d({_al_u8217_o,_al_u8229_o}),
    .sr(rst_pad),
    .f({_al_u8218_o,open_n59752}),
    .q({open_n59756,data_rd[50]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(B*A)))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~C*~(D*~(B*A)))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .INIT_LUTF0(16'b0000100000001111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0000100000001111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8219|_al_u8220  (
    .a({uncache_data[58],_al_u7995_o}),
    .b({uncache_data[50],_al_u8219_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/c_stb_lutinv }),
    .d({_al_u8127_o,\exu/n59_lutinv }),
    .f({_al_u8219_o,_al_u8220_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8222|_al_u8221  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [50]}),
    .b({_al_u3570_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [50],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8222_o,\exu/alu_au/n31 [50]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~B*~(C*D))"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0000001100110011),
    .MODE("LOGIC"))
    \_al_u8223|_al_u8240  (
    .b({rd_data_or,rd_data_or}),
    .c(ds1[50:49]),
    .d({rd_data_ds1,rd_data_ds1}),
    .f({_al_u8223_o,_al_u8240_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8224|_al_u3572  (
    .a({_al_u8223_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[50],ds1[50]}),
    .d({ds2[50],ds2[50]}),
    .f({_al_u8224_o,\exu/alu_au/n55 [50]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8226|_al_u8225  (
    .a({_al_u8222_o,and_clr}),
    .b({_al_u8224_o,rd_data_and}),
    .c({_al_u2855_o,ds1[50]}),
    .d({\exu/alu_au/n33 [50],ds2[50]}),
    .f({_al_u8226_o,\exu/alu_au/n33 [50]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000110010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8227|_al_u8229  (
    .a({open_n59875,\exu/n57 [50]}),
    .b({data_rd[50],_al_u2855_o}),
    .c({data_rd[51],_al_u8228_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [50],_al_u8229_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8228|_al_u8234  (
    .b({data_rd[50],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[49]}),
    .d({data_rd[49],\exu/n59_lutinv }),
    .f({_al_u8228_o,_al_u8234_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~A*~(C*~B))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0100010100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u8231|_al_u8233  (
    .a({open_n59926,_al_u8231_o}),
    .b({open_n59927,_al_u8232_o}),
    .c({_al_u8127_o,\exu/lsu/mux27_b56_sel_is_3_o }),
    .d({_al_u8093_o,\exu/n60_lutinv }),
    .f({_al_u8231_o,_al_u8233_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b0000001111001111),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b0000001111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8232|_al_u8707  (
    .a({open_n59948,uncache_data[49]}),
    .b({_al_u3224_o,uncache_data[33]}),
    .c({\biu/l1d_out [49],addr_ex[0]}),
    .d({uncache_data[49],addr_ex[1]}),
    .f({_al_u8232_o,_al_u8707_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8235|exu/reg1_b49  (
    .a({_al_u8125_o,_al_u8235_o}),
    .b({_al_u8126_o,_al_u8237_o}),
    .c({_al_u8233_o,_al_u8243_o}),
    .clk(clk_pad),
    .d({_al_u8234_o,_al_u8246_o}),
    .sr(rst_pad),
    .f({_al_u8235_o,open_n59986}),
    .q({open_n59990,data_rd[49]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u8236|_al_u8556  (
    .a({uncache_data[57],uncache_data[49]}),
    .b({uncache_data[49],uncache_data[41]}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,addr_ex[0]}),
    .d({_al_u8127_o,addr_ex[1]}),
    .f({_al_u8236_o,_al_u8556_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8239|_al_u8238  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [49]}),
    .b({_al_u3585_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [49],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8239_o,\exu/alu_au/n31 [49]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8241|_al_u3587  (
    .a({_al_u8240_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[49],ds1[49]}),
    .d({ds2[49],ds2[49]}),
    .f({_al_u8241_o,\exu/alu_au/n55 [49]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8243|_al_u8242  (
    .a({_al_u8239_o,and_clr}),
    .b({_al_u8241_o,rd_data_and}),
    .c({_al_u2855_o,ds1[49]}),
    .d({\exu/alu_au/n33 [49],ds2[49]}),
    .f({_al_u8243_o,\exu/alu_au/n33 [49]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000110010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8244|_al_u8246  (
    .a({open_n60079,\exu/n57 [49]}),
    .b({data_rd[49],_al_u2855_o}),
    .c({data_rd[50],_al_u8245_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [49],_al_u8246_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8245|_al_u8251  (
    .b({data_rd[49],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[48]}),
    .d({data_rd[48],\exu/n59_lutinv }),
    .f({_al_u8245_o,_al_u8251_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111010100111111),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111010100111111),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8249|_al_u8576  (
    .a({open_n60130,uncache_data[48]}),
    .b({_al_u3224_o,uncache_data[40]}),
    .c({uncache_data[48],addr_ex[0]}),
    .d({\biu/l1d_out [48],addr_ex[1]}),
    .f({_al_u8249_o,_al_u8576_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u8250|_al_u8248  (
    .b({_al_u8249_o,_al_u8127_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/n60_lutinv }),
    .d({_al_u8248_o,_al_u8109_o}),
    .f({_al_u8250_o,_al_u8248_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*B*~A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1011111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8252|exu/reg1_b48  (
    .a({_al_u8125_o,_al_u8252_o}),
    .b({_al_u8126_o,_al_u8254_o}),
    .c({_al_u8250_o,_al_u8260_o}),
    .clk(clk_pad),
    .d({_al_u8251_o,_al_u8263_o}),
    .sr(rst_pad),
    .f({_al_u8252_o,open_n60194}),
    .q({open_n60198,data_rd[48]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(B*A)))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b0000100000001111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u8253|_al_u8254  (
    .a({uncache_data[56],_al_u7995_o}),
    .b({uncache_data[48],_al_u8253_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,\exu/c_stb_lutinv }),
    .d({_al_u8127_o,\exu/n59_lutinv }),
    .f({_al_u8253_o,_al_u8254_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8256|_al_u8255  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [48]}),
    .b({_al_u3593_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [48],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8256_o,\exu/alu_au/n31 [48]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8258|_al_u3595  (
    .a({_al_u8257_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[48],ds1[48]}),
    .d({ds2[48],ds2[48]}),
    .f({_al_u8258_o,\exu/alu_au/n55 [48]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8260|_al_u8259  (
    .a({_al_u8256_o,and_clr}),
    .b({_al_u8258_o,rd_data_and}),
    .c({_al_u2855_o,ds1[48]}),
    .d({\exu/alu_au/n33 [48],ds2[48]}),
    .f({_al_u8260_o,\exu/alu_au/n33 [48]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110010001000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u8261|_al_u8263  (
    .a({open_n60279,\exu/n57 [48]}),
    .b({data_rd[48],_al_u2855_o}),
    .c({data_rd[49],_al_u8262_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [48],_al_u8263_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8262|_al_u8270  (
    .b({data_rd[48],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[47]}),
    .d({data_rd[47],\exu/n59_lutinv }),
    .f({_al_u8262_o,_al_u8270_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8266|_al_u8305  (
    .c({\exu/lsu/n2_lutinv ,\exu/lsu/n2_lutinv }),
    .d({_al_u8129_o,_al_u8164_o}),
    .f({_al_u8266_o,_al_u8305_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(C*~(D*~(~B*~A)))"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b0001000011110000),
    .MODE("LOGIC"))
    \_al_u8269|_al_u8268  (
    .a({_al_u8265_o,open_n60350}),
    .b({_al_u8266_o,\exu/lsu/mux27_b56_sel_is_3_o }),
    .c({_al_u8268_o,\exu/n60_lutinv }),
    .d({unsign,_al_u8267_o}),
    .f({_al_u8269_o,_al_u8268_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*B*~A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1011111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8271|exu/reg1_b47  (
    .a({_al_u8125_o,_al_u8271_o}),
    .b({_al_u8126_o,_al_u8274_o}),
    .c({_al_u8269_o,_al_u8280_o}),
    .clk(clk_pad),
    .d({_al_u8270_o,_al_u8283_o}),
    .sr(rst_pad),
    .f({_al_u8271_o,open_n60388}),
    .q({open_n60392,data_rd[47]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b0000101000001100),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b0000101000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8272|_al_u8428  (
    .a({uncache_data[63],uncache_data[63]}),
    .b({uncache_data[47],uncache_data[47]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u8272_o,_al_u8428_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*A)))"),
    //.LUTF1("(D*~(~A*~(C*B)))"),
    //.LUTG0("(~C*~(D*~(~B*A)))"),
    //.LUTG1("(D*~(~A*~(C*B)))"),
    .INIT_LUTF0(16'b0000001000001111),
    .INIT_LUTF1(16'b1110101000000000),
    .INIT_LUTG0(16'b0000001000001111),
    .INIT_LUTG1(16'b1110101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8273|_al_u8274  (
    .a({_al_u8272_o,_al_u7995_o}),
    .b({uncache_data[55],\exu/lsu/n59 [47]}),
    .c({\exu/lsu/n2_lutinv ,\exu/c_stb_lutinv }),
    .d({unsign,\exu/n59_lutinv }),
    .f({\exu/lsu/n59 [47],_al_u8274_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8276|_al_u8275  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [47]}),
    .b({_al_u3601_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [47],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8276_o,\exu/alu_au/n31 [47]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8278|_al_u8277  (
    .a({_al_u8277_o,open_n60461}),
    .b({rd_data_xor,rd_data_or}),
    .c({ds1[47],ds1[47]}),
    .d({ds2[47],rd_data_ds1}),
    .f({_al_u8278_o,_al_u8277_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8280|_al_u8279  (
    .a({_al_u8276_o,and_clr}),
    .b({_al_u8278_o,rd_data_and}),
    .c({_al_u2855_o,ds1[47]}),
    .d({\exu/alu_au/n33 [47],ds2[47]}),
    .f({_al_u8280_o,\exu/alu_au/n33 [47]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110010001000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u8281|_al_u8283  (
    .a({open_n60506,\exu/n57 [47]}),
    .b({data_rd[47],_al_u2855_o}),
    .c({data_rd[48],_al_u8282_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [47],_al_u8283_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8282|_al_u8289  (
    .b({data_rd[47],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[46]}),
    .d({data_rd[46],\exu/n59_lutinv }),
    .f({_al_u8282_o,_al_u8289_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b0000001111001111),
    .MODE("LOGIC"))
    \_al_u8286|_al_u8611  (
    .a({open_n60549,uncache_data[46]}),
    .b({_al_u3224_o,uncache_data[38]}),
    .c({\biu/l1d_out [46],addr_ex[0]}),
    .d({uncache_data[46],addr_ex[1]}),
    .f({_al_u8286_o,_al_u8611_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b1111010111001111),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u8288|_al_u8285  (
    .a({open_n60570,_al_u8011_o}),
    .b({_al_u8287_o,_al_u8146_o}),
    .c({unsign,addr_ex[0]}),
    .d({_al_u8285_o,addr_ex[1]}),
    .f({_al_u8288_o,_al_u8285_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8290|exu/reg1_b46  (
    .a({_al_u8125_o,_al_u8290_o}),
    .b({_al_u8126_o,_al_u8293_o}),
    .c({_al_u8288_o,_al_u8299_o}),
    .clk(clk_pad),
    .d({_al_u8289_o,_al_u8302_o}),
    .sr(rst_pad),
    .f({_al_u8290_o,open_n60604}),
    .q({open_n60608,data_rd[46]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(D*~(~A*~(C*B)))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b1110101000000000),
    .MODE("LOGIC"))
    \_al_u8292|_al_u8291  (
    .a({_al_u8291_o,uncache_data[62]}),
    .b({uncache_data[54],uncache_data[46]}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({\exu/lsu/n59 [46],_al_u8291_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8295|_al_u8294  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [46]}),
    .b({_al_u3609_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [46],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8295_o,\exu/alu_au/n31 [46]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8297|_al_u3611  (
    .a({_al_u8296_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[46],ds1[46]}),
    .d({ds2[46],ds2[46]}),
    .f({_al_u8297_o,\exu/alu_au/n55 [46]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8299|_al_u8298  (
    .a({_al_u8295_o,and_clr}),
    .b({_al_u8297_o,rd_data_and}),
    .c({_al_u2855_o,ds1[46]}),
    .d({\exu/alu_au/n33 [46],ds2[46]}),
    .f({_al_u8299_o,\exu/alu_au/n33 [46]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000110010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8300|_al_u8302  (
    .a({open_n60697,\exu/n57 [46]}),
    .b({data_rd[46],_al_u2855_o}),
    .c({data_rd[47],_al_u8301_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [46],_al_u8302_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8301|_al_u8309  (
    .b({data_rd[46],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[45]}),
    .d({data_rd[45],\exu/n59_lutinv }),
    .f({_al_u8301_o,_al_u8309_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*~(~B*~A)))"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("(C*~(D*~(~B*~A)))"),
    //.LUTG1("(C*~B*~D)"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b0001000011110000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8304|_al_u8308  (
    .a({open_n60748,_al_u8304_o}),
    .b({_al_u8028_o,_al_u8305_o}),
    .c({\exu/lsu/n5_lutinv ,_al_u8307_o}),
    .d({_al_u8027_o,unsign}),
    .f({_al_u8304_o,_al_u8308_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1100101000000000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1100101000000000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8306|_al_u8465  (
    .a({open_n60773,\biu/l1d_out [45]}),
    .b({uncache_data[45],uncache_data[45]}),
    .c({_al_u3224_o,_al_u3224_o}),
    .d({\biu/l1d_out [45],\exu/lsu/n2_lutinv }),
    .f({_al_u8306_o,_al_u8465_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(C*~(B*D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(C*~(B*D))"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b0011000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8307|_al_u8780  (
    .a({open_n60798,_al_u8306_o}),
    .b({\exu/lsu/mux27_b56_sel_is_3_o ,_al_u8779_o}),
    .c({\exu/n60_lutinv ,addr_ex[0]}),
    .d({_al_u8306_o,addr_ex[1]}),
    .f({_al_u8307_o,_al_u8780_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8310|exu/reg1_b45  (
    .a({_al_u8125_o,_al_u8310_o}),
    .b({_al_u8126_o,_al_u8313_o}),
    .c({_al_u8308_o,_al_u8319_o}),
    .clk(clk_pad),
    .d({_al_u8309_o,_al_u8322_o}),
    .sr(rst_pad),
    .f({_al_u8310_o,open_n60836}),
    .q({open_n60840,data_rd[45]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(D*~(~A*~(C*B)))"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(D*~(~A*~(C*B)))"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b1110101000000000),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b1110101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8312|_al_u8311  (
    .a({_al_u8311_o,uncache_data[61]}),
    .b({uncache_data[53],uncache_data[45]}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({\exu/lsu/n59 [45],_al_u8311_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8315|_al_u8314  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [45]}),
    .b({_al_u3617_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [45],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8315_o,\exu/alu_au/n31 [45]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8317|_al_u3619  (
    .a({_al_u8316_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[45],ds1[45]}),
    .d({ds2[45],ds2[45]}),
    .f({_al_u8317_o,\exu/alu_au/n55 [45]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8319|_al_u8318  (
    .a({_al_u8315_o,and_clr}),
    .b({_al_u8317_o,rd_data_and}),
    .c({_al_u2855_o,ds1[45]}),
    .d({\exu/alu_au/n33 [45],ds2[45]}),
    .f({_al_u8319_o,\exu/alu_au/n33 [45]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000110010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8320|_al_u8322  (
    .a({open_n60937,\exu/n57 [45]}),
    .b({data_rd[45],_al_u2855_o}),
    .c({data_rd[46],_al_u8321_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [45],_al_u8322_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8321|_al_u8329  (
    .b({data_rd[45],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[44]}),
    .d({data_rd[44],\exu/n59_lutinv }),
    .f({_al_u8321_o,_al_u8329_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("(D*~(~B*~(C*A)))"),
    .INIT_LUT0(16'b1100101000000000),
    .INIT_LUT1(16'b1110110000000000),
    .MODE("LOGIC"))
    \_al_u8325|_al_u8324  (
    .a({_al_u8180_o,\biu/l1d_out [60]}),
    .b({_al_u8324_o,uncache_data[60]}),
    .c({\exu/lsu/n2_lutinv ,_al_u3224_o}),
    .d({unsign,\exu/lsu/n5_lutinv }),
    .f({_al_u8325_o,_al_u8324_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u8326|_al_u8494  (
    .a({open_n61008,uncache_data[52]}),
    .b({open_n61009,uncache_data[44]}),
    .c({_al_u3224_o,addr_ex[0]}),
    .d({uncache_data[44],addr_ex[1]}),
    .f({_al_u8326_o,_al_u8494_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~(~B*~A))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b0000111000000000),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8327|_al_u8485  (
    .a({open_n61030,\biu/l1d_out [44]}),
    .b({_al_u3224_o,_al_u3224_o}),
    .c({_al_u8326_o,_al_u8326_o}),
    .d({\biu/l1d_out [44],\exu/lsu/n2_lutinv }),
    .f({_al_u8327_o,_al_u8485_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(D*~A*~(C*B))"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b0001010100000000),
    .MODE("LOGIC"))
    \_al_u8328|_al_u8799  (
    .a({_al_u8325_o,_al_u8327_o}),
    .b({_al_u8327_o,_al_u8798_o}),
    .c({\exu/lsu/mux27_b56_sel_is_3_o ,addr_ex[0]}),
    .d({\exu/n60_lutinv ,addr_ex[1]}),
    .f({_al_u8328_o,_al_u8799_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*B*~A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1011111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8330|exu/reg1_b44  (
    .a({_al_u8125_o,_al_u8330_o}),
    .b({_al_u8126_o,_al_u8333_o}),
    .c({_al_u8328_o,_al_u8339_o}),
    .clk(clk_pad),
    .d({_al_u8329_o,_al_u8342_o}),
    .sr(rst_pad),
    .f({_al_u8330_o,open_n61088}),
    .q({open_n61092,data_rd[44]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(D*~(~A*~(C*B)))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b1110101000000000),
    .MODE("LOGIC"))
    \_al_u8332|_al_u8331  (
    .a({_al_u8331_o,uncache_data[60]}),
    .b({uncache_data[52],uncache_data[44]}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({\exu/lsu/n59 [44],_al_u8331_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8335|_al_u8334  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [44]}),
    .b({_al_u3625_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [44],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8335_o,\exu/alu_au/n31 [44]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8337|_al_u3627  (
    .a({_al_u8336_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[44],ds1[44]}),
    .d({ds2[44],ds2[44]}),
    .f({_al_u8337_o,\exu/alu_au/n55 [44]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8339|_al_u8338  (
    .a({_al_u8335_o,and_clr}),
    .b({_al_u8337_o,rd_data_and}),
    .c({_al_u2855_o,ds1[44]}),
    .d({\exu/alu_au/n33 [44],ds2[44]}),
    .f({_al_u8339_o,\exu/alu_au/n33 [44]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110010001000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u8340|_al_u8342  (
    .a({open_n61173,\exu/n57 [44]}),
    .b({data_rd[44],_al_u2855_o}),
    .c({data_rd[45],_al_u8341_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [44],_al_u8342_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8341|_al_u8348  (
    .b({data_rd[44],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[43]}),
    .d({data_rd[43],\exu/n59_lutinv }),
    .f({_al_u8341_o,_al_u8348_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b1111101011001111),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u8346|_al_u8664  (
    .a({open_n61216,_al_u8345_o}),
    .b({\exu/lsu/mux27_b56_sel_is_3_o ,_al_u8508_o}),
    .c({\exu/n60_lutinv ,addr_ex[0]}),
    .d({_al_u8345_o,addr_ex[1]}),
    .f({_al_u8346_o,_al_u8664_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b1111101000111111),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u8347|_al_u8344  (
    .a({open_n61237,_al_u8061_o}),
    .b({_al_u8346_o,_al_u8198_o}),
    .c({unsign,addr_ex[0]}),
    .d({_al_u8344_o,addr_ex[1]}),
    .f({_al_u8347_o,_al_u8344_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*B*~A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1011111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8349|exu/reg1_b43  (
    .a({_al_u8125_o,_al_u8349_o}),
    .b({_al_u8126_o,_al_u8352_o}),
    .c({_al_u8347_o,_al_u8358_o}),
    .clk(clk_pad),
    .d({_al_u8348_o,_al_u8361_o}),
    .sr(rst_pad),
    .f({_al_u8349_o,open_n61275}),
    .q({open_n61279,data_rd[43]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(D*~(~A*~(C*B)))"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(D*~(~A*~(C*B)))"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b1110101000000000),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b1110101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8351|_al_u8350  (
    .a({_al_u8350_o,uncache_data[59]}),
    .b({uncache_data[51],uncache_data[43]}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({\exu/lsu/n59 [43],_al_u8350_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8354|_al_u8353  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [43]}),
    .b({_al_u3633_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [43],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8354_o,\exu/alu_au/n31 [43]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8356|_al_u8355  (
    .a({_al_u8355_o,open_n61324}),
    .b({rd_data_xor,rd_data_or}),
    .c({ds1[43],ds1[43]}),
    .d({ds2[43],rd_data_ds1}),
    .f({_al_u8356_o,_al_u8355_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8358|_al_u8357  (
    .a({_al_u8354_o,and_clr}),
    .b({_al_u8356_o,rd_data_and}),
    .c({_al_u2855_o,ds1[43]}),
    .d({\exu/alu_au/n33 [43],ds2[43]}),
    .f({_al_u8358_o,\exu/alu_au/n33 [43]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110010001000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u8359|_al_u8361  (
    .a({open_n61369,\exu/n57 [43]}),
    .b({data_rd[43],_al_u2855_o}),
    .c({data_rd[44],_al_u8360_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [43],_al_u8361_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8360|_al_u8367  (
    .b({data_rd[43],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[42]}),
    .d({data_rd[42],\exu/n59_lutinv }),
    .f({_al_u8360_o,_al_u8367_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(C*~(B*~D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(C*~(B*~D))"),
    .INIT_LUTF0(16'b1111101000111111),
    .INIT_LUTF1(16'b1111000000110000),
    .INIT_LUTG0(16'b1111101000111111),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8365|_al_u8683  (
    .a({open_n61412,_al_u8364_o}),
    .b({\exu/lsu/mux27_b56_sel_is_3_o ,_al_u8531_o}),
    .c({\exu/n60_lutinv ,addr_ex[0]}),
    .d({_al_u8364_o,addr_ex[1]}),
    .f({_al_u8365_o,_al_u8683_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b1111101011001111),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b1111101011001111),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8366|_al_u8363  (
    .a({open_n61437,_al_u8077_o}),
    .b({_al_u8365_o,_al_u8215_o}),
    .c({unsign,addr_ex[0]}),
    .d({_al_u8363_o,addr_ex[1]}),
    .f({_al_u8366_o,_al_u8363_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8368|exu/reg1_b42  (
    .a({_al_u8125_o,_al_u8368_o}),
    .b({_al_u8126_o,_al_u8371_o}),
    .c({_al_u8366_o,_al_u8377_o}),
    .clk(clk_pad),
    .d({_al_u8367_o,_al_u8380_o}),
    .sr(rst_pad),
    .f({_al_u8368_o,open_n61475}),
    .q({open_n61479,data_rd[42]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(D*~(~A*~(C*B)))"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(D*~(~A*~(C*B)))"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b1110101000000000),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b1110101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8370|_al_u8369  (
    .a({_al_u8369_o,uncache_data[58]}),
    .b({uncache_data[50],uncache_data[42]}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({\exu/lsu/n59 [42],_al_u8369_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8373|_al_u8372  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [42]}),
    .b({_al_u3641_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [42],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8373_o,\exu/alu_au/n31 [42]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*D))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b0000001100110011),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8375|_al_u8374  (
    .a({_al_u8374_o,open_n61528}),
    .b({rd_data_xor,rd_data_or}),
    .c({ds1[42],ds1[42]}),
    .d({ds2[42],rd_data_ds1}),
    .f({_al_u8375_o,_al_u8374_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8377|_al_u8376  (
    .a({_al_u8373_o,and_clr}),
    .b({_al_u8375_o,rd_data_and}),
    .c({_al_u2855_o,ds1[42]}),
    .d({\exu/alu_au/n33 [42],ds2[42]}),
    .f({_al_u8377_o,\exu/alu_au/n33 [42]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000110010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8378|_al_u8380  (
    .a({open_n61573,\exu/n57 [42]}),
    .b({data_rd[42],_al_u2855_o}),
    .c({data_rd[43],_al_u8379_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [42],_al_u8380_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8379|_al_u8386  (
    .b({data_rd[42],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[41]}),
    .d({data_rd[41],\exu/n59_lutinv }),
    .f({_al_u8379_o,_al_u8386_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b1111010111001111),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b1111010111001111),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8385|_al_u8382  (
    .a({open_n61624,_al_u8093_o}),
    .b({_al_u8384_o,_al_u8232_o}),
    .c({unsign,addr_ex[0]}),
    .d({_al_u8382_o,addr_ex[1]}),
    .f({_al_u8385_o,_al_u8382_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111101111110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8387|exu/reg1_b41  (
    .a({_al_u8125_o,_al_u8387_o}),
    .b({_al_u8126_o,_al_u8390_o}),
    .c({_al_u8385_o,_al_u8393_o}),
    .clk(clk_pad),
    .d({_al_u8386_o,_al_u8399_o}),
    .sr(rst_pad),
    .f({_al_u8387_o,open_n61662}),
    .q({open_n61666,data_rd[41]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(D*~(~A*~(C*B)))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b1110101000000000),
    .MODE("LOGIC"))
    \_al_u8389|_al_u8388  (
    .a({_al_u8388_o,uncache_data[57]}),
    .b({uncache_data[49],uncache_data[41]}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({\exu/lsu/n59 [41],_al_u8388_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b0000000011100100),
    .MODE("LOGIC"))
    \_al_u8391|_al_u8393  (
    .a({\exu/mux27_b32_sel_is_1_o ,open_n61687}),
    .b({data_rd[41],_al_u2855_o}),
    .c({data_rd[42],_al_u8392_o}),
    .d({shift_l,_al_u8391_o}),
    .f({_al_u8391_o,_al_u8393_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b1100101000000000),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b1100101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8392|_al_u8405  (
    .a({data_rd[40],open_n61708}),
    .b({data_rd[41],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[40]}),
    .d({shift_l,\exu/n59_lutinv }),
    .f({_al_u8392_o,_al_u8405_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8395|_al_u8394  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [41]}),
    .b({_al_u3649_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [41],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8395_o,\exu/alu_au/n31 [41]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8397|_al_u3651  (
    .a({_al_u8396_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[41],ds1[41]}),
    .d({ds2[41],ds2[41]}),
    .f({_al_u8397_o,\exu/alu_au/n55 [41]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8399|_al_u8398  (
    .a({_al_u8395_o,and_clr}),
    .b({_al_u8397_o,rd_data_and}),
    .c({_al_u2855_o,ds1[41]}),
    .d({\exu/alu_au/n33 [41],ds2[41]}),
    .f({_al_u8399_o,\exu/alu_au/n33 [41]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b0000001111001111),
    .MODE("LOGIC"))
    \_al_u8402|_al_u8725  (
    .a({open_n61805,uncache_data[40]}),
    .b({_al_u3224_o,uncache_data[24]}),
    .c({\biu/l1d_out [40],addr_ex[0]}),
    .d({uncache_data[40],addr_ex[1]}),
    .f({_al_u8402_o,_al_u8725_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(B*~(C*~D))"),
    .INIT_LUT0(16'b1111101000111111),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"))
    \_al_u8404|_al_u8401  (
    .a({open_n61826,_al_u8109_o}),
    .b({_al_u8403_o,_al_u8249_o}),
    .c({unsign,addr_ex[0]}),
    .d({_al_u8401_o,addr_ex[1]}),
    .f({_al_u8404_o,_al_u8401_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D*~(B*~A)))"),
    //.LUTF1("(D*~(C*B*~A))"),
    //.LUTG0("~(~C*~(D*~(B*~A)))"),
    //.LUTG1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101111110000),
    .INIT_LUTF1(16'b1011111100000000),
    .INIT_LUTG0(16'b1111101111110000),
    .INIT_LUTG1(16'b1011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8406|exu/reg1_b40  (
    .a({_al_u8125_o,_al_u8406_o}),
    .b({_al_u8126_o,_al_u8409_o}),
    .c({_al_u8404_o,_al_u8412_o}),
    .clk(clk_pad),
    .d({_al_u8405_o,_al_u8418_o}),
    .sr(rst_pad),
    .f({_al_u8406_o,open_n61864}),
    .q({open_n61868,data_rd[40]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(D*~(~A*~(C*B)))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b1110101000000000),
    .MODE("LOGIC"))
    \_al_u8408|_al_u8407  (
    .a({_al_u8407_o,uncache_data[56]}),
    .b({uncache_data[48],uncache_data[40]}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({\exu/lsu/n59 [40],_al_u8407_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*~D))"),
    //.LUTF1("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    //.LUTG0("(B*~(~C*~D))"),
    //.LUTG1("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT_LUTF0(16'b1100110011000000),
    .INIT_LUTF1(16'b0000000011100100),
    .INIT_LUTG0(16'b1100110011000000),
    .INIT_LUTG1(16'b0000000011100100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8410|_al_u8412  (
    .a({\exu/mux27_b32_sel_is_1_o ,open_n61889}),
    .b({data_rd[40],_al_u2855_o}),
    .c({data_rd[41],_al_u8411_o}),
    .d({shift_l,_al_u8410_o}),
    .f({_al_u8410_o,_al_u8412_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b1100101000000000),
    .MODE("LOGIC"))
    \_al_u8411|_al_u8426  (
    .a({data_rd[39],open_n61914}),
    .b({data_rd[40],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[39]}),
    .d({shift_l,\exu/n59_lutinv }),
    .f({_al_u8411_o,_al_u8426_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8414|_al_u8413  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [40]}),
    .b({_al_u3657_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [40],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8414_o,\exu/alu_au/n31 [40]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8416|_al_u3659  (
    .a({_al_u8415_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[40],ds1[40]}),
    .d({ds2[40],ds2[40]}),
    .f({_al_u8416_o,\exu/alu_au/n55 [40]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8418|_al_u8417  (
    .a({_al_u8414_o,and_clr}),
    .b({_al_u8416_o,rd_data_and}),
    .c({_al_u2855_o,ds1[40]}),
    .d({\exu/alu_au/n33 [40],ds2[40]}),
    .f({_al_u8418_o,\exu/alu_au/n33 [40]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~A)*~(B)*~(D)+~(C*~A)*B*~(D)+~(~(C*~A))*B*D+~(C*~A)*B*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~(C*~A)*~(B)*~(D)+~(C*~A)*B*~(D)+~(~(C*~A))*B*D+~(C*~A)*B*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b1100110010101111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100110010101111),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8424|_al_u8425  (
    .a({_al_u8420_o,_al_u7979_o}),
    .b({_al_u8421_o,_al_u8424_o}),
    .c({_al_u8422_o,ex_size[2]}),
    .d({_al_u8423_o,unsign}),
    .f({_al_u8424_o,_al_u8425_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D*~(B*~A)))"),
    //.LUTF1("(D*~(C*~B*A))"),
    //.LUTG0("~(~C*~(D*~(B*~A)))"),
    //.LUTG1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101111110000),
    .INIT_LUTF1(16'b1101111100000000),
    .INIT_LUTG0(16'b1111101111110000),
    .INIT_LUTG1(16'b1101111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8427|exu/reg1_b39  (
    .a({_al_u7905_o,_al_u8427_o}),
    .b({_al_u7973_o,_al_u8431_o}),
    .c({_al_u8425_o,_al_u8434_o}),
    .clk(clk_pad),
    .d({_al_u8426_o,_al_u8440_o}),
    .sr(rst_pad),
    .f({_al_u8427_o,open_n62036}),
    .q({open_n62040,data_rd[39]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(A*~(D*~(~C*~B)))"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(A*~(D*~(~C*~B)))"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b0000001010101010),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b0000001010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8430|_al_u8429  (
    .a({_al_u7995_o,uncache_data[55]}),
    .b({_al_u8428_o,uncache_data[39]}),
    .c({_al_u8429_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8430_o,_al_u8429_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~D))"),
    //.LUT1("(~B*~(C*~D))"),
    .INIT_LUT0(16'b0011001100000011),
    .INIT_LUT1(16'b0011001100000011),
    .MODE("LOGIC"))
    \_al_u8431|_al_u8579  (
    .b({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .c({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .d({_al_u8430_o,_al_u8578_o}),
    .f({_al_u8431_o,_al_u8579_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*~D))"),
    //.LUTF1("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    //.LUTG0("(B*~(~C*~D))"),
    //.LUTG1("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT_LUTF0(16'b1100110011000000),
    .INIT_LUTF1(16'b0000000011100100),
    .INIT_LUTG0(16'b1100110011000000),
    .INIT_LUTG1(16'b0000000011100100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8432|_al_u8434  (
    .a({\exu/mux27_b32_sel_is_1_o ,open_n62087}),
    .b({data_rd[39],_al_u2855_o}),
    .c({data_rd[40],_al_u8433_o}),
    .d({shift_l,_al_u8432_o}),
    .f({_al_u8432_o,_al_u8434_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b1100101000000000),
    .MODE("LOGIC"))
    \_al_u8433|_al_u8447  (
    .a({data_rd[38],open_n62112}),
    .b({data_rd[39],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[38]}),
    .d({shift_l,\exu/n59_lutinv }),
    .f({_al_u8433_o,_al_u8447_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8436|_al_u8435  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [39]}),
    .b({_al_u3672_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [39],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8436_o,\exu/alu_au/n31 [39]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8438|_al_u3674  (
    .a({_al_u8437_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[39],ds1[39]}),
    .d({ds2[39],ds2[39]}),
    .f({_al_u8438_o,\exu/alu_au/n55 [39]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8440|_al_u8439  (
    .a({_al_u8436_o,and_clr}),
    .b({_al_u8438_o,rd_data_and}),
    .c({_al_u2855_o,ds1[39]}),
    .d({\exu/alu_au/n33 [39],ds2[39]}),
    .f({_al_u8440_o,\exu/alu_au/n33 [39]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~D))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~(B*~D))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8443|_al_u8287  (
    .b({open_n62199,\exu/lsu/mux27_b56_sel_is_3_o }),
    .c({_al_u8127_o,\exu/n60_lutinv }),
    .d({_al_u8286_o,_al_u8286_o}),
    .f({_al_u8443_o,_al_u8287_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(C*~(B*D))"),
    //.LUTG0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(C*~(B*D))"),
    .INIT_LUTF0(16'b0000000010101100),
    .INIT_LUTF1(16'b0011000011110000),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b0011000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8445|_al_u8606  (
    .a({open_n62224,_al_u8444_o}),
    .b({\exu/lsu/mux27_b56_sel_is_3_o ,_al_u8605_o}),
    .c({\exu/n60_lutinv ,addr_ex[0]}),
    .d({_al_u8444_o,addr_ex[1]}),
    .f({_al_u8445_o,_al_u8606_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    //.LUT1("(C*~B*~(D*A))"),
    .INIT_LUT0(16'b1010001100000000),
    .INIT_LUT1(16'b0001000000110000),
    .MODE("LOGIC"))
    \_al_u8446|_al_u8442  (
    .a({_al_u8442_o,_al_u8011_o}),
    .b({_al_u8443_o,_al_u8146_o}),
    .c({_al_u8445_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8446_o,_al_u8442_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8448|exu/reg1_b38  (
    .a({_al_u8125_o,_al_u8448_o}),
    .b({_al_u8126_o,_al_u8452_o}),
    .c({_al_u8446_o,_al_u8458_o}),
    .clk(clk_pad),
    .d({_al_u8447_o,_al_u8461_o}),
    .sr(rst_pad),
    .f({_al_u8448_o,open_n62282}),
    .q({open_n62286,data_rd[38]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(A*~(D*~(C*B)))"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b1000000010101010),
    .MODE("LOGIC"))
    \_al_u8451|_al_u8450  (
    .a({_al_u7995_o,uncache_data[54]}),
    .b({_al_u8449_o,uncache_data[46]}),
    .c({_al_u8450_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8451_o,_al_u8450_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~D))"),
    //.LUT1("(~B*~(C*~D))"),
    .INIT_LUT0(16'b0011001100000011),
    .INIT_LUT1(16'b0011001100000011),
    .MODE("LOGIC"))
    \_al_u8452|_al_u8559  (
    .b({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .c({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .d({_al_u8451_o,_al_u8558_o}),
    .f({_al_u8452_o,_al_u8559_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8454|_al_u8453  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [38]}),
    .b({_al_u3680_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [38],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8454_o,\exu/alu_au/n31 [38]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8456|_al_u3682  (
    .a({_al_u8455_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[38],ds1[38]}),
    .d({ds2[38],ds2[38]}),
    .f({_al_u8456_o,\exu/alu_au/n55 [38]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8458|_al_u8457  (
    .a({_al_u8454_o,and_clr}),
    .b({_al_u8456_o,rd_data_and}),
    .c({_al_u2855_o,ds1[38]}),
    .d({\exu/alu_au/n33 [38],ds2[38]}),
    .f({_al_u8458_o,\exu/alu_au/n33 [38]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110001000100),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000110001000100),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8459|_al_u8461  (
    .a({open_n62397,_al_u8459_o}),
    .b({data_rd[38],_al_u2855_o}),
    .c({data_rd[39],_al_u8460_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({_al_u8459_o,_al_u8461_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8460|_al_u8469  (
    .b({data_rd[38],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[37]}),
    .d({data_rd[37],\exu/n59_lutinv }),
    .f({_al_u8460_o,_al_u8469_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~A)*~(B)*~(D)+~(C*~A)*B*~(D)+~(~(C*~A))*B*D+~(C*~A)*B*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~(C*~A)*~(B)*~(D)+~(C*~A)*B*~(D)+~(~(C*~A))*B*D+~(C*~A)*B*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b1100110010101111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100110010101111),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8467|_al_u8468  (
    .a({_al_u8463_o,_al_u7979_o}),
    .b({_al_u8464_o,_al_u8467_o}),
    .c({_al_u8465_o,ex_size[2]}),
    .d({_al_u8466_o,unsign}),
    .f({_al_u8467_o,_al_u8468_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1101111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8470|exu/reg1_b37  (
    .a({_al_u7905_o,_al_u8470_o}),
    .b({_al_u7973_o,_al_u8474_o}),
    .c({_al_u8468_o,_al_u8480_o}),
    .clk(clk_pad),
    .d({_al_u8469_o,_al_u8483_o}),
    .sr(rst_pad),
    .f({_al_u8470_o,open_n62485}),
    .q({open_n62489,data_rd[37]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(A*~(D*~(C*B)))"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b1000000010101010),
    .MODE("LOGIC"))
    \_al_u8473|_al_u8472  (
    .a({_al_u7995_o,uncache_data[61]}),
    .b({_al_u8471_o,uncache_data[37]}),
    .c({_al_u8472_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8473_o,_al_u8472_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8474|_al_u8539  (
    .b({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .c({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .d({_al_u8473_o,_al_u8538_o}),
    .f({_al_u8474_o,_al_u8539_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8476|_al_u8475  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [37]}),
    .b({_al_u3688_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [37],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8476_o,\exu/alu_au/n31 [37]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8478|_al_u3690  (
    .a({_al_u8477_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[37],ds1[37]}),
    .d({ds2[37],ds2[37]}),
    .f({_al_u8478_o,\exu/alu_au/n55 [37]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8480|_al_u8479  (
    .a({_al_u8476_o,and_clr}),
    .b({_al_u8478_o,rd_data_and}),
    .c({_al_u2855_o,ds1[37]}),
    .d({\exu/alu_au/n33 [37],ds2[37]}),
    .f({_al_u8480_o,\exu/alu_au/n33 [37]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"))
    \_al_u8481|_al_u8483  (
    .a({open_n62608,_al_u8481_o}),
    .b({data_rd[37],_al_u2855_o}),
    .c({data_rd[38],_al_u8482_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({_al_u8481_o,_al_u8483_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8482|_al_u8492  (
    .b({data_rd[37],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[36]}),
    .d({data_rd[36],\exu/n59_lutinv }),
    .f({_al_u8482_o,_al_u8492_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(~B*D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*~(~B*D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000110000001111),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000110000001111),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8488|_al_u8267  (
    .b({open_n62657,_al_u3224_o}),
    .c({_al_u3224_o,_al_u7974_o}),
    .d({uncache_data[36],\biu/l1d_out [47]}),
    .f({_al_u8488_o,_al_u8267_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTF1("(D*~(~C*~(~B*A)))"),
    //.LUTG0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG1("(D*~(~C*~(~B*A)))"),
    .INIT_LUTF0(16'b1011000010000000),
    .INIT_LUTF1(16'b1111001000000000),
    .INIT_LUTG0(16'b1011000010000000),
    .INIT_LUTG1(16'b1111001000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8489|_al_u8904  (
    .a({\biu/l1d_out [36],uncache_data[6]}),
    .b({_al_u3224_o,_al_u3224_o}),
    .c({_al_u8488_o,\exu/lsu/n0_lutinv }),
    .d({\exu/lsu/n0_lutinv ,\biu/l1d_out [6]}),
    .f({_al_u8489_o,_al_u8904_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~A)*~(B)*~(D)+~(C*~A)*B*~(D)+~(~(C*~A))*B*D+~(C*~A)*B*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b1100110010101111),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u8490|_al_u8491  (
    .a({_al_u8485_o,_al_u7979_o}),
    .b({_al_u8486_o,_al_u8490_o}),
    .c({_al_u8487_o,ex_size[2]}),
    .d({_al_u8489_o,unsign}),
    .f({_al_u8490_o,_al_u8491_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1101111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1101111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8493|exu/reg1_b36  (
    .a({_al_u7905_o,_al_u8493_o}),
    .b({_al_u7973_o,_al_u8497_o}),
    .c({_al_u8491_o,_al_u8503_o}),
    .clk(clk_pad),
    .d({_al_u8492_o,_al_u8506_o}),
    .sr(rst_pad),
    .f({_al_u8493_o,open_n62743}),
    .q({open_n62747,data_rd[36]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(A*~(D*~(C*B)))"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b1000000010101010),
    .MODE("LOGIC"))
    \_al_u8496|_al_u8495  (
    .a({_al_u7995_o,uncache_data[60]}),
    .b({_al_u8494_o,uncache_data[36]}),
    .c({_al_u8495_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8496_o,_al_u8495_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8497|_al_u8518  (
    .b({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .c({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .d({_al_u8496_o,_al_u8517_o}),
    .f({_al_u8497_o,_al_u8518_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8499|_al_u8498  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [36]}),
    .b({_al_u3696_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [36],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8499_o,\exu/alu_au/n31 [36]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8501|_al_u3698  (
    .a({_al_u8500_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[36],ds1[36]}),
    .d({ds2[36],ds2[36]}),
    .f({_al_u8501_o,\exu/alu_au/n55 [36]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8503|_al_u8502  (
    .a({_al_u8499_o,and_clr}),
    .b({_al_u8501_o,rd_data_and}),
    .c({_al_u2855_o,ds1[36]}),
    .d({\exu/alu_au/n33 [36],ds2[36]}),
    .f({_al_u8503_o,\exu/alu_au/n33 [36]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000110010001000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u8504|_al_u8506  (
    .a({open_n62854,\exu/n57 [36]}),
    .b({data_rd[36],_al_u2855_o}),
    .c({data_rd[37],_al_u8505_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [36],_al_u8506_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8505|_al_u8513  (
    .b({data_rd[36],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[35]}),
    .d({data_rd[35],\exu/n59_lutinv }),
    .f({_al_u8505_o,_al_u8513_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000110000111111),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000110000111111),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8509|_al_u8508  (
    .b({open_n62899,_al_u3224_o}),
    .c({\exu/lsu/n0_lutinv ,uncache_data[35]}),
    .d({_al_u8508_o,\biu/l1d_out [35]}),
    .f({_al_u8509_o,_al_u8508_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(B*~D))"),
    //.LUTG0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(B*~D))"),
    .INIT_LUTF0(16'b0000001111001111),
    .INIT_LUTF1(16'b1111000000110000),
    .INIT_LUTG0(16'b0000001111001111),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8511|_al_u8345  (
    .b({_al_u8127_o,_al_u3224_o}),
    .c({\exu/n60_lutinv ,\biu/l1d_out [43]}),
    .d({_al_u8345_o,uncache_data[43]}),
    .f({_al_u8511_o,_al_u8345_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    //.LUTF1("(C*~(D*~(~B*~A)))"),
    //.LUTG0("(D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    //.LUTG1("(C*~(D*~(~B*~A)))"),
    .INIT_LUTF0(16'b0101110000000000),
    .INIT_LUTF1(16'b0001000011110000),
    .INIT_LUTG0(16'b0101110000000000),
    .INIT_LUTG1(16'b0001000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8512|_al_u8510  (
    .a({_al_u8509_o,_al_u8061_o}),
    .b({_al_u8510_o,_al_u8198_o}),
    .c({_al_u8511_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8512_o,_al_u8510_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D*~(B*~A)))"),
    //.LUTF1("(D*~(C*B*~A))"),
    //.LUTG0("~(~C*~(D*~(B*~A)))"),
    //.LUTG1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101111110000),
    .INIT_LUTF1(16'b1011111100000000),
    .INIT_LUTG0(16'b1111101111110000),
    .INIT_LUTG1(16'b1011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8514|exu/reg1_b35  (
    .a({_al_u8125_o,_al_u8514_o}),
    .b({_al_u8126_o,_al_u8518_o}),
    .c({_al_u8512_o,_al_u8521_o}),
    .clk(clk_pad),
    .d({_al_u8513_o,_al_u8527_o}),
    .sr(rst_pad),
    .f({_al_u8514_o,open_n62991}),
    .q({open_n62995,data_rd[35]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(A*~(D*~(C*B)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(A*~(D*~(C*B)))"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b1000000010101010),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b1000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8517|_al_u8516  (
    .a({_al_u7995_o,uncache_data[59]}),
    .b({_al_u8515_o,uncache_data[35]}),
    .c({_al_u8516_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8517_o,_al_u8516_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b0000000011100100),
    .MODE("LOGIC"))
    \_al_u8519|_al_u8521  (
    .a({\exu/mux27_b32_sel_is_1_o ,open_n63020}),
    .b({data_rd[35],_al_u2855_o}),
    .c({data_rd[36],_al_u8520_o}),
    .d({shift_l,_al_u8519_o}),
    .f({_al_u8519_o,_al_u8521_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b1100101000000000),
    .MODE("LOGIC"))
    \_al_u8520|_al_u8534  (
    .a({data_rd[34],open_n63041}),
    .b({data_rd[35],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[34]}),
    .d({shift_l,\exu/n59_lutinv }),
    .f({_al_u8520_o,_al_u8534_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8523|_al_u8522  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [35]}),
    .b({_al_u3704_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [35],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8523_o,\exu/alu_au/n31 [35]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8525|_al_u3706  (
    .a({_al_u8524_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[35],ds1[35]}),
    .d({ds2[35],ds2[35]}),
    .f({_al_u8525_o,\exu/alu_au/n55 [35]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8527|_al_u8526  (
    .a({_al_u8523_o,and_clr}),
    .b({_al_u8525_o,rd_data_and}),
    .c({_al_u2855_o,ds1[35]}),
    .d({\exu/alu_au/n33 [35],ds2[35]}),
    .f({_al_u8527_o,\exu/alu_au/n33 [35]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000001111001111),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001111001111),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8530|_al_u8364  (
    .b({open_n63128,_al_u3224_o}),
    .c({_al_u8127_o,\biu/l1d_out [42]}),
    .d({_al_u8364_o,uncache_data[42]}),
    .f({_al_u8530_o,_al_u8364_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*D))"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b0011000011110000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u8531|_al_u8532  (
    .b({_al_u3224_o,\exu/lsu/mux27_b56_sel_is_3_o }),
    .c({\biu/l1d_out [34],\exu/n60_lutinv }),
    .d({uncache_data[34],_al_u8531_o}),
    .f({_al_u8531_o,_al_u8532_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(C*~B*~(D*A))"),
    //.LUTG0("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(C*~B*~(D*A))"),
    .INIT_LUTF0(16'b0101001100000000),
    .INIT_LUTF1(16'b0001000000110000),
    .INIT_LUTG0(16'b0101001100000000),
    .INIT_LUTG1(16'b0001000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8533|_al_u8529  (
    .a({_al_u8529_o,_al_u8077_o}),
    .b({_al_u8530_o,_al_u8215_o}),
    .c({_al_u8532_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8533_o,_al_u8529_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(D*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111101111110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8535|exu/reg1_b34  (
    .a({_al_u8125_o,_al_u8535_o}),
    .b({_al_u8126_o,_al_u8539_o}),
    .c({_al_u8533_o,_al_u8542_o}),
    .clk(clk_pad),
    .d({_al_u8534_o,_al_u8548_o}),
    .sr(rst_pad),
    .f({_al_u8535_o,open_n63212}),
    .q({open_n63216,data_rd[34]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b0000101000001100),
    .MODE("LOGIC"))
    \_al_u8536|_al_u8689  (
    .a({uncache_data[50],uncache_data[50]}),
    .b({uncache_data[34],uncache_data[34]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u8536_o,_al_u8689_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(A*~(D*~(~C*~B)))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(A*~(D*~(~C*~B)))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b0000001010101010),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b0000001010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8538|_al_u8537  (
    .a({_al_u7995_o,uncache_data[58]}),
    .b({_al_u8536_o,uncache_data[42]}),
    .c({_al_u8537_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8538_o,_al_u8537_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b0000000011100100),
    .MODE("LOGIC"))
    \_al_u8540|_al_u8542  (
    .a({\exu/mux27_b32_sel_is_1_o ,open_n63261}),
    .b({data_rd[34],_al_u2855_o}),
    .c({data_rd[35],_al_u8541_o}),
    .d({shift_l,_al_u8540_o}),
    .f({_al_u8540_o,_al_u8542_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b1100101000000000),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b1100101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8541|_al_u8554  (
    .a({data_rd[33],open_n63282}),
    .b({data_rd[34],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[33]}),
    .d({shift_l,\exu/n59_lutinv }),
    .f({_al_u8541_o,_al_u8554_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8544|_al_u8543  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [34]}),
    .b({_al_u3712_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [34],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8544_o,\exu/alu_au/n31 [34]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b0101110111010000),
    .MODE("LOGIC"))
    \_al_u8546|_al_u3714  (
    .a({_al_u8545_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[34],ds1[34]}),
    .d({ds2[34],ds2[34]}),
    .f({_al_u8546_o,\exu/alu_au/n55 [34]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8548|_al_u8547  (
    .a({_al_u8544_o,and_clr}),
    .b({_al_u8546_o,rd_data_and}),
    .c({_al_u2855_o,ds1[34]}),
    .d({\exu/alu_au/n33 [34],ds2[34]}),
    .f({_al_u8548_o,\exu/alu_au/n33 [34]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*D))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~(B*D))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0011000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8550|_al_u8384  (
    .b({open_n63377,\exu/lsu/mux27_b56_sel_is_3_o }),
    .c({\exu/lsu/n2_lutinv ,\exu/n60_lutinv }),
    .d({_al_u8383_o,_al_u8383_o}),
    .f({_al_u8550_o,_al_u8384_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    //.LUT1("(C*~(D*~(~B*~A)))"),
    .INIT_LUT0(16'b1010001100000000),
    .INIT_LUT1(16'b0001000011110000),
    .MODE("LOGIC"))
    \_al_u8553|_al_u8551  (
    .a({_al_u8550_o,_al_u8093_o}),
    .b({_al_u8551_o,_al_u8232_o}),
    .c({_al_u8552_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8553_o,_al_u8551_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1011111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8555|exu/reg1_b33  (
    .a({_al_u8125_o,_al_u8555_o}),
    .b({_al_u8126_o,_al_u8559_o}),
    .c({_al_u8553_o,_al_u8565_o}),
    .clk(clk_pad),
    .d({_al_u8554_o,_al_u8568_o}),
    .sr(rst_pad),
    .f({_al_u8555_o,open_n63435}),
    .q({open_n63439,data_rd[33]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(A*~(D*~(C*B)))"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b1000000010101010),
    .MODE("LOGIC"))
    \_al_u8558|_al_u8557  (
    .a({_al_u7995_o,uncache_data[57]}),
    .b({_al_u8556_o,uncache_data[33]}),
    .c({_al_u8557_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8558_o,_al_u8557_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*A*~(D*~B))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*A*~(D*~B))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000100000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8561|_al_u8560  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [33]}),
    .b({_al_u3720_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [33],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8561_o,\exu/alu_au/n31 [33]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8563|_al_u8562  (
    .a({_al_u8562_o,open_n63484}),
    .b({rd_data_xor,rd_data_or}),
    .c({ds1[33],ds1[33]}),
    .d({ds2[33],rd_data_ds1}),
    .f({_al_u8563_o,_al_u8562_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8565|_al_u8564  (
    .a({_al_u8561_o,and_clr}),
    .b({_al_u8563_o,rd_data_and}),
    .c({_al_u2855_o,ds1[33]}),
    .d({\exu/alu_au/n33 [33],ds2[33]}),
    .f({_al_u8565_o,\exu/alu_au/n33 [33]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000110010001000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b0000110010001000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8566|_al_u8568  (
    .a({open_n63533,\exu/n57 [33]}),
    .b({data_rd[33],_al_u2855_o}),
    .c({data_rd[34],_al_u8567_o}),
    .d({\exu/mux27_b32_sel_is_1_o ,shift_l}),
    .f({\exu/n57 [33],_al_u8568_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8567|_al_u8574  (
    .b({data_rd[33],\exu/n60_lutinv }),
    .c({ex_size[2],data_rd[32]}),
    .d({data_rd[32],\exu/n59_lutinv }),
    .f({_al_u8567_o,_al_u8574_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8570|_al_u7936  (
    .b({open_n63586,_al_u3224_o}),
    .c({\exu/lsu/n0_lutinv ,uncache_data[32]}),
    .d({_al_u7936_o,\biu/l1d_out [32]}),
    .f({_al_u8570_o,_al_u7936_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u8572|_al_u8403  (
    .b({_al_u8127_o,\exu/lsu/mux27_b56_sel_is_3_o }),
    .c({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .d({_al_u8402_o,_al_u8402_o}),
    .f({_al_u8572_o,_al_u8403_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    //.LUT1("(C*~(D*~(~B*~A)))"),
    .INIT_LUT0(16'b0101110000000000),
    .INIT_LUT1(16'b0001000011110000),
    .MODE("LOGIC"))
    \_al_u8573|_al_u8571  (
    .a({_al_u8570_o,_al_u8109_o}),
    .b({_al_u8571_o,_al_u8249_o}),
    .c({_al_u8572_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8573_o,_al_u8571_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(C*B*~A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(C*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1011111100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1011111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8575|exu/reg1_b32  (
    .a({_al_u8125_o,_al_u8575_o}),
    .b({_al_u8126_o,_al_u8579_o}),
    .c({_al_u8573_o,_al_u8585_o}),
    .clk(clk_pad),
    .d({_al_u8574_o,_al_u8588_o}),
    .sr(rst_pad),
    .f({_al_u8575_o,open_n63670}),
    .q({open_n63674,data_rd[32]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(A*~(D*~(C*B)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(A*~(D*~(C*B)))"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b1000000010101010),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b1000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8578|_al_u8577  (
    .a({_al_u7995_o,uncache_data[56]}),
    .b({_al_u8576_o,uncache_data[32]}),
    .c({_al_u8577_o,addr_ex[0]}),
    .d({unsign,addr_ex[1]}),
    .f({_al_u8578_o,_al_u8577_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(~C*A*~(D*~B))"),
    .INIT_LUT0(16'b1100000010100000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"))
    \_al_u8581|_al_u8580  (
    .a({\exu/c_stb_lutinv ,\exu/alu_au/add_64 [32]}),
    .b({_al_u3728_o,\exu/alu_au/sub_64 [31]}),
    .c({\exu/alu_au/n31 [32],rd_data_sub}),
    .d({rd_data_add,ex_size[2]}),
    .f({_al_u8581_o,\exu/alu_au/n31 [32]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*D))"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG0("(~B*~(C*D))"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0101110111010000),
    .INIT_LUTG0(16'b0000001100110011),
    .INIT_LUTG1(16'b0101110111010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8583|_al_u8582  (
    .a({_al_u8582_o,open_n63719}),
    .b({rd_data_xor,rd_data_or}),
    .c({ds1[32],ds1[32]}),
    .d({ds2[32],rd_data_ds1}),
    .f({_al_u8583_o,_al_u8582_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~C*~(~D*~B*A))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0000111100001101),
    .MODE("LOGIC"))
    \_al_u8585|_al_u8584  (
    .a({_al_u8581_o,and_clr}),
    .b({_al_u8583_o,rd_data_and}),
    .c({_al_u2855_o,ds1[32]}),
    .d({\exu/alu_au/n33 [32],ds2[32]}),
    .f({_al_u8585_o,\exu/alu_au/n33 [32]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~C*~(~D*A)))"),
    //.LUTF1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUTG0("(B*~(~C*~(~D*A)))"),
    //.LUTG1("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT_LUTF0(16'b1100000011001000),
    .INIT_LUTF1(16'b1100101000000000),
    .INIT_LUTG0(16'b1100000011001000),
    .INIT_LUTG1(16'b1100101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8587|_al_u8588  (
    .a({data_rd[31],\exu/n57 [32]}),
    .b({data_rd[32],_al_u2855_o}),
    .c({ex_size[2],_al_u8587_o}),
    .d({shift_l,shift_l}),
    .f({_al_u8587_o,_al_u8588_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(~D*~(~C*~B))"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"))
    \_al_u8591|_al_u8966  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[31],data_rd[13]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8591_o,_al_u8966_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1111110100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8592|exu/reg1_b31  (
    .a({_al_u7905_o,_al_u8592_o}),
    .b({_al_u7973_o,_al_u8594_o}),
    .c({_al_u8590_o,_al_u8600_o}),
    .clk(clk_pad),
    .d({_al_u8591_o,_al_u8603_o}),
    .sr(rst_pad),
    .f({_al_u8592_o,open_n63823}),
    .q({open_n63827,data_rd[31]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8593|_al_u8594  (
    .b({_al_u7994_o,\exu/c_stb_lutinv }),
    .c({_al_u7912_o,\exu/n59_lutinv }),
    .d({_al_u7991_o,_al_u8593_o}),
    .f({_al_u8593_o,_al_u8594_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8597|_al_u8596  (
    .a({_al_u8595_o,\exu/alu_au/sub_64 [31]}),
    .b({_al_u8596_o,rd_data_ds1}),
    .c({\exu/alu_au/add_64 [31],rd_data_sub}),
    .d({rd_data_add,ds1[31]}),
    .f({_al_u8597_o,_al_u8596_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u8600|_al_u8599  (
    .a({open_n63878,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [31],ds1[31]}),
    .d({_al_u8598_o,ds2[31]}),
    .f({_al_u8600_o,\exu/alu_au/n33 [31]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~B*A))"),
    //.LUT1("(B*~(C*~(D*~A)))"),
    .INIT_LUT0(16'b0000110100001111),
    .INIT_LUT1(16'b0100110000001100),
    .MODE("LOGIC"))
    \_al_u8602|_al_u8601  (
    .a({\exu/lsu/n56 ,data_rd[32]}),
    .b({_al_u8601_o,ex_size[2]}),
    .c({data_rd[31],shift_l}),
    .d({shift_r,shift_r}),
    .f({_al_u8602_o,_al_u8601_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(~C*~(~B*~D))"),
    //.LUTG0("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(~C*~(~B*~D))"),
    .INIT_LUTF0(16'b0101001100000000),
    .INIT_LUTF1(16'b0000111100001100),
    .INIT_LUTG0(16'b0101001100000000),
    .INIT_LUTG1(16'b0000111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8608|_al_u8607  (
    .a({open_n63919,_al_u8146_o}),
    .b({_al_u8607_o,_al_u8286_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8606_o,addr_ex[1]}),
    .f({_al_u8608_o,_al_u8607_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A*~(D*~C))"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("(B*~A*~(D*~C))"),
    //.LUTG1("(~D*~(~C*~B))"),
    .INIT_LUTF0(16'b0100000001000100),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b0100000001000100),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8609|_al_u8603  (
    .a({open_n63944,_al_u8602_o}),
    .b({\exu/n60_lutinv ,_al_u2855_o}),
    .c({data_rd[30],data_rd[30]}),
    .d({\exu/n59_lutinv ,shift_l}),
    .f({_al_u8609_o,_al_u8603_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1111110100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8610|exu/reg1_b30  (
    .a({_al_u7905_o,_al_u8610_o}),
    .b({_al_u7973_o,_al_u8614_o}),
    .c({_al_u8608_o,_al_u8620_o}),
    .clk(clk_pad),
    .d({_al_u8609_o,_al_u8622_o}),
    .sr(rst_pad),
    .f({_al_u8610_o,open_n63982}),
    .q({open_n63986,data_rd[30]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(~C*~(B*D))"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"))
    \_al_u8613|_al_u8612  (
    .a({open_n63987,uncache_data[54]}),
    .b({_al_u8612_o,uncache_data[30]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8611_o,addr_ex[1]}),
    .f({_al_u8613_o,_al_u8612_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*A)))"),
    //.LUT1("(~C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000001000001111),
    .INIT_LUT1(16'b0000001000001111),
    .MODE("LOGIC"))
    \_al_u8614|_al_u8880  (
    .a({_al_u7991_o,_al_u7991_o}),
    .b({_al_u8613_o,_al_u8879_o}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8614_o,_al_u8880_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8617|_al_u8615  (
    .a({_al_u8615_o,\exu/c_stb_lutinv }),
    .b({_al_u8616_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [30],ds1[30]}),
    .d({rd_data_add,ds2[30]}),
    .f({_al_u8617_o,_al_u8615_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u8618|_al_u3743  (
    .a({_al_u8617_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[30],ds1[30]}),
    .d({ds2[30],ds2[30]}),
    .f({_al_u8618_o,\exu/alu_au/n55 [30]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u8620|_al_u8619  (
    .a({open_n64072,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [30],ds1[30]}),
    .d({_al_u8618_o,ds2[30]}),
    .f({_al_u8620_o,\exu/alu_au/n33 [30]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8621|_al_u8622  (
    .a({open_n64093,_al_u2855_o}),
    .b({data_rd[31],\exu/n57 [30]}),
    .c({shift_r,data_rd[29]}),
    .d({data_rd[30],shift_l}),
    .f({\exu/n57 [30],_al_u8622_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1100101000000000),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8624|_al_u8466  (
    .a({open_n64114,\biu/l1d_out [37]}),
    .b({uncache_data[37],uncache_data[37]}),
    .c({_al_u3224_o,_al_u3224_o}),
    .d({\biu/l1d_out [37],\exu/lsu/n0_lutinv }),
    .f({_al_u8624_o,_al_u8466_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b0000110000111111),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8625|_al_u8631  (
    .a({open_n64135,uncache_data[45]}),
    .b({_al_u3224_o,uncache_data[29]}),
    .c({uncache_data[29],addr_ex[0]}),
    .d({\biu/l1d_out [29],addr_ex[1]}),
    .f({_al_u8625_o,_al_u8631_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(~C*~(~B*~D))"),
    //.LUTG0("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(~C*~(~B*~D))"),
    .INIT_LUTF0(16'b0000000001010011),
    .INIT_LUTF1(16'b0000111100001100),
    .INIT_LUTG0(16'b0000000001010011),
    .INIT_LUTG1(16'b0000111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8628|_al_u8626  (
    .a({open_n64160,_al_u8624_o}),
    .b({_al_u8627_o,_al_u8625_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8626_o,addr_ex[1]}),
    .f({_al_u8628_o,_al_u8626_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(~D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8629|_al_u8929  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[29],data_rd[14]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8629_o,_al_u8929_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(~C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1111110100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1111110100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8630|exu/reg1_b29  (
    .a({_al_u7905_o,_al_u8630_o}),
    .b({_al_u7973_o,_al_u8634_o}),
    .c({_al_u8628_o,_al_u8640_o}),
    .clk(clk_pad),
    .d({_al_u8629_o,_al_u8642_o}),
    .sr(rst_pad),
    .f({_al_u8630_o,open_n64228}),
    .q({open_n64232,data_rd[29]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~C*~(~B*~D))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~C*~(~B*~D))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b0000111100001100),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b0000111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8633|_al_u8632  (
    .a({open_n64233,uncache_data[53]}),
    .b({_al_u8632_o,uncache_data[37]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8631_o,addr_ex[1]}),
    .f({_al_u8633_o,_al_u8632_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*A)))"),
    //.LUTF1("(~C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*A)))"),
    //.LUTG1("(~C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000001000001111),
    .INIT_LUTF1(16'b0000001000001111),
    .INIT_LUTG0(16'b0000001000001111),
    .INIT_LUTG1(16'b0000001000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8634|_al_u8862  (
    .a({_al_u7991_o,_al_u7991_o}),
    .b({_al_u8633_o,_al_u8861_o}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8634_o,_al_u8862_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u8637|_al_u8635  (
    .a({_al_u8635_o,\exu/c_stb_lutinv }),
    .b({_al_u8636_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [29],ds1[29]}),
    .d({rd_data_add,ds2[29]}),
    .f({_al_u8637_o,_al_u8635_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8638|_al_u3757  (
    .a({_al_u8637_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[29],ds1[29]}),
    .d({ds2[29],ds2[29]}),
    .f({_al_u8638_o,\exu/alu_au/n55 [29]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8640|_al_u8639  (
    .a({open_n64326,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [29],ds1[29]}),
    .d({_al_u8638_o,ds2[29]}),
    .f({_al_u8640_o,\exu/alu_au/n33 [29]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8641|_al_u8642  (
    .a({open_n64351,_al_u2855_o}),
    .b({data_rd[30],\exu/n57 [29]}),
    .c({shift_r,data_rd[28]}),
    .d({data_rd[29],shift_l}),
    .f({\exu/n57 [29],_al_u8642_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    //.LUT1("(~C*~(~B*D))"),
    .INIT_LUT0(16'b0101000011000000),
    .INIT_LUT1(16'b0000110000001111),
    .MODE("LOGIC"))
    \_al_u8644|_al_u8994  (
    .a({open_n64376,_al_u8644_o}),
    .b({_al_u3224_o,_al_u8798_o}),
    .c({_al_u8488_o,addr_ex[0]}),
    .d({\biu/l1d_out [36],addr_ex[1]}),
    .f({_al_u8644_o,_al_u8994_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b0000001111001111),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b0000001111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8645|_al_u8652  (
    .a({open_n64397,uncache_data[44]}),
    .b({_al_u3224_o,uncache_data[28]}),
    .c({\biu/l1d_out [28],addr_ex[0]}),
    .d({uncache_data[28],addr_ex[1]}),
    .f({_al_u8645_o,_al_u8652_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(~C*~(~B*~D))"),
    //.LUTG0("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(~C*~(~B*~D))"),
    .INIT_LUTF0(16'b0000000001010011),
    .INIT_LUTF1(16'b0000111100001100),
    .INIT_LUTG0(16'b0000000001010011),
    .INIT_LUTG1(16'b0000111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8648|_al_u8646  (
    .a({open_n64422,_al_u8644_o}),
    .b({_al_u8647_o,_al_u8645_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8646_o,addr_ex[1]}),
    .f({_al_u8648_o,_al_u8646_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(~D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8649|_al_u8891  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[28],data_rd[15]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8649_o,_al_u8891_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1111110100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8650|exu/reg1_b28  (
    .a({_al_u7905_o,_al_u8650_o}),
    .b({_al_u7973_o,_al_u8654_o}),
    .c({_al_u8648_o,_al_u8660_o}),
    .clk(clk_pad),
    .d({_al_u8649_o,_al_u8662_o}),
    .sr(rst_pad),
    .f({_al_u8650_o,open_n64486}),
    .q({open_n64490,data_rd[28]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8653|_al_u8651  (
    .a({open_n64491,uncache_data[52]}),
    .b({_al_u8652_o,uncache_data[36]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8651_o,addr_ex[1]}),
    .f({_al_u8653_o,_al_u8651_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*A)))"),
    //.LUTF1("(~C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*A)))"),
    //.LUTG1("(~C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000001000001111),
    .INIT_LUTF1(16'b0000001000001111),
    .INIT_LUTG0(16'b0000001000001111),
    .INIT_LUTG1(16'b0000001000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8654|_al_u8844  (
    .a({_al_u7991_o,_al_u7991_o}),
    .b({_al_u8653_o,_al_u8843_o}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8654_o,_al_u8844_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8657|_al_u8655  (
    .a({_al_u8655_o,\exu/c_stb_lutinv }),
    .b({_al_u8656_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [28],ds1[28]}),
    .d({rd_data_add,ds2[28]}),
    .f({_al_u8657_o,_al_u8655_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8658|_al_u3764  (
    .a({_al_u8657_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[28],ds1[28]}),
    .d({ds2[28],ds2[28]}),
    .f({_al_u8658_o,\exu/alu_au/n55 [28]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8660|_al_u8659  (
    .a({open_n64584,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [28],ds1[28]}),
    .d({_al_u8658_o,ds2[28]}),
    .f({_al_u8660_o,\exu/alu_au/n33 [28]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8661|_al_u8662  (
    .a({open_n64609,_al_u2855_o}),
    .b({data_rd[29],\exu/n57 [28]}),
    .c({shift_r,data_rd[27]}),
    .d({data_rd[28],shift_l}),
    .f({\exu/n57 [28],_al_u8662_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b0000010100000011),
    .INIT_LUTF1(16'b0000001111001111),
    .INIT_LUTG0(16'b0000010100000011),
    .INIT_LUTG1(16'b0000001111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8665|_al_u9029  (
    .a({open_n64630,_al_u8665_o}),
    .b({_al_u3224_o,_al_u9012_o}),
    .c({\biu/l1d_out [27],addr_ex[0]}),
    .d({uncache_data[27],addr_ex[1]}),
    .f({_al_u8665_o,_al_u9029_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(~C*~(B*D))"),
    .INIT_LUT0(16'b0101111111111100),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"))
    \_al_u8667|_al_u8666  (
    .a({open_n64655,_al_u8198_o}),
    .b({_al_u8666_o,_al_u8665_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8664_o,addr_ex[1]}),
    .f({_al_u8667_o,_al_u8666_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(~D*~(~C*~B))"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"))
    \_al_u8668|_al_u8875  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[27],data_rd[16]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8668_o,_al_u8875_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1111110100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8669|exu/reg1_b27  (
    .a({_al_u7905_o,_al_u8669_o}),
    .b({_al_u7973_o,_al_u8673_o}),
    .c({_al_u8667_o,_al_u8679_o}),
    .clk(clk_pad),
    .d({_al_u8668_o,_al_u8681_o}),
    .sr(rst_pad),
    .f({_al_u8669_o,open_n64711}),
    .q({open_n64715,data_rd[27]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~C*~(B*D))"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"))
    \_al_u8672|_al_u8671  (
    .a({open_n64716,uncache_data[43]}),
    .b({_al_u8671_o,uncache_data[35]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8670_o,addr_ex[1]}),
    .f({_al_u8672_o,_al_u8671_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*A)))"),
    //.LUT1("(~C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000001000001111),
    .INIT_LUT1(16'b0000001000001111),
    .MODE("LOGIC"))
    \_al_u8673|_al_u8825  (
    .a({_al_u7991_o,_al_u7991_o}),
    .b({_al_u8672_o,_al_u8824_o}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8673_o,_al_u8825_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u8676|_al_u8674  (
    .a({_al_u8674_o,\exu/c_stb_lutinv }),
    .b({_al_u8675_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [27],ds1[27]}),
    .d({rd_data_add,ds2[27]}),
    .f({_al_u8676_o,_al_u8674_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u8677|_al_u3771  (
    .a({_al_u8676_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[27],ds1[27]}),
    .d({ds2[27],ds2[27]}),
    .f({_al_u8677_o,\exu/alu_au/n55 [27]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u8679|_al_u8678  (
    .a({open_n64797,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [27],ds1[27]}),
    .d({_al_u8677_o,ds2[27]}),
    .f({_al_u8679_o,\exu/alu_au/n33 [27]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8680|_al_u8681  (
    .a({open_n64818,_al_u2855_o}),
    .b({data_rd[28],\exu/n57 [27]}),
    .c({shift_r,data_rd[26]}),
    .d({data_rd[27],shift_l}),
    .f({\exu/n57 [27],_al_u8681_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTF1("(~C*~(B*D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    //.LUTG1("(~C*~(B*D))"),
    .INIT_LUTF0(16'b1010111111110011),
    .INIT_LUTF1(16'b0000001100001111),
    .INIT_LUTG0(16'b1010111111110011),
    .INIT_LUTG1(16'b0000001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8686|_al_u8685  (
    .a({open_n64843,_al_u8215_o}),
    .b({_al_u8685_o,_al_u8684_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8683_o,addr_ex[1]}),
    .f({_al_u8686_o,_al_u8685_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(~D*~(~C*~B))"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"))
    \_al_u8687|_al_u8857  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[26],data_rd[17]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8687_o,_al_u8857_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(~C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1111110100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1111110100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8688|exu/reg1_b26  (
    .a({_al_u7905_o,_al_u8688_o}),
    .b({_al_u7973_o,_al_u8692_o}),
    .c({_al_u8686_o,_al_u8698_o}),
    .clk(clk_pad),
    .d({_al_u8687_o,_al_u8700_o}),
    .sr(rst_pad),
    .f({_al_u8688_o,open_n64907}),
    .q({open_n64911,data_rd[26]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~C*~(~B*~D))"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~C*~(~B*~D))"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b0000111100001100),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b0000111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8691|_al_u8690  (
    .a({open_n64912,uncache_data[42]}),
    .b({_al_u8690_o,uncache_data[26]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8689_o,addr_ex[1]}),
    .f({_al_u8691_o,_al_u8690_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*A)))"),
    //.LUT1("(~C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000001000001111),
    .INIT_LUT1(16'b0000001000001111),
    .MODE("LOGIC"))
    \_al_u8692|_al_u8806  (
    .a({_al_u7991_o,_al_u7991_o}),
    .b({_al_u8691_o,_al_u8805_o}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8692_o,_al_u8806_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8695|_al_u8693  (
    .a({_al_u8693_o,\exu/c_stb_lutinv }),
    .b({_al_u8694_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [26],ds1[26]}),
    .d({rd_data_add,ds2[26]}),
    .f({_al_u8695_o,_al_u8693_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u8696|_al_u3778  (
    .a({_al_u8695_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[26],ds1[26]}),
    .d({ds2[26],ds2[26]}),
    .f({_al_u8696_o,\exu/alu_au/n55 [26]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u8698|_al_u8697  (
    .a({open_n65001,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [26],ds1[26]}),
    .d({_al_u8696_o,ds2[26]}),
    .f({_al_u8698_o,\exu/alu_au/n33 [26]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8699|_al_u8700  (
    .a({open_n65022,_al_u2855_o}),
    .b({data_rd[27],\exu/n57 [26]}),
    .c({shift_r,data_rd[25]}),
    .d({data_rd[26],shift_l}),
    .f({\exu/n57 [26],_al_u8700_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~C*~(B*D))"),
    .INIT_LUT0(16'b1100111111111010),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"))
    \_al_u8704|_al_u8703  (
    .a({open_n65043,_al_u7907_o}),
    .b({_al_u8703_o,_al_u8232_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8702_o,addr_ex[1]}),
    .f({_al_u8704_o,_al_u8703_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(~D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8705|_al_u8839  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[25],data_rd[18]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8705_o,_al_u8839_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(~C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1111110100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1111110100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8706|exu/reg1_b25  (
    .a({_al_u7905_o,_al_u8706_o}),
    .b({_al_u7973_o,_al_u8710_o}),
    .c({_al_u8704_o,_al_u8716_o}),
    .clk(clk_pad),
    .d({_al_u8705_o,_al_u8718_o}),
    .sr(rst_pad),
    .f({_al_u8706_o,open_n65107}),
    .q({open_n65111,data_rd[25]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8709|_al_u8708  (
    .a({open_n65112,uncache_data[41]}),
    .b({_al_u8708_o,uncache_data[25]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8707_o,addr_ex[1]}),
    .f({_al_u8709_o,_al_u8708_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*A)))"),
    //.LUTF1("(~C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*A)))"),
    //.LUTG1("(~C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000001000001111),
    .INIT_LUTF1(16'b0000001000001111),
    .INIT_LUTG0(16'b0000001000001111),
    .INIT_LUTG1(16'b0000001000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8710|_al_u8787  (
    .a({_al_u7991_o,_al_u7991_o}),
    .b({_al_u8709_o,_al_u8786_o}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8710_o,_al_u8787_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u8713|_al_u8711  (
    .a({_al_u8711_o,\exu/c_stb_lutinv }),
    .b({_al_u8712_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [25],ds1[25]}),
    .d({rd_data_add,ds2[25]}),
    .f({_al_u8713_o,_al_u8711_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8714|_al_u3785  (
    .a({_al_u8713_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[25],ds1[25]}),
    .d({ds2[25],ds2[25]}),
    .f({_al_u8714_o,\exu/alu_au/n55 [25]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8716|_al_u8715  (
    .a({open_n65201,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [25],ds1[25]}),
    .d({_al_u8714_o,ds2[25]}),
    .f({_al_u8716_o,\exu/alu_au/n33 [25]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8717|_al_u8718  (
    .a({open_n65226,_al_u2855_o}),
    .b({data_rd[26],\exu/n57 [25]}),
    .c({shift_r,data_rd[24]}),
    .d({data_rd[25],shift_l}),
    .f({\exu/n57 [25],_al_u8718_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(~C*~(~B*~D))"),
    //.LUTG0("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(~C*~(~B*~D))"),
    .INIT_LUTF0(16'b1100000010100000),
    .INIT_LUTF1(16'b0000111100001100),
    .INIT_LUTG0(16'b1100000010100000),
    .INIT_LUTG1(16'b0000111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8722|_al_u8721  (
    .a({open_n65251,_al_u7936_o}),
    .b({_al_u8721_o,_al_u8249_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8720_o,addr_ex[1]}),
    .f({_al_u8722_o,_al_u8721_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(~D*~(~C*~B))"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8723|_al_u8820  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[24],data_rd[19]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8723_o,_al_u8820_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1111110100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8724|exu/reg1_b24  (
    .a({_al_u7905_o,_al_u8724_o}),
    .b({_al_u7973_o,_al_u8728_o}),
    .c({_al_u8722_o,_al_u8734_o}),
    .clk(clk_pad),
    .d({_al_u8723_o,_al_u8736_o}),
    .sr(rst_pad),
    .f({_al_u8724_o,open_n65315}),
    .q({open_n65319,data_rd[24]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~C*~(~B*~D))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~C*~(~B*~D))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b0000111100001100),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b0000111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8727|_al_u8726  (
    .a({open_n65320,uncache_data[48]}),
    .b({_al_u8726_o,uncache_data[32]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8725_o,addr_ex[1]}),
    .f({_al_u8727_o,_al_u8726_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*A)))"),
    //.LUTF1("(~C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*A)))"),
    //.LUTG1("(~C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000001000001111),
    .INIT_LUTF1(16'b0000001000001111),
    .INIT_LUTG0(16'b0000001000001111),
    .INIT_LUTG1(16'b0000001000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8728|_al_u8768  (
    .a({_al_u7991_o,_al_u7991_o}),
    .b({_al_u8727_o,_al_u8767_o}),
    .c({\exu/c_stb_lutinv ,\exu/c_stb_lutinv }),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8728_o,_al_u8768_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8731|_al_u8729  (
    .a({_al_u8729_o,\exu/c_stb_lutinv }),
    .b({_al_u8730_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [24],ds1[24]}),
    .d({rd_data_add,ds2[24]}),
    .f({_al_u8731_o,_al_u8729_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8732|_al_u3792  (
    .a({_al_u8731_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[24],ds1[24]}),
    .d({ds2[24],ds2[24]}),
    .f({_al_u8732_o,\exu/alu_au/n55 [24]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8734|_al_u8733  (
    .a({open_n65417,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [24],ds1[24]}),
    .d({_al_u8732_o,ds2[24]}),
    .f({_al_u8734_o,\exu/alu_au/n33 [24]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8735|_al_u8736  (
    .a({open_n65442,_al_u2855_o}),
    .b({data_rd[25],\exu/n57 [24]}),
    .c({shift_r,data_rd[23]}),
    .d({data_rd[24],shift_l}),
    .f({\exu/n57 [24],_al_u8736_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000001010011),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000000001010011),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8738|_al_u8740  (
    .a({open_n65463,_al_u8738_o}),
    .b({uncache_data[31],_al_u8739_o}),
    .c({_al_u3224_o,addr_ex[0]}),
    .d({\biu/l1d_out [31],addr_ex[1]}),
    .f({_al_u8738_o,_al_u8740_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1100101000000000),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u8741|_al_u7977  (
    .a({open_n65488,\biu/l1d_out [39]}),
    .b({uncache_data[39],uncache_data[39]}),
    .c({_al_u3224_o,_al_u3224_o}),
    .d({\biu/l1d_out [39],\exu/lsu/n2_lutinv }),
    .f({_al_u8741_o,_al_u7977_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b0011010100000000),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8743|_al_u8742  (
    .a({open_n65509,_al_u8741_o}),
    .b({_al_u8742_o,_al_u8267_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8740_o,addr_ex[1]}),
    .f({_al_u8743_o,_al_u8742_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(~D*~(~C*~B))"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"))
    \_al_u8744|_al_u8801  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c({data_rd[23],data_rd[20]}),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8744_o,_al_u8801_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1111110100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8745|exu/reg1_b23  (
    .a({_al_u7905_o,_al_u8745_o}),
    .b({_al_u7973_o,_al_u8749_o}),
    .c({_al_u8743_o,_al_u8755_o}),
    .clk(clk_pad),
    .d({_al_u8744_o,_al_u8757_o}),
    .sr(rst_pad),
    .f({_al_u8745_o,open_n65565}),
    .q({open_n65569,data_rd[23]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8748|_al_u8746  (
    .a({open_n65570,uncache_data[39]}),
    .b({_al_u8747_o,uncache_data[23]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8746_o,addr_ex[1]}),
    .f({_al_u8748_o,_al_u8746_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u8752|_al_u8750  (
    .a({_al_u8750_o,\exu/c_stb_lutinv }),
    .b({_al_u8751_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [23],ds1[23]}),
    .d({rd_data_add,ds2[23]}),
    .f({_al_u8752_o,_al_u8750_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u8753|_al_u3799  (
    .a({_al_u8752_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[23],ds1[23]}),
    .d({ds2[23],ds2[23]}),
    .f({_al_u8753_o,\exu/alu_au/n55 [23]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u8755|_al_u8754  (
    .a({open_n65631,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [23],ds1[23]}),
    .d({_al_u8753_o,ds2[23]}),
    .f({_al_u8755_o,\exu/alu_au/n33 [23]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8756|_al_u8757  (
    .a({open_n65652,_al_u2855_o}),
    .b({data_rd[24],\exu/n57 [23]}),
    .c({shift_r,data_rd[22]}),
    .d({data_rd[23],shift_l}),
    .f({\exu/n57 [23],_al_u8757_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b0000001111001111),
    .MODE("LOGIC"))
    \_al_u8759|_al_u8765  (
    .a({open_n65677,uncache_data[46]}),
    .b({_al_u3224_o,uncache_data[22]}),
    .c({\biu/l1d_out [22],addr_ex[0]}),
    .d({uncache_data[22],addr_ex[1]}),
    .f({_al_u8759_o,_al_u8765_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b0101110000000000),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8762|_al_u8761  (
    .a({open_n65698,_al_u8286_o}),
    .b({_al_u8761_o,_al_u8444_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8760_o,addr_ex[1]}),
    .f({_al_u8762_o,_al_u8761_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(~D*~(~C*~B))"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"))
    \_al_u8763|_al_u8782  (
    .b({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .c(data_rd[22:21]),
    .d({\exu/n59_lutinv ,\exu/n59_lutinv }),
    .f({_al_u8763_o,_al_u8782_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(~C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1111110100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1111110100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8764|exu/reg1_b22  (
    .a({_al_u7905_o,_al_u8764_o}),
    .b({_al_u7973_o,_al_u8768_o}),
    .c({_al_u8762_o,_al_u8774_o}),
    .clk(clk_pad),
    .d({_al_u8763_o,_al_u8776_o}),
    .sr(rst_pad),
    .f({_al_u8764_o,open_n65758}),
    .q({open_n65762,data_rd[22]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~C*~(B*D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~C*~(B*D))"),
    .INIT_LUTF0(16'b1111010100111111),
    .INIT_LUTF1(16'b0000001100001111),
    .INIT_LUTG0(16'b1111010100111111),
    .INIT_LUTG1(16'b0000001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8767|_al_u8766  (
    .a({open_n65763,uncache_data[38]}),
    .b({_al_u8766_o,uncache_data[30]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8765_o,addr_ex[1]}),
    .f({_al_u8767_o,_al_u8766_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8771|_al_u8769  (
    .a({_al_u8769_o,\exu/c_stb_lutinv }),
    .b({_al_u8770_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [22],ds1[22]}),
    .d({rd_data_add,ds2[22]}),
    .f({_al_u8771_o,_al_u8769_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u8774|_al_u8773  (
    .a({open_n65812,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [22],ds1[22]}),
    .d({_al_u8772_o,ds2[22]}),
    .f({_al_u8774_o,\exu/alu_au/n33 [22]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8775|_al_u8776  (
    .a({open_n65833,_al_u2855_o}),
    .b({data_rd[23],\exu/n57 [22]}),
    .c({shift_r,data_rd[21]}),
    .d({data_rd[22],shift_l}),
    .f({\exu/n57 [22],_al_u8776_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b1111001111000000),
    .MODE("LOGIC"))
    \_al_u8779|_al_u8784  (
    .a({open_n65854,uncache_data[37]}),
    .b({_al_u3224_o,uncache_data[21]}),
    .c({uncache_data[21],addr_ex[0]}),
    .d({\biu/l1d_out [21],addr_ex[1]}),
    .f({_al_u8779_o,_al_u8784_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~C*~(B*D))"),
    .INIT_LUT0(16'b1111101011001111),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"))
    \_al_u8781|_al_u8778  (
    .a({open_n65875,_al_u8624_o}),
    .b({_al_u8780_o,_al_u8625_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8778_o,addr_ex[1]}),
    .f({_al_u8781_o,_al_u8778_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(~C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1111110100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1111110100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8783|exu/reg1_b21  (
    .a({_al_u7905_o,_al_u8783_o}),
    .b({_al_u7973_o,_al_u8787_o}),
    .c({_al_u8781_o,_al_u8793_o}),
    .clk(clk_pad),
    .d({_al_u8782_o,_al_u8795_o}),
    .sr(rst_pad),
    .f({_al_u8783_o,open_n65913}),
    .q({open_n65917,data_rd[21]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8786|_al_u8785  (
    .a({open_n65918,uncache_data[45]}),
    .b({_al_u8785_o,uncache_data[29]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8784_o,addr_ex[1]}),
    .f({_al_u8786_o,_al_u8785_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u8790|_al_u8788  (
    .a({_al_u8788_o,\exu/c_stb_lutinv }),
    .b({_al_u8789_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [21],ds1[21]}),
    .d({rd_data_add,ds2[21]}),
    .f({_al_u8790_o,_al_u8788_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u8791|_al_u3813  (
    .a({_al_u8790_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[21],ds1[21]}),
    .d({ds2[21],ds2[21]}),
    .f({_al_u8791_o,\exu/alu_au/n55 [21]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8793|_al_u8792  (
    .a({open_n65979,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [21],ds1[21]}),
    .d({_al_u8791_o,ds2[21]}),
    .f({_al_u8793_o,\exu/alu_au/n33 [21]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8794|_al_u8795  (
    .a({open_n66004,_al_u2855_o}),
    .b({data_rd[22],\exu/n57 [21]}),
    .c({shift_r,data_rd[20]}),
    .d({data_rd[21],shift_l}),
    .f({\exu/n57 [21],_al_u8795_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8798|_al_u8804  (
    .a({open_n66029,uncache_data[36]}),
    .b({_al_u3224_o,uncache_data[20]}),
    .c({\biu/l1d_out [20],addr_ex[0]}),
    .d({uncache_data[20],addr_ex[1]}),
    .f({_al_u8798_o,_al_u8804_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~C*~(B*D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~C*~(B*D))"),
    .INIT_LUTF0(16'b1111101011001111),
    .INIT_LUTF1(16'b0000001100001111),
    .INIT_LUTG0(16'b1111101011001111),
    .INIT_LUTG1(16'b0000001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8800|_al_u8797  (
    .a({open_n66054,_al_u8644_o}),
    .b({_al_u8799_o,_al_u8645_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8797_o,addr_ex[1]}),
    .f({_al_u8800_o,_al_u8797_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1111110100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8802|exu/reg1_b20  (
    .a({_al_u7905_o,_al_u8802_o}),
    .b({_al_u7973_o,_al_u8806_o}),
    .c({_al_u8800_o,_al_u8812_o}),
    .clk(clk_pad),
    .d({_al_u8801_o,_al_u8814_o}),
    .sr(rst_pad),
    .f({_al_u8802_o,open_n66092}),
    .q({open_n66096,data_rd[20]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8805|_al_u8803  (
    .a({open_n66097,uncache_data[44]}),
    .b({_al_u8804_o,uncache_data[28]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8803_o,addr_ex[1]}),
    .f({_al_u8805_o,_al_u8803_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8809|_al_u8807  (
    .a({_al_u8807_o,\exu/c_stb_lutinv }),
    .b({_al_u8808_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [20],ds1[20]}),
    .d({rd_data_add,ds2[20]}),
    .f({_al_u8809_o,_al_u8807_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8810|_al_u3820  (
    .a({_al_u8809_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[20],ds1[20]}),
    .d({ds2[20],ds2[20]}),
    .f({_al_u8810_o,\exu/alu_au/n55 [20]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8812|_al_u8811  (
    .a({open_n66166,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [20],ds1[20]}),
    .d({_al_u8810_o,ds2[20]}),
    .f({_al_u8812_o,\exu/alu_au/n33 [20]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8813|_al_u8814  (
    .a({open_n66191,_al_u2855_o}),
    .b({data_rd[21],\exu/n57 [20]}),
    .c({shift_r,data_rd[19]}),
    .d({data_rd[20],shift_l}),
    .f({\exu/n57 [20],_al_u8814_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b0000001111001111),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b0000001111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8816|_al_u8823  (
    .a({open_n66212,uncache_data[43]}),
    .b({_al_u3224_o,uncache_data[19]}),
    .c({\biu/l1d_out [19],addr_ex[0]}),
    .d({uncache_data[19],addr_ex[1]}),
    .f({_al_u8816_o,_al_u8823_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b0101001100000000),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8819|_al_u8818  (
    .a({open_n66237,_al_u8345_o}),
    .b({_al_u8818_o,_al_u8508_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8817_o,addr_ex[1]}),
    .f({_al_u8819_o,_al_u8818_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(~C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1111110100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1111110100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8821|exu/reg1_b19  (
    .a({_al_u7905_o,_al_u8821_o}),
    .b({_al_u7973_o,_al_u8825_o}),
    .c({_al_u8819_o,_al_u8831_o}),
    .clk(clk_pad),
    .d({_al_u8820_o,_al_u8833_o}),
    .sr(rst_pad),
    .f({_al_u8821_o,open_n66275}),
    .q({open_n66279,data_rd[19]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~C*~(B*D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~C*~(B*D))"),
    .INIT_LUTF0(16'b1111010100111111),
    .INIT_LUTF1(16'b0000001100001111),
    .INIT_LUTG0(16'b1111010100111111),
    .INIT_LUTG1(16'b0000001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8824|_al_u8822  (
    .a({open_n66280,uncache_data[35]}),
    .b({_al_u8823_o,uncache_data[27]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8822_o,addr_ex[1]}),
    .f({_al_u8824_o,_al_u8822_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u8828|_al_u8826  (
    .a({_al_u8826_o,\exu/c_stb_lutinv }),
    .b({_al_u8827_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [19],ds1[19]}),
    .d({rd_data_add,ds2[19]}),
    .f({_al_u8828_o,_al_u8826_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u8829|_al_u3834  (
    .a({_al_u8828_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[19],ds1[19]}),
    .d({ds2[19],ds2[19]}),
    .f({_al_u8829_o,\exu/alu_au/n55 [19]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u8831|_al_u8830  (
    .a({open_n66345,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [19],ds1[19]}),
    .d({_al_u8829_o,ds2[19]}),
    .f({_al_u8831_o,\exu/alu_au/n33 [19]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8832|_al_u8833  (
    .a({open_n66366,_al_u2855_o}),
    .b({data_rd[20],\exu/n57 [19]}),
    .c({shift_r,data_rd[18]}),
    .d({data_rd[19],shift_l}),
    .f({\exu/n57 [19],_al_u8833_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b1111001111000000),
    .MODE("LOGIC"))
    \_al_u8835|_al_u8842  (
    .a({open_n66391,uncache_data[34]}),
    .b({_al_u3224_o,uncache_data[18]}),
    .c({uncache_data[18],addr_ex[0]}),
    .d({\biu/l1d_out [18],addr_ex[1]}),
    .f({_al_u8835_o,_al_u8842_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    //.LUTF1("(~C*~(~B*~D))"),
    //.LUTG0("(D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    //.LUTG1("(~C*~(~B*~D))"),
    .INIT_LUTF0(16'b0101110000000000),
    .INIT_LUTF1(16'b0000111100001100),
    .INIT_LUTG0(16'b0101110000000000),
    .INIT_LUTG1(16'b0000111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8838|_al_u8837  (
    .a({open_n66412,_al_u8364_o}),
    .b({_al_u8837_o,_al_u8531_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8836_o,addr_ex[1]}),
    .f({_al_u8838_o,_al_u8837_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(~C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1111110100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1111110100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8840|exu/reg1_b18  (
    .a({_al_u7905_o,_al_u8840_o}),
    .b({_al_u7973_o,_al_u8844_o}),
    .c({_al_u8838_o,_al_u8850_o}),
    .clk(clk_pad),
    .d({_al_u8839_o,_al_u8852_o}),
    .sr(rst_pad),
    .f({_al_u8840_o,open_n66454}),
    .q({open_n66458,data_rd[18]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~C*~(~B*~D))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~C*~(~B*~D))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b0000111100001100),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b0000111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8843|_al_u8841  (
    .a({open_n66459,uncache_data[42]}),
    .b({_al_u8842_o,uncache_data[26]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8841_o,addr_ex[1]}),
    .f({_al_u8843_o,_al_u8841_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8847|_al_u8845  (
    .a({_al_u8845_o,\exu/c_stb_lutinv }),
    .b({_al_u8846_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [18],ds1[18]}),
    .d({rd_data_add,ds2[18]}),
    .f({_al_u8847_o,_al_u8845_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u8848|_al_u3841  (
    .a({_al_u8847_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[18],ds1[18]}),
    .d({ds2[18],ds2[18]}),
    .f({_al_u8848_o,\exu/alu_au/n55 [18]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u8850|_al_u8849  (
    .a({open_n66528,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [18],ds1[18]}),
    .d({_al_u8848_o,ds2[18]}),
    .f({_al_u8850_o,\exu/alu_au/n33 [18]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8851|_al_u8852  (
    .a({open_n66549,_al_u2855_o}),
    .b({data_rd[19],\exu/n57 [18]}),
    .c({shift_r,data_rd[17]}),
    .d({data_rd[18],shift_l}),
    .f({\exu/n57 [18],_al_u8852_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~C*~(B*D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~C*~(B*D))"),
    .INIT_LUTF0(16'b1111101011001111),
    .INIT_LUTF1(16'b0000001100001111),
    .INIT_LUTG0(16'b1111101011001111),
    .INIT_LUTG1(16'b0000001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8856|_al_u8854  (
    .a({open_n66570,_al_u7906_o}),
    .b({_al_u8855_o,_al_u7907_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8854_o,addr_ex[1]}),
    .f({_al_u8856_o,_al_u8854_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1111110100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8858|exu/reg1_b17  (
    .a({_al_u7905_o,_al_u8858_o}),
    .b({_al_u7973_o,_al_u8862_o}),
    .c({_al_u8856_o,_al_u8868_o}),
    .clk(clk_pad),
    .d({_al_u8857_o,_al_u8870_o}),
    .sr(rst_pad),
    .f({_al_u8858_o,open_n66608}),
    .q({open_n66612,data_rd[17]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~C*~(B*D))"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b0000001100001111),
    .MODE("LOGIC"))
    \_al_u8861|_al_u8860  (
    .a({open_n66613,uncache_data[33]}),
    .b({_al_u8860_o,uncache_data[25]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8859_o,addr_ex[1]}),
    .f({_al_u8861_o,_al_u8860_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u8865|_al_u8863  (
    .a({_al_u8863_o,\exu/c_stb_lutinv }),
    .b({_al_u8864_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [17],ds1[17]}),
    .d({rd_data_add,ds2[17]}),
    .f({_al_u8865_o,_al_u8863_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8866|_al_u3848  (
    .a({_al_u8865_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[17],ds1[17]}),
    .d({ds2[17],ds2[17]}),
    .f({_al_u8866_o,\exu/alu_au/n55 [17]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8868|_al_u8867  (
    .a({open_n66678,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [17],ds1[17]}),
    .d({_al_u8866_o,ds2[17]}),
    .f({_al_u8868_o,\exu/alu_au/n33 [17]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8869|_al_u8870  (
    .a({open_n66703,_al_u2855_o}),
    .b({data_rd[18],\exu/n57 [17]}),
    .c({shift_r,data_rd[16]}),
    .d({data_rd[17],shift_l}),
    .f({\exu/n57 [17],_al_u8870_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b0011101000000000),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8874|_al_u8872  (
    .a({open_n66728,_al_u7936_o}),
    .b({_al_u8873_o,_al_u8402_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8872_o,addr_ex[1]}),
    .f({_al_u8874_o,_al_u8872_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b1111110100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8876|exu/reg1_b16  (
    .a({_al_u7905_o,_al_u8876_o}),
    .b({_al_u7973_o,_al_u8880_o}),
    .c({_al_u8874_o,_al_u8886_o}),
    .clk(clk_pad),
    .d({_al_u8875_o,_al_u8888_o}),
    .sr(rst_pad),
    .f({_al_u8876_o,open_n66762}),
    .q({open_n66766,data_rd[16]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~C*~(~B*~D))"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b0000111100001100),
    .MODE("LOGIC"))
    \_al_u8879|_al_u8878  (
    .a({open_n66767,uncache_data[40]}),
    .b({_al_u8878_o,uncache_data[24]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({_al_u8877_o,addr_ex[1]}),
    .f({_al_u8879_o,_al_u8878_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8883|_al_u8881  (
    .a({_al_u8881_o,\exu/c_stb_lutinv }),
    .b({_al_u8882_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [16],ds1[16]}),
    .d({rd_data_add,ds2[16]}),
    .f({_al_u8883_o,_al_u8881_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8884|_al_u3855  (
    .a({_al_u8883_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[16],ds1[16]}),
    .d({ds2[16],ds2[16]}),
    .f({_al_u8884_o,\exu/alu_au/n55 [16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8886|_al_u8885  (
    .a({open_n66836,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [16],ds1[16]}),
    .d({_al_u8884_o,ds2[16]}),
    .f({_al_u8886_o,\exu/alu_au/n33 [16]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8887|_al_u8888  (
    .a({open_n66861,_al_u2855_o}),
    .b({data_rd[17],\exu/n57 [16]}),
    .c({shift_r,data_rd[15]}),
    .d({data_rd[16],shift_l}),
    .f({\exu/n57 [16],_al_u8888_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(D*~(~C*~B*A))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(D*~(~C*~B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b1111110100000000),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b1111110100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8892|exu/reg1_b15  (
    .a({_al_u7905_o,_al_u8892_o}),
    .b({_al_u7973_o,_al_u8894_o}),
    .c({_al_u8890_o,_al_u8900_o}),
    .clk(clk_pad),
    .d({_al_u8891_o,_al_u8902_o}),
    .sr(rst_pad),
    .f({_al_u8892_o,open_n66899}),
    .q({open_n66903,data_rd[15]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(D*~(~C*~B))"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(D*~(~C*~B))"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8893|_al_u8894  (
    .b({_al_u7990_o,\exu/c_stb_lutinv }),
    .c({_al_u7912_o,\exu/n59_lutinv }),
    .d({_al_u7991_o,_al_u8893_o}),
    .f({_al_u8893_o,_al_u8894_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u8897|_al_u8895  (
    .a({_al_u8895_o,\exu/c_stb_lutinv }),
    .b({_al_u8896_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [15],ds1[15]}),
    .d({rd_data_add,ds2[15]}),
    .f({_al_u8897_o,_al_u8895_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u8898|_al_u3862  (
    .a({_al_u8897_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[15],ds1[15]}),
    .d({ds2[15],ds2[15]}),
    .f({_al_u8898_o,\exu/alu_au/n55 [15]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u8900|_al_u8899  (
    .a({open_n66970,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [15],ds1[15]}),
    .d({_al_u8898_o,ds2[15]}),
    .f({_al_u8900_o,\exu/alu_au/n33 [15]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8901|_al_u8902  (
    .a({open_n66991,_al_u2855_o}),
    .b({data_rd[16],\exu/n57 [15]}),
    .c({shift_r,data_rd[14]}),
    .d({data_rd[15],shift_l}),
    .f({\exu/n57 [15],_al_u8902_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8905|_al_u8925  (
    .a({open_n67016,uncache_data[38]}),
    .b({_al_u3224_o,uncache_data[14]}),
    .c({\biu/l1d_out [14],addr_ex[0]}),
    .d({uncache_data[14],addr_ex[1]}),
    .f({_al_u8905_o,_al_u8925_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b0000000010100011),
    .INIT_LUT1(16'b1111101000111111),
    .MODE("LOGIC"))
    \_al_u8906|_al_u8760  (
    .a({_al_u8759_o,_al_u8605_o}),
    .b({_al_u8905_o,_al_u8759_o}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u8906_o,_al_u8760_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(B*~A*~(D*C))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"))
    \_al_u8907|_al_u8923  (
    .a({_al_u8904_o,_al_u8605_o}),
    .b({_al_u8906_o,_al_u8905_o}),
    .c({_al_u8605_o,addr_ex[0]}),
    .d({\exu/lsu/n8_lutinv ,addr_ex[1]}),
    .f({_al_u8907_o,_al_u8923_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u8908|_al_u9052  (
    .c({data_rd[6],data_rd[2]}),
    .d({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .f({_al_u8908_o,_al_u9052_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(~D*~(~C*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b0000000011110100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8909|exu/reg1_b6  (
    .a({_al_u8907_o,_al_u8909_o}),
    .b({_al_u7953_o,_al_u8912_o}),
    .c({_al_u8908_o,_al_u8918_o}),
    .clk(clk_pad),
    .d({\exu/n59_lutinv ,_al_u8920_o}),
    .sr(rst_pad),
    .f({_al_u8909_o,open_n67118}),
    .q({open_n67122,data_rd[6]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~D*~(C*~(B*A)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~D*~(C*~(B*A)))"),
    .INIT_LUTF0(16'b1111010100111111),
    .INIT_LUTF1(16'b0000000010001111),
    .INIT_LUTG0(16'b1111010100111111),
    .INIT_LUTG1(16'b0000000010001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8912|_al_u8911  (
    .a({_al_u8910_o,uncache_data[22]}),
    .b({_al_u8911_o,uncache_data[14]}),
    .c({_al_u7956_o,addr_ex[0]}),
    .d({\exu/c_stb_lutinv ,addr_ex[1]}),
    .f({_al_u8912_o,_al_u8911_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8915|_al_u8913  (
    .a({_al_u8913_o,\exu/c_stb_lutinv }),
    .b({_al_u8914_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [6],ds1[6]}),
    .d({rd_data_add,ds2[6]}),
    .f({_al_u8915_o,_al_u8913_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u8916|_al_u3491  (
    .a({_al_u8915_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[6],ds1[6]}),
    .d({ds2[6],ds2[6]}),
    .f({_al_u8916_o,\exu/alu_au/n55 [6]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u8918|_al_u8917  (
    .a({open_n67191,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [6],ds1[6]}),
    .d({_al_u8916_o,ds2[6]}),
    .f({_al_u8918_o,\exu/alu_au/n33 [6]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8919|_al_u8920  (
    .a({open_n67212,_al_u2855_o}),
    .b({data_rd[7],\exu/n57 [6]}),
    .c({shift_r,data_rd[5]}),
    .d({data_rd[6],shift_l}),
    .f({\exu/n57 [6],_al_u8920_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    //.LUTF1("(~(~D*C)*~(~B*~A))"),
    //.LUTG0("(C*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    //.LUTG1("(~(~D*C)*~(~B*~A))"),
    .INIT_LUTF0(16'b1010000000110000),
    .INIT_LUTF1(16'b1110111000001110),
    .INIT_LUTG0(16'b1010000000110000),
    .INIT_LUTG1(16'b1110111000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8924|_al_u8922  (
    .a({_al_u8922_o,_al_u8444_o}),
    .b({_al_u8923_o,_al_u8759_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u8924_o,_al_u8922_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(~D*C)*~(B*A))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(~D*C)*~(B*A))"),
    .INIT_LUTF0(16'b1111010100111111),
    .INIT_LUTF1(16'b0111011100000111),
    .INIT_LUTG0(16'b1111010100111111),
    .INIT_LUTG1(16'b0111011100000111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8927|_al_u8926  (
    .a({_al_u8925_o,uncache_data[30]}),
    .b({_al_u8926_o,uncache_data[22]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u8927_o,_al_u8926_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*~A)))"),
    //.LUT1("(C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000000100001111),
    .INIT_LUT1(16'b0010000011110000),
    .MODE("LOGIC"))
    \_al_u8930|_al_u8928  (
    .a({_al_u7905_o,\exu/lsu/n52 [10]}),
    .b({_al_u8924_o,_al_u8927_o}),
    .c({_al_u8928_o,\exu/c_stb_lutinv }),
    .d({_al_u8929_o,\exu/n59_lutinv }),
    .f({_al_u8930_o,_al_u8928_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u8933|_al_u8931  (
    .a({_al_u8931_o,\exu/c_stb_lutinv }),
    .b({_al_u8932_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [14],ds1[14]}),
    .d({rd_data_add,ds2[14]}),
    .f({_al_u8933_o,_al_u8931_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(B*~D))"),
    //.LUT1("(~B*~(A*~(D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111100),
    .INIT_LUT1(16'b0011000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8935|exu/reg1_b14  (
    .a({_al_u8934_o,open_n67321}),
    .b({_al_u2855_o,_al_u8935_o}),
    .c({\exu/alu_au/alu_and [14],_al_u8937_o}),
    .clk(clk_pad),
    .d({rd_data_and,_al_u8930_o}),
    .sr(rst_pad),
    .f({_al_u8935_o,open_n67335}),
    .q({open_n67339,data_rd[14]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8936|_al_u8937  (
    .a({open_n67340,_al_u2855_o}),
    .b({data_rd[15],\exu/n57 [14]}),
    .c({shift_r,data_rd[13]}),
    .d({data_rd[14],shift_l}),
    .f({\exu/n57 [14],_al_u8937_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000110000111111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u8939|_al_u8942  (
    .b({open_n67363,_al_u3224_o}),
    .c({\biu/l1d_out [5],uncache_data[13]}),
    .d({_al_u3224_o,\biu/l1d_out [13]}),
    .f({_al_u8939_o,_al_u8942_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(~(C*~B)*~(D*~A))"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b1000101011001111),
    .MODE("LOGIC"))
    \_al_u8941|_al_u8940  (
    .a({_al_u8625_o,open_n67384}),
    .b({_al_u8939_o,_al_u3224_o}),
    .c({_al_u8940_o,\exu/lsu/n0_lutinv }),
    .d({\exu/lsu/n8_lutinv ,uncache_data[5]}),
    .f({_al_u8941_o,_al_u8940_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000010100000011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000010100000011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8943|_al_u8959  (
    .a({open_n67405,_al_u8625_o}),
    .b({open_n67406,_al_u8942_o}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[0]}),
    .d({_al_u8942_o,addr_ex[1]}),
    .f({_al_u8943_o,_al_u8959_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u8945|_al_u9015  (
    .c({data_rd[5],data_rd[3]}),
    .d({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .f({_al_u8945_o,_al_u9015_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(~D*~(~C*~(B*~A)))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(~D*~(~C*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b0000000011110100),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b0000000011110100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8946|exu/reg1_b5  (
    .a({_al_u8944_o,_al_u8946_o}),
    .b({_al_u7953_o,_al_u8949_o}),
    .c({_al_u8945_o,_al_u8955_o}),
    .clk(clk_pad),
    .d({\exu/n59_lutinv ,_al_u8957_o}),
    .sr(rst_pad),
    .f({_al_u8946_o,open_n67472}),
    .q({open_n67476,data_rd[5]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b0000110000001010),
    .MODE("LOGIC"))
    \_al_u8947|_al_u8962  (
    .a({uncache_data[5],uncache_data[29]}),
    .b({uncache_data[21],uncache_data[21]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u8947_o,_al_u8962_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~D*~(C*~(~B*~A)))"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b0000000000011111),
    .MODE("LOGIC"))
    \_al_u8949|_al_u8948  (
    .a({_al_u8947_o,uncache_data[29]}),
    .b({_al_u8948_o,uncache_data[13]}),
    .c({_al_u7956_o,addr_ex[0]}),
    .d({\exu/c_stb_lutinv ,addr_ex[1]}),
    .f({_al_u8949_o,_al_u8948_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8952|_al_u8950  (
    .a({_al_u8950_o,\exu/c_stb_lutinv }),
    .b({_al_u8951_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [5],ds1[5]}),
    .d({rd_data_add,ds2[5]}),
    .f({_al_u8952_o,_al_u8950_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8953|_al_u3578  (
    .a({_al_u8952_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[5],ds1[5]}),
    .d({ds2[5],ds2[5]}),
    .f({_al_u8953_o,\exu/alu_au/n55 [5]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8955|_al_u8954  (
    .a({open_n67565,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [5],ds1[5]}),
    .d({_al_u8953_o,ds2[5]}),
    .f({_al_u8955_o,\exu/alu_au/n33 [5]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8956|_al_u8957  (
    .a({open_n67590,_al_u2855_o}),
    .b({data_rd[6],\exu/n57 [5]}),
    .c({shift_r,data_rd[4]}),
    .d({data_rd[5],shift_l}),
    .f({\exu/n57 [5],_al_u8957_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    //.LUTF1("(~(~D*C)*~(~B*~A))"),
    //.LUTG0("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    //.LUTG1("(~(~D*C)*~(~B*~A))"),
    .INIT_LUTF0(16'b0101000011000000),
    .INIT_LUTF1(16'b1110111000001110),
    .INIT_LUTG0(16'b0101000011000000),
    .INIT_LUTG1(16'b1110111000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8961|_al_u8960  (
    .a({_al_u8959_o,_al_u8624_o}),
    .b({_al_u8960_o,_al_u8779_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u8961_o,_al_u8960_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(~(~D*C)*~(B*A))"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b0111011100000111),
    .MODE("LOGIC"))
    \_al_u8964|_al_u8963  (
    .a({_al_u8962_o,uncache_data[37]}),
    .b({_al_u8963_o,uncache_data[13]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u8964_o,_al_u8963_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*~A)))"),
    //.LUT1("(C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000000100001111),
    .INIT_LUT1(16'b0010000011110000),
    .MODE("LOGIC"))
    \_al_u8967|_al_u8965  (
    .a({_al_u7905_o,\exu/lsu/n52 [10]}),
    .b({_al_u8961_o,_al_u8964_o}),
    .c({_al_u8965_o,\exu/c_stb_lutinv }),
    .d({_al_u8966_o,\exu/n59_lutinv }),
    .f({_al_u8967_o,_al_u8965_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8970|_al_u8968  (
    .a({_al_u8968_o,\exu/c_stb_lutinv }),
    .b({_al_u8969_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [13],ds1[13]}),
    .d({rd_data_add,ds2[13]}),
    .f({_al_u8970_o,_al_u8968_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(B*~D))"),
    //.LUT1("(~B*~(A*~(D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111100),
    .INIT_LUT1(16'b0011000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8972|exu/reg1_b13  (
    .a({_al_u8971_o,open_n67703}),
    .b({_al_u2855_o,_al_u8972_o}),
    .c({\exu/alu_au/alu_and [13],_al_u8974_o}),
    .clk(clk_pad),
    .d({rd_data_and,_al_u8967_o}),
    .sr(rst_pad),
    .f({_al_u8972_o,open_n67717}),
    .q({open_n67721,data_rd[13]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u8973|_al_u8974  (
    .a({open_n67722,_al_u2855_o}),
    .b({data_rd[14],\exu/n57 [13]}),
    .c({shift_r,data_rd[12]}),
    .d({data_rd[13],shift_l}),
    .f({\exu/n57 [13],_al_u8974_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u8977|_al_u8998  (
    .a({open_n67743,uncache_data[28]}),
    .b({_al_u3224_o,uncache_data[12]}),
    .c({\biu/l1d_out [12],addr_ex[0]}),
    .d({uncache_data[12],addr_ex[1]}),
    .f({_al_u8977_o,_al_u8998_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b1111010100111111),
    .MODE("LOGIC"))
    \_al_u8978|_al_u8982  (
    .a({_al_u8798_o,uncache_data[20]}),
    .b({_al_u8977_o,uncache_data[12]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u8978_o,_al_u8982_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUT1("(B*~A*~(D*~C))"),
    .INIT_LUT0(16'b1011000010000000),
    .INIT_LUT1(16'b0100000001000100),
    .MODE("LOGIC"))
    \_al_u8979|_al_u8976  (
    .a({_al_u8976_o,uncache_data[4]}),
    .b({_al_u8978_o,_al_u3224_o}),
    .c({_al_u8645_o,\exu/lsu/n0_lutinv }),
    .d({\exu/lsu/n8_lutinv ,\biu/l1d_out [4]}),
    .f({_al_u8979_o,_al_u8976_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(~D*~(~C*~(B*~A)))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(~D*~(~C*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b0000000011110100),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b0000000011110100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u8981|exu/reg1_b4  (
    .a({_al_u8979_o,_al_u8981_o}),
    .b({_al_u7953_o,_al_u8984_o}),
    .c({_al_u8980_o,_al_u8990_o}),
    .clk(clk_pad),
    .d({\exu/n59_lutinv ,_al_u8992_o}),
    .sr(rst_pad),
    .f({_al_u8981_o,open_n67821}),
    .q({open_n67825,data_rd[4]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUT1("(~D*~(C*~(B*A)))"),
    .INIT_LUT0(16'b0011111111110101),
    .INIT_LUT1(16'b0000000010001111),
    .MODE("LOGIC"))
    \_al_u8984|_al_u8983  (
    .a({_al_u8982_o,uncache_data[4]}),
    .b({_al_u8983_o,uncache_data[28]}),
    .c({_al_u7956_o,addr_ex[0]}),
    .d({\exu/c_stb_lutinv ,addr_ex[1]}),
    .f({_al_u8984_o,_al_u8983_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u8987|_al_u8985  (
    .a({_al_u8985_o,\exu/c_stb_lutinv }),
    .b({_al_u8986_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [4],ds1[4]}),
    .d({rd_data_add,ds2[4]}),
    .f({_al_u8987_o,_al_u8985_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8988|_al_u3665  (
    .a({_al_u8987_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[4],ds1[4]}),
    .d({ds2[4],ds2[4]}),
    .f({_al_u8988_o,\exu/alu_au/n55 [4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8990|_al_u8989  (
    .a({open_n67890,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [4],ds1[4]}),
    .d({_al_u8988_o,ds2[4]}),
    .f({_al_u8990_o,\exu/alu_au/n33 [4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8991|_al_u8992  (
    .a({open_n67915,_al_u2855_o}),
    .b({data_rd[5],\exu/n57 [4]}),
    .c({shift_r,data_rd[3]}),
    .d({data_rd[4],shift_l}),
    .f({\exu/n57 [4],_al_u8992_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    //.LUT1("(~(~D*C)*~(~B*~A))"),
    .INIT_LUT0(16'b0000010100001100),
    .INIT_LUT1(16'b1110111000001110),
    .MODE("LOGIC"))
    \_al_u8996|_al_u8995  (
    .a({_al_u8994_o,_al_u8645_o}),
    .b({_al_u8995_o,_al_u8977_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u8996_o,_al_u8995_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~(~D*C)*~(~B*~A))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~(~D*C)*~(~B*~A))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b1110111000001110),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b1110111000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u8999|_al_u8997  (
    .a({_al_u8997_o,uncache_data[36]}),
    .b({_al_u8998_o,uncache_data[20]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u8999_o,_al_u8997_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*~A)))"),
    //.LUTF1("(C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*~A)))"),
    //.LUTG1("(C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000000100001111),
    .INIT_LUTF1(16'b0010000011110000),
    .INIT_LUTG0(16'b0000000100001111),
    .INIT_LUTG1(16'b0010000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9002|_al_u9000  (
    .a({_al_u7905_o,\exu/lsu/n52 [10]}),
    .b({_al_u8996_o,_al_u8999_o}),
    .c({_al_u9000_o,\exu/c_stb_lutinv }),
    .d({_al_u9001_o,\exu/n59_lutinv }),
    .f({_al_u9002_o,_al_u9000_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u9005|_al_u9003  (
    .a({_al_u9003_o,\exu/c_stb_lutinv }),
    .b({_al_u9004_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [12],ds1[12]}),
    .d({rd_data_add,ds2[12]}),
    .f({_al_u9005_o,_al_u9003_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(B*~D))"),
    //.LUTF1("(~B*~(A*~(D*C)))"),
    //.LUTG0("~(~C*~(B*~D))"),
    //.LUTG1("(~B*~(A*~(D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111100),
    .INIT_LUTF1(16'b0011000100010001),
    .INIT_LUTG0(16'b1111000011111100),
    .INIT_LUTG1(16'b0011000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9007|exu/reg1_b12  (
    .a({_al_u9006_o,open_n68028}),
    .b({_al_u2855_o,_al_u9007_o}),
    .c({\exu/alu_au/alu_and [12],_al_u9009_o}),
    .clk(clk_pad),
    .d({rd_data_and,_al_u9002_o}),
    .sr(rst_pad),
    .f({_al_u9007_o,open_n68046}),
    .q({open_n68050,data_rd[12]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9008|_al_u9009  (
    .a({open_n68051,_al_u2855_o}),
    .b({data_rd[13],\exu/n57 [12]}),
    .c({shift_r,data_rd[11]}),
    .d({data_rd[12],shift_l}),
    .f({\exu/n57 [12],_al_u9009_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b0000001111001111),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b0000001111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9012|_al_u9032  (
    .a({open_n68076,uncache_data[27]}),
    .b({_al_u3224_o,uncache_data[11]}),
    .c({\biu/l1d_out [11],addr_ex[0]}),
    .d({uncache_data[11],addr_ex[1]}),
    .f({_al_u9012_o,_al_u9032_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b1111010100111111),
    .INIT_LUTF1(16'b1111101011001111),
    .INIT_LUTG0(16'b1111010100111111),
    .INIT_LUTG1(16'b1111101011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9013|_al_u9017  (
    .a({_al_u8816_o,uncache_data[19]}),
    .b({_al_u9012_o,uncache_data[11]}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u9013_o,_al_u9017_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(B*~A*~(D*~C))"),
    //.LUTG0("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(B*~A*~(D*~C))"),
    .INIT_LUTF0(16'b0000000001010011),
    .INIT_LUTF1(16'b0100000001000100),
    .INIT_LUTG0(16'b0000000001010011),
    .INIT_LUTG1(16'b0100000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9014|_al_u8817  (
    .a({_al_u9011_o,_al_u8665_o}),
    .b({_al_u9013_o,_al_u8816_o}),
    .c({_al_u8665_o,addr_ex[0]}),
    .d({\exu/lsu/n8_lutinv ,addr_ex[1]}),
    .f({_al_u9014_o,_al_u8817_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(~D*~(~C*~(B*~A)))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(~D*~(~C*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b0000000011110100),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b0000000011110100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9016|exu/reg1_b3  (
    .a({_al_u9014_o,_al_u9016_o}),
    .b({_al_u7953_o,_al_u9019_o}),
    .c({_al_u9015_o,_al_u9025_o}),
    .clk(clk_pad),
    .d({\exu/n59_lutinv ,_al_u9027_o}),
    .sr(rst_pad),
    .f({_al_u9016_o,open_n68166}),
    .q({open_n68170,data_rd[3]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTF1("(~D*~(C*~(B*A)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    //.LUTG1("(~D*~(C*~(B*A)))"),
    .INIT_LUTF0(16'b0011111111110101),
    .INIT_LUTF1(16'b0000000010001111),
    .INIT_LUTG0(16'b0011111111110101),
    .INIT_LUTG1(16'b0000000010001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9019|_al_u9018  (
    .a({_al_u9017_o,uncache_data[3]}),
    .b({_al_u9018_o,uncache_data[27]}),
    .c({_al_u7956_o,addr_ex[0]}),
    .d({\exu/c_stb_lutinv ,addr_ex[1]}),
    .f({_al_u9019_o,_al_u9018_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u9022|_al_u9020  (
    .a({_al_u9020_o,\exu/c_stb_lutinv }),
    .b({_al_u9021_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [3],ds1[3]}),
    .d({rd_data_add,ds2[3]}),
    .f({_al_u9022_o,_al_u9020_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u9023|_al_u3750  (
    .a({_al_u9022_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[3],ds1[3]}),
    .d({ds2[3],ds2[3]}),
    .f({_al_u9023_o,\exu/alu_au/n55 [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u9025|_al_u9024  (
    .a({open_n68235,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [3],ds1[3]}),
    .d({_al_u9023_o,ds2[3]}),
    .f({_al_u9025_o,\exu/alu_au/n33 [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u9026|_al_u9027  (
    .a({open_n68256,_al_u2855_o}),
    .b({data_rd[4],\exu/n57 [3]}),
    .c({shift_r,data_rd[2]}),
    .d({data_rd[3],shift_l}),
    .f({\exu/n57 [3],_al_u9027_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~(~D*C)*~(~B*~A))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b1110111000001110),
    .MODE("LOGIC"))
    \_al_u9031|_al_u9030  (
    .a({_al_u9029_o,_al_u8508_o}),
    .b({_al_u9030_o,_al_u8816_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u9031_o,_al_u9030_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~(~D*C)*~(~B*~A))"),
    //.LUTG0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~(~D*C)*~(~B*~A))"),
    .INIT_LUTF0(16'b1010000011000000),
    .INIT_LUTF1(16'b1110111000001110),
    .INIT_LUTG0(16'b1010000011000000),
    .INIT_LUTG1(16'b1110111000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9034|_al_u9033  (
    .a({_al_u9032_o,uncache_data[35]}),
    .b({_al_u9033_o,uncache_data[19]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u9034_o,_al_u9033_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D*~(~B*~A)))"),
    //.LUTF1("(C*~(D*~(~B*A)))"),
    //.LUTG0("(~C*~(D*~(~B*~A)))"),
    //.LUTG1("(C*~(D*~(~B*A)))"),
    .INIT_LUTF0(16'b0000000100001111),
    .INIT_LUTF1(16'b0010000011110000),
    .INIT_LUTG0(16'b0000000100001111),
    .INIT_LUTG1(16'b0010000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9037|_al_u9035  (
    .a({_al_u7905_o,\exu/lsu/n52 [10]}),
    .b({_al_u9031_o,_al_u9034_o}),
    .c({_al_u9035_o,\exu/c_stb_lutinv }),
    .d({_al_u9036_o,\exu/n59_lutinv }),
    .f({_al_u9037_o,_al_u9035_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9040|_al_u9038  (
    .a({_al_u9038_o,\exu/c_stb_lutinv }),
    .b({_al_u9039_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [11],ds1[11]}),
    .d({rd_data_add,ds2[11]}),
    .f({_al_u9040_o,_al_u9038_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(B*~D))"),
    //.LUTF1("(~B*~(A*~(D*C)))"),
    //.LUTG0("~(~C*~(B*~D))"),
    //.LUTG1("(~B*~(A*~(D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111100),
    .INIT_LUTF1(16'b0011000100010001),
    .INIT_LUTG0(16'b1111000011111100),
    .INIT_LUTG1(16'b0011000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9042|exu/reg1_b11  (
    .a({_al_u9041_o,open_n68369}),
    .b({_al_u2855_o,_al_u9042_o}),
    .c({\exu/alu_au/alu_and [11],_al_u9044_o}),
    .clk(clk_pad),
    .d({rd_data_and,_al_u9037_o}),
    .sr(rst_pad),
    .f({_al_u9042_o,open_n68387}),
    .q({open_n68391,data_rd[11]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1010000010001000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1010000010001000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9043|_al_u9044  (
    .a({open_n68392,_al_u2855_o}),
    .b({data_rd[12],\exu/n57 [11]}),
    .c({shift_r,data_rd[10]}),
    .d({data_rd[11],shift_l}),
    .f({\exu/n57 [11],_al_u9044_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUT1("(C*~(B*~D))"),
    .INIT_LUT0(16'b0101111111110011),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"))
    \_al_u9047|_al_u9054  (
    .a({open_n68417,uncache_data[26]}),
    .b({_al_u3224_o,uncache_data[2]}),
    .c({\exu/lsu/n0_lutinv ,addr_ex[0]}),
    .d({uncache_data[2],addr_ex[1]}),
    .f({_al_u9047_o,_al_u9054_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(~(C*~B)*~(D*A))"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b0100010111001111),
    .MODE("LOGIC"))
    \_al_u9048|_al_u8684  (
    .a({_al_u8684_o,open_n68438}),
    .b({_al_u9046_o,_al_u3224_o}),
    .c({_al_u9047_o,\biu/l1d_out [26]}),
    .d({\exu/lsu/n8_lutinv ,uncache_data[26]}),
    .f({_al_u9048_o,_al_u8684_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9049|_al_u9070  (
    .a({open_n68459,uncache_data[26]}),
    .b({_al_u3224_o,uncache_data[10]}),
    .c({uncache_data[10],addr_ex[0]}),
    .d({\biu/l1d_out [10],addr_ex[1]}),
    .f({_al_u9049_o,_al_u9070_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000010101100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u9050|_al_u9067  (
    .a({open_n68484,_al_u8835_o}),
    .b({open_n68485,_al_u9049_o}),
    .c({\exu/lsu/n2_lutinv ,addr_ex[0]}),
    .d({_al_u9049_o,addr_ex[1]}),
    .f({_al_u9050_o,_al_u9067_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUT1("(~B*A*~(D*C))"),
    .INIT_LUT0(16'b0000000010101100),
    .INIT_LUT1(16'b0000001000100010),
    .MODE("LOGIC"))
    \_al_u9051|_al_u8836  (
    .a({_al_u9048_o,_al_u8684_o}),
    .b({_al_u9050_o,_al_u8835_o}),
    .c({_al_u8835_o,addr_ex[0]}),
    .d({\exu/lsu/n5_lutinv ,addr_ex[1]}),
    .f({_al_u9051_o,_al_u8836_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(~D*~(~C*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b0000000011110100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9053|exu/reg1_b2  (
    .a({_al_u9051_o,_al_u9053_o}),
    .b({_al_u7953_o,_al_u9056_o}),
    .c({_al_u9052_o,_al_u9062_o}),
    .clk(clk_pad),
    .d({\exu/n59_lutinv ,_al_u9064_o}),
    .sr(rst_pad),
    .f({_al_u9053_o,open_n68539}),
    .q({open_n68543,data_rd[2]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~D*~(C*~(B*A)))"),
    .INIT_LUT0(16'b1111010100111111),
    .INIT_LUT1(16'b0000000010001111),
    .MODE("LOGIC"))
    \_al_u9056|_al_u9055  (
    .a({_al_u9054_o,uncache_data[18]}),
    .b({_al_u9055_o,uncache_data[10]}),
    .c({_al_u7956_o,addr_ex[0]}),
    .d({\exu/c_stb_lutinv ,addr_ex[1]}),
    .f({_al_u9056_o,_al_u9055_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9059|_al_u9057  (
    .a({_al_u9057_o,\exu/c_stb_lutinv }),
    .b({_al_u9058_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [2],ds1[2]}),
    .d({rd_data_add,ds2[2]}),
    .f({_al_u9059_o,_al_u9057_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(A*~(B*(D@C)))"),
    //.LUTG0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(A*~(B*(D@C)))"),
    .INIT_LUTF0(16'b1100010010000000),
    .INIT_LUTF1(16'b1010001000101010),
    .INIT_LUTG0(16'b1100010010000000),
    .INIT_LUTG1(16'b1010001000101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9060|_al_u3827  (
    .a({_al_u9059_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[2],ds1[2]}),
    .d({ds2[2],ds2[2]}),
    .f({_al_u9060_o,\exu/alu_au/n55 [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*(D@A))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0100000010000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u9062|_al_u9061  (
    .a({open_n68612,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [2],ds1[2]}),
    .d({_al_u9060_o,ds2[2]}),
    .f({_al_u9062_o,\exu/alu_au/n33 [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u9063|_al_u9064  (
    .a({open_n68633,_al_u2855_o}),
    .b({data_rd[3],\exu/n57 [2]}),
    .c({shift_r,data_rd[1]}),
    .d({data_rd[2],shift_l}),
    .f({\exu/n57 [2],_al_u9064_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUT1("(~(~D*C)*~(~B*~A))"),
    .INIT_LUT0(16'b1010110000000000),
    .INIT_LUT1(16'b1110111000001110),
    .MODE("LOGIC"))
    \_al_u9068|_al_u9066  (
    .a({_al_u9066_o,_al_u8531_o}),
    .b({_al_u9067_o,_al_u8684_o}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u9068_o,_al_u9066_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(~(~D*C)*~(~B*~A))"),
    .INIT_LUT0(16'b1010000011000000),
    .INIT_LUT1(16'b1110111000001110),
    .MODE("LOGIC"))
    \_al_u9071|_al_u9069  (
    .a({_al_u9069_o,uncache_data[34]}),
    .b({_al_u9070_o,uncache_data[18]}),
    .c({_al_u7912_o,addr_ex[0]}),
    .d({ex_size[1],addr_ex[1]}),
    .f({_al_u9071_o,_al_u9069_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~(~B*~A)))"),
    //.LUT1("(C*~(D*~(~B*A)))"),
    .INIT_LUT0(16'b0000000100001111),
    .INIT_LUT1(16'b0010000011110000),
    .MODE("LOGIC"))
    \_al_u9074|_al_u9072  (
    .a({_al_u7905_o,\exu/lsu/n52 [10]}),
    .b({_al_u9068_o,_al_u9071_o}),
    .c({_al_u9072_o,\exu/c_stb_lutinv }),
    .d({_al_u9073_o,\exu/n59_lutinv }),
    .f({_al_u9074_o,_al_u9072_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B*~(~D*~C)))"),
    //.LUT1("(B*A*~(D*C))"),
    .INIT_LUT0(16'b0010001000101010),
    .INIT_LUT1(16'b0000100010001000),
    .MODE("LOGIC"))
    \_al_u9077|_al_u9075  (
    .a({_al_u9075_o,\exu/c_stb_lutinv }),
    .b({_al_u9076_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [10],ds1[10]}),
    .d({rd_data_add,ds2[10]}),
    .f({_al_u9077_o,_al_u9075_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(B*~D))"),
    //.LUT1("(~B*~(A*~(D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111100),
    .INIT_LUT1(16'b0011000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9079|exu/reg1_b10  (
    .a({_al_u9078_o,open_n68734}),
    .b({_al_u2855_o,_al_u9079_o}),
    .c({\exu/alu_au/alu_and [10],_al_u9081_o}),
    .clk(clk_pad),
    .d({rd_data_and,_al_u9074_o}),
    .sr(rst_pad),
    .f({_al_u9079_o,open_n68748}),
    .q({open_n68752,data_rd[10]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u9080|_al_u9081  (
    .a({open_n68753,_al_u2855_o}),
    .b({data_rd[11],\exu/n57 [10]}),
    .c({shift_r,data_rd[9]}),
    .d({data_rd[10],shift_l}),
    .f({\exu/n57 [10],_al_u9081_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTF1("(C*~(B*~D))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    //.LUTG1("(C*~(B*~D))"),
    .INIT_LUTF0(16'b0101111111110011),
    .INIT_LUTF1(16'b1111000000110000),
    .INIT_LUTG0(16'b0101111111110011),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9084|_al_u9090  (
    .a({open_n68774,uncache_data[25]}),
    .b({_al_u3224_o,uncache_data[1]}),
    .c({\exu/lsu/n0_lutinv ,addr_ex[0]}),
    .d({uncache_data[1],addr_ex[1]}),
    .f({_al_u9084_o,_al_u9090_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~(C*~B)*~(D*~A))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1000101011001111),
    .MODE("LOGIC"))
    \_al_u9085|_al_u9083  (
    .a({_al_u7907_o,open_n68799}),
    .b({_al_u9083_o,open_n68800}),
    .c({_al_u9084_o,\biu/l1d_out [1]}),
    .d({\exu/lsu/n8_lutinv ,_al_u3224_o}),
    .f({_al_u9085_o,_al_u9083_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~B*A*~(D*C))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000001000100010),
    .MODE("LOGIC"))
    \_al_u9087|_al_u9086  (
    .a({_al_u9085_o,open_n68821}),
    .b({_al_u9086_o,open_n68822}),
    .c({_al_u7910_o,\exu/lsu/n2_lutinv }),
    .d({\exu/lsu/n5_lutinv ,_al_u7909_o}),
    .f({_al_u9087_o,_al_u9086_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(B*~A)))"),
    //.LUTF1("(~D*~(~C*~(B*~A)))"),
    //.LUTG0("~(~D*~(C*~(B*~A)))"),
    //.LUTG1("(~D*~(~C*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110110000),
    .INIT_LUTF1(16'b0000000011110100),
    .INIT_LUTG0(16'b1111111110110000),
    .INIT_LUTG1(16'b0000000011110100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9089|exu/reg1_b1  (
    .a({_al_u9087_o,_al_u9089_o}),
    .b({_al_u7953_o,_al_u9092_o}),
    .c({_al_u9088_o,_al_u9098_o}),
    .clk(clk_pad),
    .d({\exu/n59_lutinv ,_al_u9100_o}),
    .sr(rst_pad),
    .f({_al_u9089_o,open_n68860}),
    .q({open_n68864,data_rd[1]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~D*~(C*~(B*A)))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~D*~(C*~(B*A)))"),
    .INIT_LUTF0(16'b1111001101011111),
    .INIT_LUTF1(16'b0000000010001111),
    .INIT_LUTG0(16'b1111001101011111),
    .INIT_LUTG1(16'b0000000010001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9092|_al_u9091  (
    .a({_al_u9090_o,uncache_data[9]}),
    .b({_al_u9091_o,uncache_data[17]}),
    .c({_al_u7956_o,addr_ex[0]}),
    .d({\exu/c_stb_lutinv ,addr_ex[1]}),
    .f({_al_u9092_o,_al_u9091_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9095|_al_u9093  (
    .a({_al_u9093_o,\exu/c_stb_lutinv }),
    .b({_al_u9094_o,rd_data_or}),
    .c({\exu/alu_au/add_64 [1],ds1[1]}),
    .d({rd_data_add,ds2[1]}),
    .f({_al_u9095_o,_al_u9093_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(A*~(B*(D@C)))"),
    .INIT_LUT0(16'b1100010010000000),
    .INIT_LUT1(16'b1010001000101010),
    .MODE("LOGIC"))
    \_al_u9096|_al_u3909  (
    .a({_al_u9095_o,\exu/alu_au/ds1_light_than_ds2_lutinv }),
    .b({rd_data_xor,mem_csr_data_min}),
    .c({ds1[1],ds1[1]}),
    .d({ds2[1],ds2[1]}),
    .f({_al_u9096_o,\exu/alu_au/n55 [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9098|_al_u9097  (
    .a({open_n68933,and_clr}),
    .b({_al_u2855_o,rd_data_and}),
    .c({\exu/alu_au/n33 [1],ds1[1]}),
    .d({_al_u9096_o,ds2[1]}),
    .f({_al_u9098_o,\exu/alu_au/n33 [1]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u9099|_al_u9100  (
    .a({open_n68958,_al_u2855_o}),
    .b({data_rd[2],\exu/n57 [1]}),
    .c({shift_r,data_rd[0]}),
    .d({data_rd[1],shift_l}),
    .f({\exu/n57 [1],_al_u9100_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUTF0(16'b0000000010101100),
    .INIT_LUTF1(16'b1111010111001111),
    .INIT_LUTG0(16'b0000000010101100),
    .INIT_LUTG1(16'b1111010111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9103|_al_u8873  (
    .a({_al_u7933_o,_al_u7932_o}),
    .b({_al_u7935_o,_al_u7933_o}),
    .c({addr_ex[0],addr_ex[0]}),
    .d({addr_ex[1],addr_ex[1]}),
    .f({_al_u9103_o,_al_u8873_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTF1("(B*~A*~(D*C))"),
    //.LUTG0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG1("(B*~A*~(D*C))"),
    .INIT_LUTF0(16'b1011000010000000),
    .INIT_LUTF1(16'b0000010001000100),
    .INIT_LUTG0(16'b1011000010000000),
    .INIT_LUTG1(16'b0000010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9104|_al_u9102  (
    .a({_al_u9102_o,uncache_data[0]}),
    .b({_al_u9103_o,_al_u3224_o}),
    .c({_al_u7932_o,\exu/lsu/n0_lutinv }),
    .d({\exu/lsu/n8_lutinv ,\biu/l1d_out [0]}),
    .f({_al_u9104_o,_al_u9102_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9105|_al_u8980  (
    .c({data_rd[0],data_rd[4]}),
    .d({\exu/n60_lutinv ,\exu/n60_lutinv }),
    .f({_al_u9105_o,_al_u8980_o}));
  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(~D*~(~C*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b0000000011110100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9106|exu/reg1_b0  (
    .a({_al_u9104_o,_al_u9106_o}),
    .b({_al_u7953_o,_al_u9110_o}),
    .c({_al_u9105_o,_al_u9117_o}),
    .clk(clk_pad),
    .d({\exu/n59_lutinv ,_al_u9119_o}),
    .sr(rst_pad),
    .f({_al_u9106_o,open_n69068}),
    .q({open_n69072,data_rd[0]}));  // ../../RTL/CPU/EX/exu.v(327)
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(D*~(C*B))"),
    .INIT_LUT0(16'b1111001101011111),
    .INIT_LUT1(16'b0011111100000000),
    .MODE("LOGIC"))
    \_al_u9108|_al_u9107  (
    .a({open_n69073,uncache_data[8]}),
    .b({uncache_data[24],uncache_data[16]}),
    .c({\exu/lsu/n8_lutinv ,addr_ex[0]}),
    .d({_al_u9107_o,addr_ex[1]}),
    .f({_al_u9108_o,_al_u9107_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~(~B*A)))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000101111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u9109|_al_u9110  (
    .a({open_n69094,_al_u9108_o}),
    .b({open_n69095,\exu/lsu/n22 [0]}),
    .c({\exu/lsu/n0_lutinv ,_al_u7956_o}),
    .d({uncache_data[0],\exu/c_stb_lutinv }),
    .f({\exu/lsu/n22 [0],_al_u9110_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(B*~(~D*~C)))"),
    //.LUTF1("(B*A*~(D*C))"),
    //.LUTG0("(A*~(B*~(~D*~C)))"),
    //.LUTG1("(B*A*~(D*C))"),
    .INIT_LUTF0(16'b0010001000101010),
    .INIT_LUTF1(16'b0000100010001000),
    .INIT_LUTG0(16'b0010001000101010),
    .INIT_LUTG1(16'b0000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9113|_al_u9111  (
    .a({_al_u9111_o,\exu/c_stb_lutinv }),
    .b({_al_u9112_o,rd_data_or}),
    .c({\exu/alu_au/sub_64 [0],ds1[0]}),
    .d({rd_data_sub,ds2[0]}),
    .f({_al_u9113_o,_al_u9111_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*(D@A))"),
    //.LUTF1("(~C*~(~D*~B*A))"),
    //.LUTG0("(C*B*(D@A))"),
    //.LUTG1("(~C*~(~D*~B*A))"),
    .INIT_LUTF0(16'b0100000010000000),
    .INIT_LUTF1(16'b0000111100001101),
    .INIT_LUTG0(16'b0100000010000000),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9117|_al_u9116  (
    .a({_al_u9114_o,and_clr}),
    .b({\exu/alu_au/n39 [0],rd_data_and}),
    .c({_al_u2855_o,ds1[0]}),
    .d({\exu/alu_au/n33 [0],ds2[0]}),
    .f({_al_u9117_o,\exu/alu_au/n33 [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u9118|_al_u9119  (
    .b({data_rd[1],_al_u9118_o}),
    .c({shift_r,shift_l}),
    .d({data_rd[0],_al_u2855_o}),
    .f({_al_u9118_o,_al_u9119_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9121|_al_u3418  (
    .c({cache_reset,store}),
    .d({cache_flush,_al_u3181_o}),
    .f({_al_u9121_o,\exu/store_addr_mis }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~D)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(C*B*~D)"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0000000011000000),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000000011000000),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9122|_al_u2854  (
    .b({_al_u9121_o,\exu/c_stb_lutinv }),
    .c({amo,ex_valid}),
    .d({_al_u2852_o,_al_u2852_o}),
    .f({_al_u9122_o,\exu/n49 }));
  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*~(C*B*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111100000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0111111100000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9124|exu/valid_reg  (
    .a({open_n69240,_al_u9149_o}),
    .b({\exu/n17_lutinv ,ex_more_exception_neg_lutinv}),
    .c({ex_valid,\exu/n17_lutinv }),
    .clk(clk_pad),
    .d({\exu/c_stb_lutinv ,ex_valid}),
    .sr(\exu/n86 ),
    .f({\exu/n19 ,open_n69258}),
    .q({open_n69262,wb_valid}));  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(268)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(~C*B))"),
    //.LUT1("(~C*B*~(~D*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100001100),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9125|exu/reg8_b2  (
    .a({_al_u9122_o,open_n69263}),
    .b({\exu/n19 ,\exu/main_state [2]}),
    .c({load,_al_u9131_o}),
    .ce(ex_nop),
    .clk(clk_pad),
    .d({store,_al_u9125_o}),
    .sr(rst_pad),
    .f({_al_u9125_o,open_n69276}),
    .q({open_n69280,\exu/main_state [2]}));  // ../../RTL/CPU/EX/exu.v(268)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*~D)"),
    //.LUT1("(~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000011000000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"))
    \_al_u9126|_al_u9707  (
    .a({_al_u6309_o,open_n69281}),
    .b({_al_u6320_o,_al_u4399_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [7],\biu/cache_ctrl_logic/l1i_pte [7]}),
    .d({\biu/cache_ctrl_logic/l1d_pte [7],\biu/cache_ctrl_logic/n100 [4]}),
    .f({_al_u9126_o,_al_u9707_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~(~A*~(~D*B)))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~(~A*~(~D*B)))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000101000001110),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000101000001110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9127|_al_u2849  (
    .a({\biu/cache_ctrl_logic/n100 [4],open_n69302}),
    .b({_al_u3222_o,open_n69303}),
    .c({_al_u2848_o,rst_pad}),
    .d({_al_u7150_o,_al_u2848_o}),
    .f({_al_u9127_o,\biu/cache_ctrl_logic/u128_sel_is_0_o }));
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~C*B*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000110000000000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9130|exu/reg5_b31  (
    .b({_al_u9128_o,addr_ex[31]}),
    .c({_al_u9129_o,ex_exc_code[31]}),
    .clk(clk_pad),
    .d({ex_more_exception_neg_lutinv,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({_al_u9130_o,open_n69347}),
    .q({open_n69351,wb_exc_code[31]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~((D*~A)*~(B)*~(C)+(D*~A)*B*~(C)+~((D*~A))*B*C+(D*~A)*B*C)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~((D*~A)*~(B)*~(C)+(D*~A)*B*~(C)+~((D*~A))*B*C+(D*~A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0011101000111111),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0011101000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9133|exu/reg5_b22  (
    .a({_al_u9131_o,open_n69352}),
    .b({ex_more_exception_neg_lutinv,addr_ex[22]}),
    .c({_al_u2910_o,ex_exc_code[22]}),
    .clk(clk_pad),
    .d({\exu/main_state [3],ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({_al_u9133_o,open_n69370}),
    .q({open_n69374,wb_exc_code[22]}));  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*B*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"))
    \_al_u9136|_al_u2852  (
    .b({_al_u2852_o,open_n69377}),
    .c({amo,shift_r}),
    .d({_al_u9135_o,shift_l}),
    .f({\exu/n138_lutinv ,_al_u2852_o}));
  // ../../RTL/CPU/EX/exu.v(268)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*D)"),
    //.LUT1("(~C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111111),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9137|exu/reg8_b3  (
    .b({_al_u2852_o,open_n69400}),
    .c({\exu/n138_lutinv ,_al_u9137_o}),
    .ce(ex_nop),
    .clk(clk_pad),
    .d({_al_u9134_o,_al_u9133_o}),
    .sr(rst_pad),
    .f({_al_u9137_o,open_n69413}),
    .q({open_n69417,\exu/main_state [3]}));  // ../../RTL/CPU/EX/exu.v(268)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u9141|_al_u9143  (
    .a({\exu/shift_count [4],open_n69418}),
    .b({\exu/shift_count [5],_al_u9141_o}),
    .c({\exu/shift_count [6],_al_u9142_o}),
    .d({\exu/shift_count [7],_al_u2855_o}),
    .f({_al_u9141_o,\exu/shift_multi_ready }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(~D*~(~C*B))"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"))
    \_al_u9144|_al_u9142  (
    .a({open_n69439,\exu/shift_count [0]}),
    .b({\exu/shift_multi_ready ,\exu/shift_count [1]}),
    .c({_al_u2852_o,\exu/shift_count [2]}),
    .d({\exu/n138_lutinv ,\exu/shift_count [3]}),
    .f({_al_u9144_o,_al_u9142_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*~A)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(~D*~C*B*~A)"),
    //.LUTG1("(~D*~C*B*A)"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000000000000100),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9145|_al_u9139  (
    .a({\exu/main_state [0],\exu/main_state [0]}),
    .b({\exu/main_state [1],\exu/main_state [1]}),
    .c({\exu/main_state [2],\exu/main_state [2]}),
    .d({\exu/main_state [3],\exu/main_state [3]}),
    .f({\exu/c_load_1_lutinv ,_al_u9139_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~D)"),
    //.LUTF1("(B*~(D*~(~C*~A)))"),
    //.LUTG0("(C*B*~D)"),
    //.LUTG1("(B*~(D*~(~C*~A)))"),
    .INIT_LUTF0(16'b0000000011000000),
    .INIT_LUTF1(16'b0000010011001100),
    .INIT_LUTG0(16'b0000000011000000),
    .INIT_LUTG1(16'b0000010011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9146|_al_u9140  (
    .a({\exu/n10 ,open_n69484}),
    .b({_al_u9144_o,_al_u3224_o}),
    .c({\exu/c_load_1_lutinv ,_al_u9139_o}),
    .d({load,\biu/cache_ctrl_logic/n100 [4]}),
    .f({_al_u9146_o,\exu/n10 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000001100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9147|_al_u9135  (
    .b({open_n69511,load}),
    .c({_al_u9121_o,store}),
    .d({\exu/c_fence_lutinv ,_al_u9121_o}),
    .f({_al_u9147_o,_al_u9135_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~B*~D))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .INIT_LUT0(16'b1111000011000000),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"))
    \_al_u9148|_al_u6256  (
    .a({_al_u6254_o,open_n69532}),
    .b({_al_u6255_o,_al_u6255_o}),
    .c({amo,store}),
    .d({store,_al_u6254_o}),
    .f({_al_u9148_o,write}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*~(B*A)))"),
    //.LUTF1("(B*~(~A*~(D*~C)))"),
    //.LUTG0("(C*~(D*~(B*A)))"),
    //.LUTG1("(B*~(~A*~(D*~C)))"),
    .INIT_LUTF0(16'b1000000011110000),
    .INIT_LUTF1(16'b1000110010001000),
    .INIT_LUTG0(16'b1000000011110000),
    .INIT_LUTG1(16'b1000110010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9149|_al_u9128  (
    .a({_al_u9128_o,_al_u6426_o}),
    .b({_al_u9146_o,_al_u9126_o}),
    .c({_al_u9147_o,_al_u9127_o}),
    .d({_al_u9148_o,\biu/cache_ctrl_logic/n55_lutinv }),
    .f({_al_u9149_o,_al_u9128_o}));
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9152|exu/reg5_b21  (
    .b({_al_u9129_o,addr_ex[21]}),
    .c({_al_u2910_o,ex_exc_code[21]}),
    .clk(clk_pad),
    .d({ex_more_exception_neg_lutinv,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({_al_u9152_o,open_n69596}),
    .q({open_n69600,wb_exc_code[21]}));  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*D))"),
    //.LUT1("(~B*~(~C*~D))"),
    .INIT_LUT0(16'b0000001100001111),
    .INIT_LUT1(16'b0011001100110000),
    .MODE("LOGIC"))
    \_al_u9155|_al_u9154  (
    .b({_al_u9152_o,\exu/main_state [0]}),
    .c({_al_u9154_o,\exu/main_state [1]}),
    .d({_al_u9151_o,_al_u9153_o}),
    .f({_al_u9155_o,_al_u9154_o}));
  // ../../RTL/CPU/EX/exu.v(268)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*D))"),
    //.LUT1("(~D*~(~C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001100),
    .INIT_LUT1(16'b0000000011110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9156|exu/reg8_b1  (
    .b({\exu/n19 ,_al_u9156_o}),
    .c({load,\exu/n19 }),
    .ce(ex_nop),
    .clk(clk_pad),
    .d({\exu/n10 ,_al_u9155_o}),
    .sr(rst_pad),
    .f({_al_u9156_o,open_n69637}),
    .q({open_n69641,\exu/main_state [1]}));  // ../../RTL/CPU/EX/exu.v(268)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(B*C*~(D)+~(B)*~(C)*D))"),
    //.LUT1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b0000000101000000),
    .INIT_LUT1(16'b1011110000110000),
    .MODE("LOGIC"))
    \_al_u9158|_al_u9131  (
    .a({_al_u9130_o,_al_u9130_o}),
    .b({_al_u9153_o,\exu/main_state [0]}),
    .c({\exu/main_state [0],\exu/main_state [1]}),
    .d({\exu/main_state [1],\exu/main_state [2]}),
    .f({_al_u9158_o,_al_u9131_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9159|_al_u9151  (
    .c({\exu/shift_multi_ready ,_al_u6255_o}),
    .d({_al_u9158_o,_al_u9130_o}),
    .f({_al_u9159_o,_al_u9151_o}));
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000001111001111),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000001111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9160|exu/reg5_b59  (
    .b({_al_u2910_o,open_n69692}),
    .c({_al_u9139_o,addr_ex[59]}),
    .clk(clk_pad),
    .d({ex_more_exception_neg_lutinv,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({_al_u9160_o,open_n69710}),
    .q({open_n69714,wb_exc_code[59]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(268)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~B*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("~(~C*~B*~D)"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111100),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111111111111100),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9161|exu/reg8_b0  (
    .b({open_n69717,_al_u9161_o}),
    .c({_al_u9128_o,_al_u9162_o}),
    .ce(ex_nop),
    .clk(clk_pad),
    .d({_al_u9160_o,_al_u9159_o}),
    .sr(rst_pad),
    .f({_al_u9161_o,open_n69734}),
    .q({open_n69738,\exu/main_state [0]}));  // ../../RTL/CPU/EX/exu.v(268)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9162|_al_u9134  (
    .b({open_n69741,load}),
    .c({_al_u2852_o,store}),
    .d({_al_u9134_o,\exu/n19 }),
    .f({_al_u9162_o,_al_u9134_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B*~D)"),
    //.LUT1("~(C@D)"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b1111000000001111),
    .MODE("LOGIC"))
    \_al_u9165|_al_u2691  (
    .b({open_n69768,wb_rd_index[3]}),
    .c({wb_rd_index[2],wb_rd_index[4]}),
    .d({id_rs2_index[2],wb_rd_index[2]}),
    .f({_al_u9165_o,_al_u2691_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~D)"),
    //.LUTF1("(D*B*~(C*~A))"),
    //.LUTG0("~(C*~D)"),
    //.LUTG1("(D*B*~(C*~A))"),
    .INIT_LUTF0(16'b1111111100001111),
    .INIT_LUTF1(16'b1000110000000000),
    .INIT_LUTG0(16'b1111111100001111),
    .INIT_LUTG1(16'b1000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9166|_al_u2689  (
    .a({id_rs2_index[4],open_n69789}),
    .b({_al_u5144_o,open_n69790}),
    .c({wb_rd_index[4],id_valid}),
    .d({id_valid,rst_pad}),
    .f({_al_u9166_o,\ins_dec/n107 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C@B)*~(~D*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(C@B)*~(~D*A))"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1100001101000001),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1100001101000001),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9168|_al_u9164  (
    .a({_al_u9164_o,id_rs2_index[4]}),
    .b({_al_u9165_o,id_rs2_index[0]}),
    .c({_al_u9166_o,wb_rd_index[0]}),
    .d({_al_u9167_o,wb_rd_index[4]}),
    .f({_al_u9168_o,_al_u9164_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*D)"),
    //.LUTF1("(D*~(~C*~B*A))"),
    //.LUTG0("(~C*~B*D)"),
    //.LUTG1("(D*~(~C*~B*A))"),
    .INIT_LUTF0(16'b0000001100000000),
    .INIT_LUTF1(16'b1111110100000000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111110100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9169|_al_u4873  (
    .a({_al_u4872_o,open_n69839}),
    .b({id_rs1_index[4],id_rs1_index[4]}),
    .c({id_rs1_index[3],id_rs1_index[3]}),
    .d({id_valid,_al_u4872_o}),
    .f({\pip_ctrl/n34 ,\cu_ru/n45_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C@B)*~(D@A))"),
    //.LUTF1("(C@D)"),
    //.LUTG0("(~(C@B)*~(D@A))"),
    //.LUTG1("(C@D)"),
    .INIT_LUTF0(16'b1000001001000001),
    .INIT_LUTF1(16'b0000111111110000),
    .INIT_LUTG0(16'b1000001001000001),
    .INIT_LUTG1(16'b0000111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9172|_al_u9167  (
    .a({open_n69864,id_rs2_index[3]}),
    .b({open_n69865,id_rs2_index[1]}),
    .c({wb_rd_index[1],wb_rd_index[1]}),
    .d({id_rs1_index[1],wb_rd_index[3]}),
    .f({\pip_ctrl/eq2/xor_i0[1]_i1[1]_o_lutinv ,_al_u9167_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u9174|_al_u4173  (
    .c({wb_rd_index[3],id_ins[18]}),
    .d({id_ins[18],_al_u3214_o}),
    .f({_al_u9174_o,_al_u4173_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*~B*~(D@A))"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*~B*~(D@A))"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000001000000001),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000001000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9175|_al_u9173  (
    .a({id_rs1_index[2],open_n69914}),
    .b({_al_u9173_o,open_n69915}),
    .c({_al_u9174_o,wb_rd_index[4]}),
    .d({wb_rd_index[2],id_ins[19]}),
    .f({_al_u9175_o,_al_u9173_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*B)*~(D*~A))"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(~(~C*B)*~(D*~A))"),
    //.LUTG1("(D*~C*B*A)"),
    .INIT_LUTF0(16'b1010001011110011),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b1010001011110011),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9176|_al_u9171  (
    .a({_al_u9170_o,id_rs1_index[4]}),
    .b({_al_u9171_o,id_rs1_index[0]}),
    .c({\pip_ctrl/eq2/xor_i0[1]_i1[1]_o_lutinv ,wb_rd_index[0]}),
    .d({_al_u9175_o,wb_rd_index[4]}),
    .f({_al_u9176_o,_al_u9171_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~A*~(D*~B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*~A*~(D*~B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000010000000101),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9177|_al_u9189  (
    .a({open_n69964,_al_u9149_o}),
    .b({\pip_ctrl/n34 ,_al_u9177_o}),
    .c({_al_u9176_o,\pip_ctrl/id_ex_war_lutinv }),
    .d({_al_u9168_o,_al_u9188_o}),
    .f({_al_u9177_o,_al_u9189_o}));
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(~D*A))"),
    //.LUT1("(D*B*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111101000101),
    .INIT_LUT1(16'b1000110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9179|exu/reg7_b4  (
    .a({id_rs2_index[4],id_rs2_index[4]}),
    .b({_al_u5144_o,id_rs2_index[2]}),
    .c({ex_rd_index[4],ex_rd_index[2]}),
    .clk(clk_pad),
    .d({id_valid,ex_rd_index[4]}),
    .mi({open_n70000,ex_rd_index[4]}),
    .sr(rst_pad),
    .f({_al_u9179_o,_al_u9180_o}),
    .q({open_n70004,wb_rd_index[4]}));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C@B)*~(D@A))"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(~(C@B)*~(D@A))"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000001001000001),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b1000001001000001),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9181|exu/reg7_b1  (
    .a({id_rs2_index[1],id_rs1_index[4]}),
    .b({id_rs2_index[0],id_rs1_index[1]}),
    .c({ex_rd_index[0],ex_rd_index[1]}),
    .clk(clk_pad),
    .d({ex_rd_index[1],ex_rd_index[4]}),
    .mi({open_n70009,ex_rd_index[1]}),
    .sr(rst_pad),
    .f({_al_u9181_o,_al_u9183_o}),
    .q({open_n70024,wb_rd_index[1]}));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~C*B)*~(D@A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~C*B)*~(D@A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001001010001),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1010001001010001),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9182|exu/reg7_b3  (
    .a({_al_u9178_o,id_rs2_index[3]}),
    .b({_al_u9179_o,id_rs2_index[2]}),
    .c({_al_u9180_o,ex_rd_index[2]}),
    .clk(clk_pad),
    .d({_al_u9181_o,ex_rd_index[3]}),
    .mi({open_n70029,ex_rd_index[3]}),
    .sr(rst_pad),
    .f({_al_u9182_o,_al_u9178_o}),
    .q({open_n70044,wb_rd_index[3]}));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*~(~B*~(C*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1110110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9187|exu/gpr_write_reg  (
    .a({\pip_ctrl/n34 ,open_n70045}),
    .b({_al_u9182_o,open_n70046}),
    .c({\pip_ctrl/n36_lutinv ,ex_valid}),
    .clk(clk_pad),
    .d({_al_u9186_o,ex_gpr_write}),
    .mi({open_n70058,ex_gpr_write}),
    .sr(rst_pad),
    .f({\pip_ctrl/id_ex_war_lutinv ,_al_u9186_o}),
    .q({open_n70062,wb_gpr_write}));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(D*~(C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0111111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9194|exu/reg5_b47  (
    .a({ex_more_exception_neg_lutinv,open_n70063}),
    .b({_al_u9193_o,open_n70064}),
    .c({\exu/n17_lutinv ,addr_ex[47]}),
    .clk(clk_pad),
    .d({ex_valid,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .f({\pip_ctrl/ex_exception ,open_n70078}),
    .q({open_n70082,wb_exc_code[47]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*~B*~A))"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(D*~(C*~B*~A))"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110111100000000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1110111100000000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u9195|ins_dec/valid_reg  (
    .a({open_n70083,id_ill_ins}),
    .b({\pip_ctrl/ex_exception ,\ins_dec/n302 }),
    .c({ex_nop,_al_u9190_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\pip_ctrl/id_exception ,id_valid}),
    .mi({open_n70087,id_valid}),
    .sr(\ins_dec/u478_sel_is_0_o ),
    .f({_al_u9195_o,\pip_ctrl/id_exception }),
    .q({open_n70102,ex_valid}));  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u9197|_al_u3928  (
    .c({ex_nop,_al_u2932_o}),
    .d({\pip_ctrl/ex_exception ,_al_u2931_o}),
    .f({_al_u9197_o,_al_u3928_o}));
  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*A*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000100000001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9198|ins_dec/ins_acc_fault_reg  (
    .a({_al_u9197_o,open_n70127}),
    .b({_al_u9177_o,open_n70128}),
    .c({\pip_ctrl/id_ex_war_lutinv ,_al_u9197_o}),
    .ce(\ins_dec/u461_sel_is_0_o ),
    .clk(clk_pad),
    .d({_al_u9188_o,_al_u9189_o}),
    .mi({open_n70139,id_ins_acc_fault}),
    .sr(\ins_dec/n107 ),
    .f({id_nop_neg_lutinv,\ins_dec/u461_sel_is_0_o }),
    .q({open_n70143,ex_ins_acc_fault}));  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u9199|_al_u9200  (
    .c({_al_u9149_o,\ins_dec/n107 }),
    .d({id_nop_neg_lutinv,id_nop_neg_lutinv}),
    .f({id_hold,\ins_dec/u478_sel_is_0_o }));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9204|ins_fetch/reg0_b0  (
    .c({_al_u9195_o,_al_u9195_o}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u9189_o,_al_u9189_o}),
    .mi({open_n70175,addr_if[0]}),
    .sr(rst_pad),
    .f({_al_u9204_o,if_hold}),
    .q({open_n70190,id_ins_pc[0]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9207|biu/cache_ctrl_logic/reg0_b24  (
    .a({\biu/cache_ctrl_logic/l1i_va [18],\ins_fetch/n27 }),
    .b({\biu/cache_ctrl_logic/l1i_va [24],pip_flush}),
    .c({addr_if[18],\ins_fetch/n1 [22]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[24],addr_if[24]}),
    .mi({open_n70194,addr_if[24]}),
    .sr(rst_pad),
    .f({_al_u9207_o,_al_u9579_o}),
    .q({open_n70209,\biu/cache_ctrl_logic/l1i_va [24]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9209|ins_fetch/reg0_b58  (
    .a({_al_u9205_o,\biu/cache_ctrl_logic/l1i_va [13]}),
    .b({_al_u9206_o,\biu/cache_ctrl_logic/l1i_va [58]}),
    .c({_al_u9207_o,addr_if[13]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u9208_o,addr_if[58]}),
    .mi({open_n70213,addr_if[58]}),
    .sr(rst_pad),
    .f({_al_u9209_o,_al_u9205_o}),
    .q({open_n70228,id_ins_pc[58]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u9218|_al_u6725  (
    .a({_al_u9214_o,open_n70229}),
    .b({_al_u9215_o,open_n70230}),
    .c({_al_u9216_o,_al_u2837_o}),
    .d({_al_u9217_o,_al_u2835_o}),
    .f({_al_u9218_o,_al_u6725_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9219|biu/cache_ctrl_logic/reg3_b17  (
    .a({\biu/cache_ctrl_logic/l1i_va [17],\biu/cache_ctrl_logic/l1i_va [17]}),
    .b({\biu/cache_ctrl_logic/l1i_va [21],\biu/cache_ctrl_logic/l1i_va [24]}),
    .c({addr_if[17],addr_ex[17]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_if[21],addr_ex[24]}),
    .mi({open_n70261,addr_ex[17]}),
    .sr(rst_pad),
    .f({_al_u9219_o,_al_u6418_o}),
    .q({open_n70265,\biu/cache_ctrl_logic/l1d_va [17]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9221|biu/cache_ctrl_logic/reg0_b44  (
    .a({\biu/cache_ctrl_logic/l1i_va [32],\ins_fetch/n27 }),
    .b({\biu/cache_ctrl_logic/l1i_va [44],pip_flush}),
    .c({addr_if[32],\ins_fetch/n1 [42]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[44],addr_if[44]}),
    .mi({open_n70269,addr_if[44]}),
    .sr(rst_pad),
    .f({_al_u9221_o,_al_u9437_o}),
    .q({open_n70284,\biu/cache_ctrl_logic/l1i_va [44]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9222|biu/cache_ctrl_logic/reg0_b30  (
    .a({\biu/cache_ctrl_logic/l1i_va [16],\ins_fetch/n27 }),
    .b({\biu/cache_ctrl_logic/l1i_va [30],pip_flush}),
    .c({addr_if[16],\ins_fetch/n1 [28]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[30],addr_if[30]}),
    .mi({open_n70295,addr_if[30]}),
    .sr(rst_pad),
    .f({_al_u9222_o,_al_u9537_o}),
    .q({open_n70299,\biu/cache_ctrl_logic/l1i_va [30]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9228|biu/cache_ctrl_logic/reg3_b60  (
    .a({_al_u9224_o,open_n70300}),
    .b({_al_u9225_o,\biu/cache_ctrl_logic/l1i_va [60]}),
    .c({_al_u9226_o,addr_ex[60]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u9227_o,_al_u6396_o}),
    .mi({open_n70304,addr_ex[60]}),
    .sr(rst_pad),
    .f({_al_u9228_o,_al_u6397_o}),
    .q({open_n70319,\biu/cache_ctrl_logic/l1d_va [60]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*~C))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000010001000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9229|ins_fetch/reg0_b37  (
    .a({_al_u9211_o,_al_u9209_o}),
    .b({_al_u9218_o,_al_u9210_o}),
    .c({_al_u9223_o,\biu/cache_ctrl_logic/l1i_va [37]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u9228_o,addr_if[37]}),
    .mi({open_n70330,addr_if[37]}),
    .sr(rst_pad),
    .f({_al_u9229_o,_al_u9211_o}),
    .q({open_n70334,id_ins_pc[37]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9238|ins_fetch/reg0_b20  (
    .a({open_n70335,\biu/cache_ctrl_logic/l1i_va [20]}),
    .b({_al_u9236_o,\biu/cache_ctrl_logic/l1i_va [56]}),
    .c({_al_u9237_o,addr_if[20]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u9235_o,addr_if[56]}),
    .mi({open_n70346,addr_if[20]}),
    .sr(rst_pad),
    .f({_al_u9238_o,_al_u9236_o}),
    .q({open_n70350,id_ins_pc[20]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(B*A*~(D@C))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000001000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9242|ins_fetch/reg0_b27  (
    .a({open_n70351,_al_u9231_o}),
    .b({_al_u9238_o,_al_u9232_o}),
    .c({_al_u9241_o,\biu/cache_ctrl_logic/l1i_va [27]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u9233_o,addr_if[27]}),
    .mi({open_n70362,addr_if[27]}),
    .sr(rst_pad),
    .f({_al_u9242_o,_al_u9233_o}),
    .q({open_n70366,id_ins_pc[27]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9244|biu/cache_ctrl_logic/reg0_b42  (
    .a({open_n70367,\ins_fetch/n27 }),
    .b({open_n70368,pip_flush}),
    .c({addr_if[42],\ins_fetch/n1 [40]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_va [42],addr_if[42]}),
    .mi({open_n70372,addr_if[42]}),
    .sr(rst_pad),
    .f({_al_u9244_o,_al_u9449_o}),
    .q({open_n70387,\biu/cache_ctrl_logic/l1i_va [42]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9250|_al_u9264  (
    .a({_al_u9246_o,_al_u9229_o}),
    .b({_al_u9247_o,_al_u9242_o}),
    .c({_al_u9248_o,_al_u9253_o}),
    .d({_al_u9249_o,_al_u9263_o}),
    .f({_al_u9250_o,_al_u9264_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100110001),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9253|biu/cache_ctrl_logic/reg3_b40  (
    .a({_al_u9245_o,\biu/cache_ctrl_logic/l1i_va [40]}),
    .b({_al_u9250_o,\biu/cache_ctrl_logic/l1i_va [50]}),
    .c({_al_u9251_o,addr_ex[40]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u9252_o,addr_ex[50]}),
    .mi({open_n70422,addr_ex[40]}),
    .sr(rst_pad),
    .f({_al_u9253_o,_al_u6417_o}),
    .q({open_n70426,\biu/cache_ctrl_logic/l1d_va [40]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9258|ins_fetch/reg0_b54  (
    .a({_al_u9254_o,\biu/cache_ctrl_logic/l1i_va [54]}),
    .b({_al_u9255_o,\biu/cache_ctrl_logic/l1i_va [62]}),
    .c({_al_u9256_o,addr_if[54]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u9257_o,addr_if[62]}),
    .mi({open_n70430,addr_if[54]}),
    .sr(rst_pad),
    .f({_al_u9258_o,_al_u9257_o}),
    .q({open_n70445,id_ins_pc[54]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9263|ins_fetch/reg0_b52  (
    .a({_al_u9258_o,open_n70446}),
    .b({_al_u9260_o,\biu/cache_ctrl_logic/l1i_va [52]}),
    .c({_al_u9261_o,addr_if[52]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u9262_o,_al_u9259_o}),
    .mi({open_n70450,addr_if[52]}),
    .sr(rst_pad),
    .f({_al_u9263_o,_al_u9260_o}),
    .q({open_n70465,id_ins_pc[52]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*~D)"),
    //.LUTF1("(~C*B*~(D*A))"),
    //.LUTG0("(~C*B*~D)"),
    //.LUTG1("(~C*B*~(D*A))"),
    .INIT_LUTF0(16'b0000000000001100),
    .INIT_LUTF1(16'b0000010000001100),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000010000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9265|_al_u6317  (
    .a({\biu/bus_unit/mmu/n7_lutinv ,open_n70466}),
    .b({_al_u6319_o,priv[1]}),
    .c({\biu/bus_unit/mmu/n8_lutinv ,priv[3]}),
    .d({\biu/cache_ctrl_logic/l1i_pte [4],priv[0]}),
    .f({_al_u9265_o,\biu/bus_unit/mmu/n8_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(C*~B*D)"),
    .INIT_LUT0(16'b1100111011101010),
    .INIT_LUT1(16'b0011000000000000),
    .MODE("LOGIC"))
    \_al_u9266|_al_u7151  (
    .a({open_n70491,_al_u2835_o}),
    .b({\biu/cache_ctrl_logic/statu [0],_al_u2838_o}),
    .c(\biu/cache_ctrl_logic/statu [1:0]),
    .d({_al_u2838_o,\biu/cache_ctrl_logic/statu [1]}),
    .f({_al_u9266_o,_al_u7151_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*B*~(D*~A))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*B*~(D*~A))"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b1000000011000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b1000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9270|_al_u9271  (
    .a({\biu/cache_ctrl_logic/n100 [4],open_n70512}),
    .b({_al_u7149_o,open_n70513}),
    .c({_al_u4399_o,_al_u3224_o}),
    .d({\biu/cache_ctrl_logic/l1i_pte [7],_al_u9270_o}),
    .f({_al_u9270_o,_al_u9271_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~C*~(D*B)))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1010100010100000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u9275|_al_u9273  (
    .a({open_n70538,\biu/cache_ctrl_logic/n100 [4]}),
    .b({_al_u9274_o,_al_u7149_o}),
    .c({\biu/cache_ctrl_logic/statu [3],_al_u3945_o}),
    .d({_al_u9273_o,_al_u7150_o}),
    .f({_al_u9275_o,_al_u9273_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(A*~(~D*~(C*~B)))"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b1010101000100000),
    .MODE("LOGIC"))
    \_al_u9276|_al_u9272  (
    .a({_al_u9271_o,open_n70559}),
    .b({_al_u9272_o,\biu/cache_ctrl_logic/n97_lutinv }),
    .c({_al_u9275_o,\biu/cache_ctrl_logic/l1d_pte [7]}),
    .d({_al_u4399_o,\biu/cache_ctrl_logic/n100 [4]}),
    .f({_al_u9276_o,_al_u9272_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~D))"),
    //.LUTF1("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("(~C*~(B*~D))"),
    //.LUTG1("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .INIT_LUTF0(16'b0000111100000011),
    .INIT_LUTF1(16'b1100111100000011),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b1100111100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9279|_al_u9277  (
    .b({_al_u9277_o,_al_u3224_o}),
    .c({_al_u9278_o,_al_u4834_o}),
    .d({_al_u9276_o,_al_u7163_o}),
    .f({_al_u9279_o,_al_u9277_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(~B*~(~C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u9282|biu/cache_ctrl_logic/reg8_b3  (
    .b({_al_u7193_o,_al_u9284_o}),
    .c({_al_u7162_o,_al_u9287_o}),
    .clk(clk_pad),
    .d({_al_u9281_o,\biu/cache_ctrl_logic/n128 [3]}),
    .sr(\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ),
    .f({\biu/cache_ctrl_logic/n128 [3],open_n70621}),
    .q({open_n70625,\biu/cache_ctrl_logic/statu [3]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9287|_al_u9286  (
    .c({_al_u9286_o,\biu/cache_ctrl_logic/l1i_pte [7]}),
    .d({_al_u9285_o,_al_u7162_o}),
    .f({_al_u9287_o,_al_u9286_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u9291|_al_u9290  (
    .a({open_n70654,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({open_n70655,\cu_ru/trap_target_m }),
    .c({_al_u4138_o,\cu_ru/stvec [0]}),
    .d({_al_u9290_o,\cu_ru/mtvec [0]}),
    .f({\cu_ru/mux34_b0_sel_is_2_o ,_al_u9290_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000000100001011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u9292|_al_u9559  (
    .a({open_n70676,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [13],\cu_ru/tvec [29]}),
    .c({\cu_ru/n43 [9],_al_u6055_o}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/n43 [25]}),
    .f({_al_u9292_o,_al_u9559_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9293|ins_fetch/reg2_b11  (
    .a({_al_u9292_o,_al_u9289_o}),
    .b({_al_u6055_o,_al_u9293_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[11],_al_u9294_o}),
    .sr(rst_pad),
    .f({_al_u9293_o,open_n70714}),
    .q({open_n70718,addr_if[11]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT_LUTF0(16'b0001010110111111),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9294|_al_u9516  (
    .a({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [11],\cu_ru/sepc [33]}),
    .d({\cu_ru/mepc [11],\cu_ru/mepc [33]}),
    .f({_al_u9294_o,_al_u9516_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9296|ins_fetch/reg2_b60  (
    .a({\ins_fetch/n27 ,_al_u9330_o}),
    .b({pip_flush,_al_u9332_o}),
    .c({\ins_fetch/n1 [8],pip_flush}),
    .clk(clk_pad),
    .d({addr_if[10],_al_u9333_o}),
    .sr(rst_pad),
    .f({_al_u9296_o,open_n70756}),
    .q({open_n70760,addr_if[60]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u9297|_al_u9665  (
    .b({\cu_ru/tvec [12],\cu_ru/tvec [14]}),
    .c({\cu_ru/n43 [8],\cu_ru/n43 [10]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .f({_al_u9297_o,_al_u9665_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000111000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9298|ins_fetch/reg2_b10  (
    .a({_al_u9297_o,_al_u9296_o}),
    .b({_al_u6055_o,_al_u9298_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[10],_al_u9299_o}),
    .sr(rst_pad),
    .f({_al_u9298_o,open_n70796}),
    .q({open_n70800,addr_if[10]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUT1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT_LUT0(16'b0001010110111111),
    .INIT_LUT1(16'b0001010110111111),
    .MODE("LOGIC"))
    \_al_u9299|_al_u9497  (
    .a({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [10],\cu_ru/sepc [36]}),
    .d({\cu_ru/mepc [10],\cu_ru/mepc [36]}),
    .f({_al_u9299_o,_al_u9497_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u9302|_al_u9646  (
    .b({\cu_ru/tvec [11],\cu_ru/tvec [17]}),
    .c({\cu_ru/n43 [7],\cu_ru/n43 [13]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .f({_al_u9302_o,_al_u9646_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9303|ins_fetch/reg2_b9  (
    .a({_al_u9302_o,_al_u9301_o}),
    .b({_al_u6055_o,_al_u9303_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[9],_al_u9304_o}),
    .sr(rst_pad),
    .f({_al_u9303_o,open_n70860}),
    .q({open_n70864,addr_if[9]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUT1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT_LUT0(16'b0001010110111111),
    .INIT_LUT1(16'b0001010110111111),
    .MODE("LOGIC"))
    \_al_u9304|_al_u9402  (
    .a({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [9],\cu_ru/sepc [50]}),
    .d({\cu_ru/mepc [9],\cu_ru/mepc [50]}),
    .f({_al_u9304_o,_al_u9402_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9307|_al_u6054  (
    .a({open_n70885,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [10],\cu_ru/trap_target_m }),
    .c({\cu_ru/n43 [6],\cu_ru/stvec [10]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mtvec [10]}),
    .f({_al_u9307_o,\cu_ru/tvec [10]}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9308|ins_fetch/reg2_b8  (
    .a({_al_u9307_o,_al_u9306_o}),
    .b({_al_u6055_o,_al_u9308_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[8],_al_u9309_o}),
    .sr(rst_pad),
    .f({_al_u9308_o,open_n70927}),
    .q({open_n70931,addr_if[8]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9309|cu_ru/m_s_scratch/reg0_b8  (
    .a({\cu_ru/m_s_status/n2 ,open_n70932}),
    .b({_al_u2844_o,\cu_ru/sepc [8]}),
    .c({\cu_ru/sepc [8],data_csr[8]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [8],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n70936,data_csr[8]}),
    .sr(rst_pad),
    .f({_al_u9309_o,_al_u5361_o}),
    .q({open_n70951,\cu_ru/mscratch [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001110100111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001110100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9312|_al_u6055  (
    .a({_al_u6055_o,open_n70952}),
    .b({_al_u2844_o,open_n70953}),
    .c({\cu_ru/sepc [63],_al_u5157_o}),
    .d({new_pc[63],\cu_ru/trap_target_m }),
    .f({_al_u9312_o,_al_u6055_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(A*~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C))"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(A*~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000100010101000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000100010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9313|ins_fetch/reg2_b63  (
    .a({pip_flush,open_n70978}),
    .b({_al_u9312_o,open_n70979}),
    .c({\cu_ru/m_s_status/n2 ,_al_u9313_o}),
    .clk(clk_pad),
    .d({\cu_ru/mepc [63],_al_u9311_o}),
    .sr(rst_pad),
    .f({_al_u9313_o,open_n70997}),
    .q({open_n71001,addr_if[63]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUT1("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT_LUT0(16'b0000000100001011),
    .INIT_LUT1(16'b0001001111011111),
    .MODE("LOGIC"))
    \_al_u9315|_al_u9670  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({_al_u6055_o,\cu_ru/tvec [4]}),
    .c({\cu_ru/add0_2_co ,_al_u6055_o}),
    .d({new_pc[62],\cu_ru/n43 [0]}),
    .f({_al_u9315_o,_al_u9670_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~B*~(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000001000110010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9316|cu_ru/m_s_scratch/reg0_b62  (
    .a({_al_u9315_o,open_n71022}),
    .b({\cu_ru/m_s_status/n2 ,\cu_ru/sepc [62]}),
    .c({_al_u2844_o,data_csr[62]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [62],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n71033,data_csr[62]}),
    .sr(rst_pad),
    .f({_al_u9316_o,_al_u5373_o}),
    .q({open_n71037,\cu_ru/mscratch [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*~D))"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("~(~B*~(C*~D))"),
    //.LUTG1("(D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011111100),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b1100110011111100),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9318|ins_fetch/reg2_b62  (
    .b({\cu_ru/m_s_status/n2 ,_al_u9317_o}),
    .c({\cu_ru/mepc [62],_al_u9318_o}),
    .clk(clk_pad),
    .d({pip_flush,_al_u9316_o}),
    .sr(rst_pad),
    .f({_al_u9318_o,open_n71057}),
    .q({open_n71061,addr_if[62]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9321|_al_u9620  (
    .b({\cu_ru/tvec [9],\cu_ru/tvec [21]}),
    .c({\cu_ru/n43 [5],\cu_ru/n43 [17]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .f({_al_u9321_o,_al_u9620_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000111000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9322|ins_fetch/reg2_b7  (
    .a({_al_u9321_o,_al_u9320_o}),
    .b({_al_u6055_o,_al_u9322_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[7],_al_u9323_o}),
    .sr(rst_pad),
    .f({_al_u9322_o,open_n71101}),
    .q({open_n71105,addr_if[7]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT_LUTF0(16'b0001010110111111),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9323|_al_u9338  (
    .a({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [7],\cu_ru/sepc [59]}),
    .d({\cu_ru/mepc [7],\cu_ru/mepc [59]}),
    .f({_al_u9323_o,_al_u9338_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9326|_al_u5998  (
    .a({open_n71130,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [63],\cu_ru/trap_target_m }),
    .c({\cu_ru/n43 [59],\cu_ru/stvec [63]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mtvec [63]}),
    .f({_al_u9326_o,\cu_ru/tvec [63]}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9327|ins_fetch/reg2_b61  (
    .a({_al_u9326_o,_al_u9325_o}),
    .b({_al_u6055_o,_al_u9327_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[61],_al_u9328_o}),
    .sr(rst_pad),
    .f({_al_u9327_o,open_n71172}),
    .q({open_n71176,addr_if[61]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010110111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9328|cu_ru/m_s_scratch/reg0_b61  (
    .a({\cu_ru/m_s_status/n2 ,open_n71177}),
    .b({_al_u2844_o,\cu_ru/sepc [61]}),
    .c({\cu_ru/sepc [61],data_csr[61]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [61],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n71188,data_csr[61]}),
    .sr(rst_pad),
    .f({_al_u9328_o,_al_u5377_o}),
    .q({open_n71192,\cu_ru/mscratch [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9331|_al_u5999  (
    .a({open_n71193,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [62],\cu_ru/trap_target_m }),
    .c({\cu_ru/n43 [58],\cu_ru/stvec [62]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mtvec [62]}),
    .f({_al_u9331_o,\cu_ru/tvec [62]}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9333|cu_ru/m_s_scratch/reg0_b60  (
    .a({\cu_ru/m_s_status/n2 ,open_n71218}),
    .b({_al_u2844_o,\cu_ru/sepc [60]}),
    .c({\cu_ru/sepc [60],data_csr[60]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [60],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n71222,data_csr[60]}),
    .sr(rst_pad),
    .f({_al_u9333_o,_al_u5381_o}),
    .q({open_n71237,\cu_ru/mscratch [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9336|_al_u9587  (
    .b({\cu_ru/tvec [61],\cu_ru/tvec [25]}),
    .c({\cu_ru/n43 [57],\cu_ru/n43 [21]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .f({_al_u9336_o,_al_u9587_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000111000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9337|ins_fetch/reg2_b59  (
    .a({_al_u9336_o,_al_u9335_o}),
    .b({_al_u6055_o,_al_u9337_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[59],_al_u9338_o}),
    .sr(rst_pad),
    .f({_al_u9337_o,open_n71277}),
    .q({open_n71281,addr_if[59]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*A))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b1110110010100000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u9341|_al_u6001  (
    .a({open_n71282,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [60],\cu_ru/trap_target_m }),
    .c({\cu_ru/n43 [56],\cu_ru/stvec [60]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mtvec [60]}),
    .f({_al_u9341_o,\cu_ru/tvec [60]}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9342|ins_fetch/reg2_b58  (
    .a({_al_u9341_o,_al_u9340_o}),
    .b({_al_u6055_o,_al_u9342_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[58],_al_u9343_o}),
    .sr(rst_pad),
    .f({_al_u9342_o,open_n71320}),
    .q({open_n71324,addr_if[58]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010110111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9343|cu_ru/m_s_scratch/reg1_b58  (
    .a({\cu_ru/m_s_status/n2 ,open_n71325}),
    .b({_al_u2844_o,\cu_ru/sepc [58]}),
    .c({\cu_ru/sepc [58],data_csr[58]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [58],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n71336,data_csr[58]}),
    .sr(rst_pad),
    .f({_al_u9343_o,_al_u5393_o}),
    .q({open_n71340,\cu_ru/sscratch [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b0000000100001011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9346|_al_u9658  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [59],\cu_ru/tvec [15]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [55],\cu_ru/n43 [11]}),
    .f({_al_u9346_o,_al_u9658_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u9347|_al_u9491  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({new_pc[57],\cu_ru/sepc [37]}),
    .d({_al_u6055_o,\cu_ru/m_s_status/n2 }),
    .f({_al_u9347_o,_al_u9491_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u9348|cu_ru/m_s_cause/reg1_b57  (
    .a({open_n71383,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({open_n71384,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [57],\cu_ru/mepc [57]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,data_csr[57]}),
    .mi({open_n71395,data_csr[57]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u9348_o,_al_u6592_o}),
    .q({open_n71399,\cu_ru/mcause [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9349|cu_ru/m_s_epc/reg0_b57  (
    .b({_al_u2844_o,_al_u5157_o}),
    .c({\cu_ru/sepc [57],_al_u5397_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/n2 [57]}),
    .sr(rst_pad),
    .f({_al_u9349_o,open_n71418}),
    .q({open_n71422,\cu_ru/sepc [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9350|ins_fetch/reg2_b57  (
    .a({_al_u9346_o,open_n71423}),
    .b({_al_u9347_o,_al_u9350_o}),
    .c({_al_u9348_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9349_o,_al_u9345_o}),
    .sr(rst_pad),
    .f({_al_u9350_o,open_n71437}),
    .q({open_n71441,addr_if[57]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b1110110010100000),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9353|_al_u6004  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [58],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [58]}),
    .d({\cu_ru/n43 [54],\cu_ru/mtvec [58]}),
    .f({_al_u9353_o,\cu_ru/tvec [58]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9354|_al_u9659  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({new_pc[56],new_pc[13]}),
    .d({_al_u6055_o,_al_u6055_o}),
    .f({_al_u9354_o,_al_u9659_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9355|_al_u9672  (
    .c({\cu_ru/mepc [56],\cu_ru/mepc [2]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9355_o,_al_u9672_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9356|_al_u9654  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [56],\cu_ru/sepc [14]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9356_o,_al_u9654_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9357|ins_fetch/reg2_b56  (
    .a({_al_u9353_o,open_n71538}),
    .b({_al_u9354_o,_al_u9357_o}),
    .c({_al_u9355_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9356_o,_al_u9352_o}),
    .sr(rst_pad),
    .f({_al_u9357_o,open_n71556}),
    .q({open_n71560,addr_if[56]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9360|_al_u6005  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [57],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [57]}),
    .d({\cu_ru/n43 [53],\cu_ru/mtvec [57]}),
    .f({_al_u9360_o,\cu_ru/tvec [57]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9361|_al_u9652  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({new_pc[55],new_pc[14]}),
    .d({_al_u6055_o,_al_u6055_o}),
    .f({_al_u9361_o,_al_u9652_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9362|_al_u9660  (
    .c({\cu_ru/mepc [55],\cu_ru/mepc [13]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9362_o,_al_u9660_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9363|cu_ru/m_s_scratch/reg1_b55  (
    .b({_al_u2844_o,\cu_ru/sepc [55]}),
    .c({\cu_ru/sepc [55],data_csr[55]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n71651,data_csr[55]}),
    .sr(rst_pad),
    .f({_al_u9363_o,_al_u5405_o}),
    .q({open_n71655,\cu_ru/sscratch [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9364|ins_fetch/reg2_b55  (
    .a({_al_u9360_o,open_n71656}),
    .b({_al_u9361_o,_al_u9364_o}),
    .c({_al_u9362_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9363_o,_al_u9359_o}),
    .sr(rst_pad),
    .f({_al_u9364_o,open_n71674}),
    .q({open_n71678,addr_if[55]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9367|_al_u6006  (
    .a({open_n71679,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [56],\cu_ru/trap_target_m }),
    .c({\cu_ru/n43 [52],\cu_ru/stvec [56]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mtvec [56]}),
    .f({_al_u9367_o,\cu_ru/tvec [56]}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9368|ins_fetch/reg2_b54  (
    .a({_al_u9367_o,_al_u9366_o}),
    .b({_al_u6055_o,_al_u9368_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[54],_al_u9369_o}),
    .sr(rst_pad),
    .f({_al_u9368_o,open_n71721}),
    .q({open_n71725,addr_if[54]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u9369|cu_ru/m_s_cause/reg1_b54  (
    .a({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2844_o,\cu_ru/trap_target_m }),
    .c({\cu_ru/sepc [54],\cu_ru/mepc [54]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [54],data_csr[54]}),
    .mi({open_n71729,data_csr[54]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u9369_o,_al_u6598_o}),
    .q({open_n71744,\cu_ru/mcause [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b0000000100001011),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b0000000100001011),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9372|_al_u9651  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [55],\cu_ru/tvec [16]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [51],\cu_ru/n43 [12]}),
    .f({_al_u9372_o,_al_u9651_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u9374|cu_ru/m_s_cause/reg1_b53  (
    .a({open_n71769,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({open_n71770,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [53],\cu_ru/mepc [53]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,data_csr[53]}),
    .mi({open_n71781,data_csr[53]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u9374_o,_al_u6600_o}),
    .q({open_n71785,\cu_ru/mcause [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u9375|_al_u9642  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [53],\cu_ru/sepc [16]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9375_o,_al_u9642_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9376|ins_fetch/reg2_b53  (
    .a({_al_u9372_o,open_n71808}),
    .b({_al_u9373_o,_al_u9376_o}),
    .c({_al_u9374_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9375_o,_al_u9371_o}),
    .sr(rst_pad),
    .f({_al_u9376_o,open_n71822}),
    .q({open_n71826,addr_if[53]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b0000000100001011),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b0000000100001011),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9379|_al_u9639  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [54],\cu_ru/tvec [18]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [50],\cu_ru/n43 [14]}),
    .f({_al_u9379_o,_al_u9639_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u9380|_al_u9593  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({new_pc[52],new_pc[22]}),
    .d({_al_u6055_o,_al_u6055_o}),
    .f({_al_u9380_o,_al_u9593_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9381|_al_u9641  (
    .c({\cu_ru/mepc [52],\cu_ru/mepc [16]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9381_o,_al_u9641_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u9382|_al_u9635  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [52],\cu_ru/sepc [17]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9382_o,_al_u9635_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9383|ins_fetch/reg2_b52  (
    .a({_al_u9379_o,open_n71923}),
    .b({_al_u9380_o,_al_u9383_o}),
    .c({_al_u9381_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9382_o,_al_u9378_o}),
    .sr(rst_pad),
    .f({_al_u9383_o,open_n71937}),
    .q({open_n71941,addr_if[52]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b0000000100001011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9386|_al_u9632  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [8],\cu_ru/tvec [19]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [4],\cu_ru/n43 [15]}),
    .f({_al_u9386_o,_al_u9632_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u9387|_al_u9532  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({new_pc[6],new_pc[31]}),
    .d({_al_u6055_o,_al_u6055_o}),
    .f({_al_u9387_o,_al_u9532_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9388|_al_u9634  (
    .c({\cu_ru/mepc [6],\cu_ru/mepc [17]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9388_o,_al_u9634_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9389|_al_u9616  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [6],\cu_ru/sepc [20]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9389_o,_al_u9616_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9390|ins_fetch/reg2_b6  (
    .a({_al_u9386_o,open_n72034}),
    .b({_al_u9387_o,_al_u9390_o}),
    .c({_al_u9388_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9389_o,_al_u9385_o}),
    .sr(rst_pad),
    .f({_al_u9390_o,open_n72048}),
    .q({open_n72052,addr_if[6]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b1110110010100000),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9393|_al_u6009  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [53],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [53]}),
    .d({\cu_ru/n43 [49],\cu_ru/mtvec [53]}),
    .f({_al_u9393_o,\cu_ru/tvec [53]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u9394|_al_u9489  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({new_pc[51],new_pc[37]}),
    .d({_al_u6055_o,_al_u6055_o}),
    .f({_al_u9394_o,_al_u9489_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9395|_al_u9627  (
    .c({\cu_ru/mepc [51],\cu_ru/mepc [18]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9395_o,_al_u9627_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u9396|_al_u9576  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [51],\cu_ru/sepc [25]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9396_o,_al_u9576_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9397|ins_fetch/reg2_b51  (
    .a({_al_u9393_o,open_n72141}),
    .b({_al_u9394_o,_al_u9397_o}),
    .c({_al_u9395_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9396_o,_al_u9392_o}),
    .sr(rst_pad),
    .f({_al_u9397_o,open_n72159}),
    .q({open_n72163,addr_if[51]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u9400|_al_u9526  (
    .b({\cu_ru/tvec [52],\cu_ru/tvec [6]}),
    .c({\cu_ru/n43 [48],\cu_ru/n43 [2]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .f({_al_u9400_o,_al_u9526_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000111000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9401|ins_fetch/reg2_b50  (
    .a({_al_u9400_o,_al_u9399_o}),
    .b({_al_u6055_o,_al_u9401_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[50],_al_u9402_o}),
    .sr(rst_pad),
    .f({_al_u9401_o,open_n72199}),
    .q({open_n72203,addr_if[50]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b0000000100001011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9405|_al_u9625  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [51],\cu_ru/tvec [20]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [47],\cu_ru/n43 [16]}),
    .f({_al_u9405_o,_al_u9625_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u9406|_al_u9439  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({new_pc[49],new_pc[44]}),
    .d({_al_u6055_o,_al_u6055_o}),
    .f({_al_u9406_o,_al_u9439_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9407|_al_u6887  (
    .a({open_n72246,\cu_ru/read_mepc_sel_lutinv }),
    .b({open_n72247,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/mepc [49],\cu_ru/mepc [49]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/stvec [49]}),
    .f({_al_u9407_o,_al_u6887_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9408|cu_ru/m_s_epc/reg0_b49  (
    .b({_al_u2844_o,_al_u5157_o}),
    .c({\cu_ru/sepc [49],_al_u5433_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/n2 [49]}),
    .sr(rst_pad),
    .f({_al_u9408_o,open_n72290}),
    .q({open_n72294,\cu_ru/sepc [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9409|ins_fetch/reg2_b49  (
    .a({_al_u9405_o,open_n72295}),
    .b({_al_u9406_o,_al_u9409_o}),
    .c({_al_u9407_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9408_o,_al_u9404_o}),
    .sr(rst_pad),
    .f({_al_u9409_o,open_n72313}),
    .q({open_n72317,addr_if[49]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b1110110010100000),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9412|_al_u6012  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [50],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [50]}),
    .d({\cu_ru/n43 [46],\cu_ru/mtvec [50]}),
    .f({_al_u9412_o,\cu_ru/tvec [50]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9413|_al_u9420  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c(new_pc[48:47]),
    .d({_al_u6055_o,_al_u6055_o}),
    .f({_al_u9413_o,_al_u9420_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u9414|cu_ru/m_s_cause/reg1_b48  (
    .a({open_n72364,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({open_n72365,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [48],\cu_ru/mepc [48]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,data_csr[48]}),
    .mi({open_n72376,data_csr[48]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u9414_o,_al_u6612_o}),
    .q({open_n72380,\cu_ru/mcause [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u9415|_al_u9569  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [48],\cu_ru/sepc [26]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9415_o,_al_u9569_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9416|ins_fetch/reg2_b48  (
    .a({_al_u9412_o,open_n72403}),
    .b({_al_u9413_o,_al_u9416_o}),
    .c({_al_u9414_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9415_o,_al_u9411_o}),
    .sr(rst_pad),
    .f({_al_u9416_o,open_n72421}),
    .q({open_n72425,addr_if[48]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9419|_al_u6014  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [49],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [49]}),
    .d({\cu_ru/n43 [45],\cu_ru/mtvec [49]}),
    .f({_al_u9419_o,\cu_ru/tvec [49]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9421|_al_u9615  (
    .c({\cu_ru/mepc [47],\cu_ru/mepc [20]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9421_o,_al_u9615_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9422|cu_ru/m_s_epc/reg0_b47  (
    .b({_al_u2844_o,_al_u5157_o}),
    .c({\cu_ru/sepc [47],_al_u5441_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/n2 [47]}),
    .sr(rst_pad),
    .f({_al_u9422_o,open_n72496}),
    .q({open_n72500,\cu_ru/sepc [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9423|ins_fetch/reg2_b47  (
    .a({_al_u9419_o,open_n72501}),
    .b({_al_u9420_o,_al_u9423_o}),
    .c({_al_u9421_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9422_o,_al_u9418_o}),
    .sr(rst_pad),
    .f({_al_u9423_o,open_n72519}),
    .q({open_n72523,addr_if[47]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u9426|_al_u9514  (
    .b({\cu_ru/tvec [48],\cu_ru/tvec [35]}),
    .c({\cu_ru/n43 [44],\cu_ru/n43 [31]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .f({_al_u9426_o,_al_u9514_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000111000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9427|ins_fetch/reg2_b46  (
    .a({_al_u9426_o,_al_u9425_o}),
    .b({_al_u6055_o,_al_u9427_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[46],_al_u9428_o}),
    .sr(rst_pad),
    .f({_al_u9427_o,open_n72559}),
    .q({open_n72563,addr_if[46]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u9428|cu_ru/m_s_cause/reg1_b46  (
    .a({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u2844_o,\cu_ru/trap_target_m }),
    .c({\cu_ru/sepc [46],\cu_ru/mepc [46]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [46],data_csr[46]}),
    .mi({open_n72567,data_csr[46]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u9428_o,_al_u6616_o}),
    .q({open_n72582,\cu_ru/mcause [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9431|_al_u6016  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [47],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [47]}),
    .d({\cu_ru/n43 [43],\cu_ru/mtvec [47]}),
    .f({_al_u9431_o,\cu_ru/tvec [47]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9433|_al_u9601  (
    .c({\cu_ru/mepc [45],\cu_ru/mepc [3]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9433_o,_al_u9601_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9434|cu_ru/m_s_scratch/reg1_b45  (
    .b({_al_u2844_o,\cu_ru/sepc [45]}),
    .c({\cu_ru/sepc [45],data_csr[45]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n72640,data_csr[45]}),
    .sr(rst_pad),
    .f({_al_u9434_o,_al_u5449_o}),
    .q({open_n72655,\cu_ru/sscratch [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9435|ins_fetch/reg2_b45  (
    .a({_al_u9431_o,open_n72656}),
    .b({_al_u9432_o,_al_u9435_o}),
    .c({_al_u9433_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9434_o,_al_u9430_o}),
    .sr(rst_pad),
    .f({_al_u9435_o,open_n72670}),
    .q({open_n72674,addr_if[45]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b0000000100001011),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b0000000100001011),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9438|_al_u9613  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [46],\cu_ru/tvec [22]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [42],\cu_ru/n43 [18]}),
    .f({_al_u9438_o,_al_u9613_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9440|_al_u9594  (
    .c({\cu_ru/mepc [44],\cu_ru/mepc [22]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9440_o,_al_u9594_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9441|_al_u9555  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [44],\cu_ru/sepc [28]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9441_o,_al_u9555_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9442|ins_fetch/reg2_b44  (
    .a({_al_u9438_o,open_n72749}),
    .b({_al_u9439_o,_al_u9442_o}),
    .c({_al_u9440_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9441_o,_al_u9437_o}),
    .sr(rst_pad),
    .f({_al_u9442_o,open_n72763}),
    .q({open_n72767,addr_if[44]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*A))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b1110110010100000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u9445|_al_u6018  (
    .a({open_n72768,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [45],\cu_ru/trap_target_m }),
    .c({\cu_ru/n43 [41],\cu_ru/stvec [45]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mtvec [45]}),
    .f({_al_u9445_o,\cu_ru/tvec [45]}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000111000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9446|ins_fetch/reg2_b43  (
    .a({_al_u9445_o,_al_u9444_o}),
    .b({_al_u6055_o,_al_u9446_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[43],_al_u9447_o}),
    .sr(rst_pad),
    .f({_al_u9446_o,open_n72802}),
    .q({open_n72806,addr_if[43]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9447|cu_ru/m_s_scratch/reg0_b43  (
    .a({\cu_ru/m_s_status/n2 ,open_n72807}),
    .b({_al_u2844_o,\cu_ru/sepc [43]}),
    .c({\cu_ru/sepc [43],data_csr[43]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [43],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n72811,data_csr[43]}),
    .sr(rst_pad),
    .f({_al_u9447_o,_al_u5457_o}),
    .q({open_n72826,\cu_ru/mscratch [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b1110110010100000),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9450|_al_u6019  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [44],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [44]}),
    .d({\cu_ru/n43 [40],\cu_ru/mtvec [44]}),
    .f({_al_u9450_o,\cu_ru/tvec [44]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9452|_al_u9582  (
    .c({\cu_ru/mepc [42],\cu_ru/mepc [24]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9452_o,_al_u9582_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*B))"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~D*~(C*B))"),
    //.LUTG1("(~D*~(C*B))"),
    .INIT_LUTF0(16'b0000000000111111),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000000000111111),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9453|_al_u9541  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [42],\cu_ru/sepc [30]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9453_o,_al_u9541_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9454|ins_fetch/reg2_b42  (
    .a({_al_u9450_o,open_n72897}),
    .b({_al_u9451_o,_al_u9454_o}),
    .c({_al_u9452_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9453_o,_al_u9449_o}),
    .sr(rst_pad),
    .f({_al_u9454_o,open_n72911}),
    .q({open_n72915,addr_if[42]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9457|_al_u9469  (
    .b({\cu_ru/tvec [7],\cu_ru/tvec [42]}),
    .c({\cu_ru/n43 [3],\cu_ru/n43 [38]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .f({_al_u9457_o,_al_u9469_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000111000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9458|ins_fetch/reg2_b5  (
    .a({_al_u9457_o,_al_u9456_o}),
    .b({_al_u6055_o,_al_u9458_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[5],_al_u9459_o}),
    .sr(rst_pad),
    .f({_al_u9458_o,open_n72955}),
    .q({open_n72959,addr_if[5]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001010110111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9459|biu/bus_unit/mmu/reg2_b17  (
    .a({\cu_ru/m_s_status/n2 ,open_n72960}),
    .b({_al_u2844_o,open_n72961}),
    .c({\cu_ru/sepc [5],_al_u3159_o}),
    .clk(clk_pad),
    .d({\cu_ru/mepc [5],_al_u3158_o}),
    .sr(rst_pad),
    .f({_al_u9459_o,open_n72975}),
    .q({open_n72979,\biu/paddress [81]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b0000000100001011),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b0000000100001011),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9462|_al_u9606  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [43],\cu_ru/tvec [23]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [39],\cu_ru/n43 [19]}),
    .f({_al_u9462_o,_al_u9606_o}));
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9464|biu/bus_unit/mmu/reg2_b53  (
    .c({\cu_ru/mepc [41],_al_u3050_o}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,_al_u3049_o}),
    .sr(rst_pad),
    .f({_al_u9464_o,open_n73021}),
    .q({open_n73025,\biu/paddress [117]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9465|cu_ru/m_s_scratch/reg0_b41  (
    .b({_al_u2844_o,\cu_ru/sepc [41]}),
    .c({\cu_ru/sepc [41],data_csr[41]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n73038,data_csr[41]}),
    .sr(rst_pad),
    .f({_al_u9465_o,_al_u5465_o}),
    .q({open_n73042,\cu_ru/mscratch [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9466|ins_fetch/reg2_b41  (
    .a({_al_u9462_o,open_n73043}),
    .b({_al_u9463_o,_al_u9466_o}),
    .c({_al_u9464_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9465_o,_al_u9461_o}),
    .sr(rst_pad),
    .f({_al_u9466_o,open_n73057}),
    .q({open_n73061,addr_if[41]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9470|ins_fetch/reg2_b40  (
    .a({_al_u9469_o,_al_u9468_o}),
    .b({_al_u6055_o,_al_u9470_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[40],_al_u9471_o}),
    .sr(rst_pad),
    .f({_al_u9470_o,open_n73079}),
    .q({open_n73083,addr_if[40]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9471|cu_ru/m_s_scratch/reg0_b40  (
    .a({\cu_ru/m_s_status/n2 ,open_n73084}),
    .b({_al_u2844_o,\cu_ru/sepc [40]}),
    .c({\cu_ru/sepc [40],data_csr[40]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [40],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n73088,data_csr[40]}),
    .sr(rst_pad),
    .f({_al_u9471_o,_al_u5469_o}),
    .q({open_n73103,\cu_ru/mscratch [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9474|_al_u6022  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [41],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [41]}),
    .d({\cu_ru/n43 [37],\cu_ru/mtvec [41]}),
    .f({_al_u9474_o,\cu_ru/tvec [41]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9476|_al_u9575  (
    .c({\cu_ru/mepc [39],\cu_ru/mepc [25]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9476_o,_al_u9575_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9477|cu_ru/m_s_scratch/reg0_b39  (
    .b({_al_u2844_o,\cu_ru/sepc [39]}),
    .c({\cu_ru/sepc [39],data_csr[39]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n73161,data_csr[39]}),
    .sr(rst_pad),
    .f({_al_u9477_o,_al_u5477_o}),
    .q({open_n73176,\cu_ru/mscratch [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9478|ins_fetch/reg2_b39  (
    .a({_al_u9474_o,open_n73177}),
    .b({_al_u9475_o,_al_u9478_o}),
    .c({_al_u9476_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9477_o,_al_u9473_o}),
    .sr(rst_pad),
    .f({_al_u9478_o,open_n73195}),
    .q({open_n73199,addr_if[39]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b1110110010100000),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9481|_al_u6023  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [40],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [40]}),
    .d({\cu_ru/n43 [36],\cu_ru/mtvec [40]}),
    .f({_al_u9481_o,\cu_ru/tvec [40]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9483|_al_u9568  (
    .c({\cu_ru/mepc [38],\cu_ru/mepc [26]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9483_o,_al_u9568_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u9484|_al_u9522  (
    .b({_al_u2844_o,_al_u2844_o}),
    .c({\cu_ru/sepc [38],\cu_ru/sepc [32]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9484_o,_al_u9522_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9485|ins_fetch/reg2_b38  (
    .a({_al_u9481_o,open_n73270}),
    .b({_al_u9482_o,_al_u9485_o}),
    .c({_al_u9483_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9484_o,_al_u9480_o}),
    .sr(rst_pad),
    .f({_al_u9485_o,open_n73284}),
    .q({open_n73288,addr_if[38]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b0000000100001011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9488|_al_u9599  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [39],\cu_ru/tvec [5]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [35],\cu_ru/n43 [1]}),
    .f({_al_u9488_o,_al_u9599_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9490|_al_u9561  (
    .c({\cu_ru/mepc [37],\cu_ru/mepc [27]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9490_o,_al_u9561_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9492|ins_fetch/reg2_b37  (
    .a({_al_u9488_o,open_n73333}),
    .b({_al_u9489_o,_al_u9492_o}),
    .c({_al_u9490_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9491_o,_al_u9487_o}),
    .sr(rst_pad),
    .f({_al_u9492_o,open_n73347}),
    .q({open_n73351,addr_if[37]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9495|_al_u6026  (
    .a({open_n73352,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [38],\cu_ru/trap_target_m }),
    .c({\cu_ru/n43 [34],\cu_ru/stvec [38]}),
    .d({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mtvec [38]}),
    .f({_al_u9495_o,\cu_ru/tvec [38]}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9496|ins_fetch/reg2_b36  (
    .a({_al_u9495_o,_al_u9494_o}),
    .b({_al_u6055_o,_al_u9496_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[36],_al_u9497_o}),
    .sr(rst_pad),
    .f({_al_u9496_o,open_n73394}),
    .q({open_n73398,addr_if[36]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("~(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b1110110010100000),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b1110110010100000),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9500|_al_u6027  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [37],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [37]}),
    .d({\cu_ru/n43 [33],\cu_ru/mtvec [37]}),
    .f({_al_u9500_o,\cu_ru/tvec [37]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9502|_al_u7221  (
    .a({open_n73423,\cu_ru/read_mtvec_sel_lutinv }),
    .b({open_n73424,\cu_ru/read_mepc_sel_lutinv }),
    .c({\cu_ru/mepc [35],\cu_ru/mepc [35]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/mtvec [35]}),
    .f({_al_u9502_o,_al_u7221_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9503|cu_ru/m_s_scratch/reg0_b35  (
    .b({_al_u2844_o,\cu_ru/sepc [35]}),
    .c({\cu_ru/sepc [35],data_csr[35]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n73450,data_csr[35]}),
    .sr(rst_pad),
    .f({_al_u9503_o,_al_u5493_o}),
    .q({open_n73465,\cu_ru/mscratch [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9504|ins_fetch/reg2_b35  (
    .a({_al_u9500_o,open_n73466}),
    .b({_al_u9501_o,_al_u9504_o}),
    .c({_al_u9502_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9503_o,_al_u9499_o}),
    .sr(rst_pad),
    .f({_al_u9504_o,open_n73484}),
    .q({open_n73488,addr_if[35]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b0000000100001011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9507|_al_u9592  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [36],\cu_ru/tvec [24]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [32],\cu_ru/n43 [20]}),
    .f({_al_u9507_o,_al_u9592_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9509|_al_u9547  (
    .c({\cu_ru/mepc [34],\cu_ru/mepc [29]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_status/n2 }),
    .f({_al_u9509_o,_al_u9547_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9510|cu_ru/m_s_epc/reg0_b34  (
    .b({_al_u2844_o,_al_u5157_o}),
    .c({\cu_ru/sepc [34],_al_u5497_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/n2 [34]}),
    .sr(rst_pad),
    .f({_al_u9510_o,open_n73551}),
    .q({open_n73555,\cu_ru/sepc [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9511|ins_fetch/reg2_b34  (
    .a({_al_u9507_o,open_n73556}),
    .b({_al_u9508_o,_al_u9511_o}),
    .c({_al_u9509_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9510_o,_al_u9506_o}),
    .sr(rst_pad),
    .f({_al_u9511_o,open_n73574}),
    .q({open_n73578,addr_if[34]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9515|ins_fetch/reg2_b33  (
    .a({_al_u9514_o,_al_u9513_o}),
    .b({_al_u6055_o,_al_u9515_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[33],_al_u9516_o}),
    .sr(rst_pad),
    .f({_al_u9515_o,open_n73596}),
    .q({open_n73600,addr_if[33]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b1110110010100000),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9519|_al_u6030  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [34],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [34]}),
    .d({\cu_ru/n43 [30],\cu_ru/mtvec [34]}),
    .f({_al_u9519_o,\cu_ru/tvec [34]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9521|_al_u7419  (
    .a({open_n73621,\cu_ru/read_time_sel_lutinv }),
    .b({open_n73622,\cu_ru/read_mepc_sel_lutinv }),
    .c({\cu_ru/mepc [32],mtime_pad[32]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/mepc [32]}),
    .f({_al_u9521_o,_al_u7419_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9523|ins_fetch/reg2_b32  (
    .a({_al_u9519_o,open_n73643}),
    .b({_al_u9520_o,_al_u9523_o}),
    .c({_al_u9521_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9522_o,_al_u9518_o}),
    .sr(rst_pad),
    .f({_al_u9523_o,open_n73661}),
    .q({open_n73665,addr_if[32]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9527|ins_fetch/reg2_b4  (
    .a({_al_u9526_o,_al_u9525_o}),
    .b({_al_u6055_o,_al_u9527_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[4],_al_u9528_o}),
    .sr(rst_pad),
    .f({_al_u9527_o,open_n73683}),
    .q({open_n73687,addr_if[4]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0001010110111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9528|cu_ru/m_s_scratch/reg0_b4  (
    .a({\cu_ru/m_s_status/n2 ,open_n73688}),
    .b({_al_u2844_o,\cu_ru/sepc [4]}),
    .c({\cu_ru/sepc [4],data_csr[4]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [4],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n73699,data_csr[4]}),
    .sr(rst_pad),
    .f({_al_u9528_o,_al_u5473_o}),
    .q({open_n73703,\cu_ru/mscratch [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b0000000100001011),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b0000000100001011),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9531|_al_u9580  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [33],\cu_ru/tvec [26]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [29],\cu_ru/n43 [22]}),
    .f({_al_u9531_o,_al_u9580_o}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9534|cu_ru/m_s_scratch/reg0_b31  (
    .b({_al_u2844_o,\cu_ru/sepc [31]}),
    .c({\cu_ru/sepc [31],data_csr[31]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n73733,data_csr[31]}),
    .sr(rst_pad),
    .f({_al_u9534_o,_al_u5509_o}),
    .q({open_n73748,\cu_ru/mscratch [31]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9535|ins_fetch/reg2_b31  (
    .a({_al_u9531_o,open_n73749}),
    .b({_al_u9532_o,_al_u9535_o}),
    .c({_al_u9533_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9534_o,_al_u9530_o}),
    .sr(rst_pad),
    .f({_al_u9535_o,open_n73767}),
    .q({open_n73771,addr_if[31]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTF1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUTG1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUTF0(16'b0000000100001011),
    .INIT_LUTF1(16'b0000000100001011),
    .INIT_LUTG0(16'b0000000100001011),
    .INIT_LUTG1(16'b0000000100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9538|_al_u9573  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [32],\cu_ru/tvec [27]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [28],\cu_ru/n43 [23]}),
    .f({_al_u9538_o,_al_u9573_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9540|_al_u7433  (
    .a({open_n73796,\cu_ru/read_mepc_sel_lutinv }),
    .b({open_n73797,\cu_ru/read_stvec_sel_lutinv }),
    .c({\cu_ru/mepc [30],\cu_ru/mepc [30]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/stvec [30]}),
    .f({_al_u9540_o,_al_u7433_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9542|ins_fetch/reg2_b30  (
    .a({_al_u9538_o,open_n73822}),
    .b({_al_u9539_o,_al_u9542_o}),
    .c({_al_u9540_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9541_o,_al_u9537_o}),
    .sr(rst_pad),
    .f({_al_u9542_o,open_n73836}),
    .q({open_n73840,addr_if[30]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*B)*~(C*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b1110110010100000),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9545|_al_u6033  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/m_s_status/u14_sel_is_2_o }),
    .b({\cu_ru/tvec [31],\cu_ru/trap_target_m }),
    .c({_al_u6055_o,\cu_ru/stvec [31]}),
    .d({\cu_ru/n43 [27],\cu_ru/mtvec [31]}),
    .f({_al_u9545_o,\cu_ru/tvec [31]}));
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9548|cu_ru/m_s_scratch/reg0_b29  (
    .b({_al_u2844_o,\cu_ru/sepc [29]}),
    .c({\cu_ru/sepc [29],data_csr[29]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n73873,data_csr[29]}),
    .sr(rst_pad),
    .f({_al_u9548_o,_al_u5521_o}),
    .q({open_n73877,\cu_ru/mscratch [29]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9549|ins_fetch/reg2_b29  (
    .a({_al_u9545_o,open_n73878}),
    .b({_al_u9546_o,_al_u9549_o}),
    .c({_al_u9547_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9548_o,_al_u9544_o}),
    .sr(rst_pad),
    .f({_al_u9549_o,open_n73892}),
    .q({open_n73896,addr_if[29]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT_LUT0(16'b0000000100001011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"))
    \_al_u9552|_al_u9566  (
    .a({\cu_ru/mux34_b0_sel_is_2_o ,\cu_ru/mux34_b0_sel_is_2_o }),
    .b({\cu_ru/tvec [30],\cu_ru/tvec [28]}),
    .c({_al_u6055_o,_al_u6055_o}),
    .d({\cu_ru/n43 [26],\cu_ru/n43 [24]}),
    .f({_al_u9552_o,_al_u9566_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(D*B)*~(C*A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0001001101011111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001001101011111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9554|_al_u7445  (
    .a({open_n73917,\cu_ru/read_time_sel_lutinv }),
    .b({open_n73918,\cu_ru/read_mepc_sel_lutinv }),
    .c({\cu_ru/mepc [28],mtime_pad[28]}),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/mepc [28]}),
    .f({_al_u9554_o,_al_u7445_o}));
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9556|ins_fetch/reg2_b28  (
    .a({_al_u9552_o,open_n73943}),
    .b({_al_u9553_o,_al_u9556_o}),
    .c({_al_u9554_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9555_o,_al_u9551_o}),
    .sr(rst_pad),
    .f({_al_u9556_o,open_n73957}),
    .q({open_n73961,addr_if[28]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9562|cu_ru/m_s_scratch/reg0_b27  (
    .b({_al_u2844_o,\cu_ru/sepc [27]}),
    .c({\cu_ru/sepc [27],data_csr[27]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n73967,data_csr[27]}),
    .sr(rst_pad),
    .f({_al_u9562_o,_al_u5529_o}),
    .q({open_n73982,\cu_ru/mscratch [27]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9563|ins_fetch/reg2_b27  (
    .a({_al_u9559_o,open_n73983}),
    .b({_al_u9560_o,_al_u9563_o}),
    .c({_al_u9561_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9562_o,_al_u9558_o}),
    .sr(rst_pad),
    .f({_al_u9563_o,open_n73997}),
    .q({open_n74001,addr_if[27]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9570|ins_fetch/reg2_b26  (
    .a({_al_u9566_o,open_n74002}),
    .b({_al_u9567_o,_al_u9570_o}),
    .c({_al_u9568_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9569_o,_al_u9565_o}),
    .sr(rst_pad),
    .f({_al_u9570_o,open_n74020}),
    .q({open_n74024,addr_if[26]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9577|ins_fetch/reg2_b25  (
    .a({_al_u9573_o,open_n74025}),
    .b({_al_u9574_o,_al_u9577_o}),
    .c({_al_u9575_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9576_o,_al_u9572_o}),
    .sr(rst_pad),
    .f({_al_u9577_o,open_n74043}),
    .q({open_n74047,addr_if[25]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9583|cu_ru/m_s_scratch/reg0_b24  (
    .b({_al_u2844_o,\cu_ru/sepc [24]}),
    .c({\cu_ru/sepc [24],data_csr[24]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n74053,data_csr[24]}),
    .sr(rst_pad),
    .f({_al_u9583_o,_al_u5541_o}),
    .q({open_n74068,\cu_ru/mscratch [24]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9584|ins_fetch/reg2_b24  (
    .a({_al_u9580_o,open_n74069}),
    .b({_al_u9581_o,_al_u9584_o}),
    .c({_al_u9582_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9583_o,_al_u9579_o}),
    .sr(rst_pad),
    .f({_al_u9584_o,open_n74087}),
    .q({open_n74091,addr_if[24]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000111000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9588|ins_fetch/reg2_b23  (
    .a({_al_u9587_o,_al_u9586_o}),
    .b({_al_u6055_o,_al_u9588_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[23],_al_u9589_o}),
    .sr(rst_pad),
    .f({_al_u9588_o,open_n74105}),
    .q({open_n74109,addr_if[23]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9589|cu_ru/m_s_scratch/reg0_b23  (
    .a({\cu_ru/m_s_status/n2 ,open_n74110}),
    .b({_al_u2844_o,\cu_ru/sepc [23]}),
    .c({\cu_ru/sepc [23],data_csr[23]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/mepc [23],\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n74114,data_csr[23]}),
    .sr(rst_pad),
    .f({_al_u9589_o,_al_u5545_o}),
    .q({open_n74129,\cu_ru/mscratch [23]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9595|cu_ru/m_s_scratch/reg0_b22  (
    .b({_al_u2844_o,\cu_ru/sepc [22]}),
    .c({\cu_ru/sepc [22],data_csr[22]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n74142,data_csr[22]}),
    .sr(rst_pad),
    .f({_al_u9595_o,_al_u5549_o}),
    .q({open_n74146,\cu_ru/mscratch [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9596|ins_fetch/reg2_b22  (
    .a({_al_u9592_o,open_n74147}),
    .b({_al_u9593_o,_al_u9596_o}),
    .c({_al_u9594_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9595_o,_al_u9591_o}),
    .sr(rst_pad),
    .f({_al_u9596_o,open_n74161}),
    .q({open_n74165,addr_if[22]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9603|ins_fetch/reg2_b3  (
    .a({_al_u9599_o,open_n74166}),
    .b({_al_u9600_o,_al_u9603_o}),
    .c({_al_u9601_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9602_o,_al_u9598_o}),
    .sr(rst_pad),
    .f({_al_u9603_o,open_n74180}),
    .q({open_n74184,addr_if[3]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9608|biu/bus_unit/mmu/reg2_b33  (
    .c({\cu_ru/mepc [21],_al_u3110_o}),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,_al_u3109_o}),
    .sr(rst_pad),
    .f({_al_u9608_o,open_n74202}),
    .q({open_n74206,\biu/paddress [97]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9609|cu_ru/m_s_scratch/reg0_b21  (
    .b({_al_u2844_o,\cu_ru/sepc [21]}),
    .c({\cu_ru/sepc [21],data_csr[21]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n74212,data_csr[21]}),
    .sr(rst_pad),
    .f({_al_u9609_o,_al_u5553_o}),
    .q({open_n74227,\cu_ru/mscratch [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9610|ins_fetch/reg2_b21  (
    .a({_al_u9606_o,open_n74228}),
    .b({_al_u9607_o,_al_u9610_o}),
    .c({_al_u9608_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9609_o,_al_u9605_o}),
    .sr(rst_pad),
    .f({_al_u9610_o,open_n74242}),
    .q({open_n74246,addr_if[21]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9617|ins_fetch/reg2_b20  (
    .a({_al_u9613_o,open_n74247}),
    .b({_al_u9614_o,_al_u9617_o}),
    .c({_al_u9615_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9616_o,_al_u9612_o}),
    .sr(rst_pad),
    .f({_al_u9617_o,open_n74265}),
    .q({open_n74269,addr_if[20]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000111000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9621|ins_fetch/reg2_b19  (
    .a({_al_u9620_o,_al_u9619_o}),
    .b({_al_u6055_o,_al_u9621_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[19],_al_u9622_o}),
    .sr(rst_pad),
    .f({_al_u9621_o,open_n74283}),
    .q({open_n74287,addr_if[19]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1100111100000011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9628|cu_ru/m_s_epc/reg0_b18  (
    .b({_al_u2844_o,_al_u5157_o}),
    .c({\cu_ru/sepc [18],_al_u5569_o}),
    .ce(\cu_ru/trap_target_m ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/n2 [18]}),
    .sr(rst_pad),
    .f({_al_u9628_o,open_n74306}),
    .q({open_n74310,\cu_ru/sepc [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9629|ins_fetch/reg2_b18  (
    .a({_al_u9625_o,open_n74311}),
    .b({_al_u9626_o,_al_u9629_o}),
    .c({_al_u9627_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9628_o,_al_u9624_o}),
    .sr(rst_pad),
    .f({_al_u9629_o,open_n74329}),
    .q({open_n74333,addr_if[18]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9636|ins_fetch/reg2_b17  (
    .a({_al_u9632_o,open_n74334}),
    .b({_al_u9633_o,_al_u9636_o}),
    .c({_al_u9634_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9635_o,_al_u9631_o}),
    .sr(rst_pad),
    .f({_al_u9636_o,open_n74352}),
    .q({open_n74356,addr_if[17]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9643|ins_fetch/reg2_b16  (
    .a({_al_u9639_o,open_n74357}),
    .b({_al_u9640_o,_al_u9643_o}),
    .c({_al_u9641_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9642_o,_al_u9638_o}),
    .sr(rst_pad),
    .f({_al_u9643_o,open_n74371}),
    .q({open_n74375,addr_if[16]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*C*~B))"),
    //.LUTF1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~A*~(D*C*~B))"),
    //.LUTG1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010101010101),
    .INIT_LUTF1(16'b0000111000000010),
    .INIT_LUTG0(16'b0100010101010101),
    .INIT_LUTG1(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9647|ins_fetch/reg2_b15  (
    .a({_al_u9646_o,_al_u9645_o}),
    .b({_al_u6055_o,_al_u9647_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[15],_al_u9648_o}),
    .sr(rst_pad),
    .f({_al_u9647_o,open_n74393}),
    .q({open_n74397,addr_if[15]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0001010110111111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9648|biu/bus_unit/mmu/reg2_b27  (
    .a({\cu_ru/m_s_status/n2 ,open_n74398}),
    .b({_al_u2844_o,open_n74399}),
    .c({\cu_ru/sepc [15],_al_u3128_o}),
    .clk(clk_pad),
    .d({\cu_ru/mepc [15],_al_u3127_o}),
    .sr(rst_pad),
    .f({_al_u9648_o,open_n74417}),
    .q({open_n74421,\biu/paddress [91]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9653|cu_ru/m_cycle_event/reg0_b14  (
    .a({open_n74422,_al_u6763_o}),
    .b({open_n74423,\cu_ru/read_mepc_sel_lutinv }),
    .c({\cu_ru/mepc [14],\cu_ru/minstret [14]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/mepc [14]}),
    .mi({open_n74427,\cu_ru/m_cycle_event/n4 [14]}),
    .sr(rst_pad),
    .f({_al_u9653_o,_al_u7467_o}),
    .q({open_n74442,\cu_ru/minstret [14]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9655|ins_fetch/reg2_b14  (
    .a({_al_u9651_o,open_n74443}),
    .b({_al_u9652_o,_al_u9655_o}),
    .c({_al_u9653_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9654_o,_al_u9650_o}),
    .sr(rst_pad),
    .f({_al_u9655_o,open_n74457}),
    .q({open_n74461,addr_if[14]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9661|cu_ru/m_s_scratch/reg1_b13  (
    .b({_al_u2844_o,\cu_ru/sepc [13]}),
    .c({\cu_ru/sepc [13],data_csr[13]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n74467,data_csr[13]}),
    .sr(rst_pad),
    .f({_al_u9661_o,_al_u5589_o}),
    .q({open_n74482,\cu_ru/sscratch [13]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~C*~(D*~(B*~A)))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~C*~(D*~(B*~A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000010000001111),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000010000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9662|ins_fetch/reg2_b13  (
    .a({_al_u9658_o,open_n74483}),
    .b({_al_u9659_o,_al_u9662_o}),
    .c({_al_u9660_o,pip_flush}),
    .clk(clk_pad),
    .d({_al_u9661_o,_al_u9657_o}),
    .sr(rst_pad),
    .f({_al_u9662_o,open_n74501}),
    .q({open_n74505,addr_if[13]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(D*C*~B))"),
    //.LUT1("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100010101010101),
    .INIT_LUT1(16'b0000111000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9666|ins_fetch/reg2_b12  (
    .a({_al_u9665_o,_al_u9664_o}),
    .b({_al_u6055_o,_al_u9666_o}),
    .c({_al_u2842_o,pip_flush}),
    .clk(clk_pad),
    .d({new_pc[12],_al_u9667_o}),
    .sr(rst_pad),
    .f({_al_u9666_o,open_n74519}),
    .q({open_n74523,addr_if[12]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/IF/ins_fetch.v(83)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b0000001000010011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b0000001000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9669|ins_fetch/reg2_b2  (
    .a({\ins_fetch/n27 ,open_n74524}),
    .b({pip_flush,_al_u9674_o}),
    .c({\ins_fetch/n1 [0],pip_flush}),
    .clk(clk_pad),
    .d({addr_if[2],_al_u9669_o}),
    .sr(rst_pad),
    .f({_al_u9669_o,open_n74542}),
    .q({open_n74546,addr_if[2]}));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~(C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9673|cu_ru/medeleg_exc_ctrl/dii_reg  (
    .b({_al_u2844_o,\cu_ru/sepc [2]}),
    .c({\cu_ru/sepc [2],data_csr[2]}),
    .ce(\cu_ru/medeleg_exc_ctrl/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_status/n2 ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .mi({open_n74559,data_csr[2]}),
    .sr(rst_pad),
    .f({_al_u9673_o,_al_u5561_o}),
    .q({open_n74563,\cu_ru/medeleg [2]}));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(~C*~(D*~(B*~A)))"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0000010000001111),
    .MODE("LOGIC"))
    \_al_u9674|_al_u9671  (
    .a({_al_u9670_o,open_n74564}),
    .b({_al_u9671_o,_al_u2844_o}),
    .c({_al_u9672_o,new_pc[2]}),
    .d({_al_u9673_o,_al_u6055_o}),
    .f({_al_u9674_o,_al_u9671_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~C*A))"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~B*~(D*~C*A))"),
    //.LUTG1("(C*~B*D)"),
    .INIT_LUTF0(16'b0011000100110011),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b0011000100110011),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9676|_al_u9284  (
    .a({open_n74585,_al_u9204_o}),
    .b({_al_u9264_o,_al_u9283_o}),
    .c({\biu/cache_ctrl_logic/n55_lutinv ,_al_u9264_o}),
    .d({_al_u9204_o,\biu/cache_ctrl_logic/n55_lutinv }),
    .f({_al_u9676_o,_al_u9284_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~B*~(D*~C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011001000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9678|biu/cache_ctrl_logic/reg5_b63  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({_al_u7151_o,\biu/cache_ctrl_logic/l1i_pte [63]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/statu [0],\biu/cache_ctrl_logic/l1d_pte [63]}),
    .mi({open_n74620,\biu/cache_ctrl_logic/pte_temp [63]}),
    .sr(rst_pad),
    .f({_al_u9678_o,_al_u5676_o}),
    .q({open_n74624,\biu/cache_ctrl_logic/l1d_pte [63]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~B*~(C*~(D*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0010001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u9679|biu/cache_ctrl_logic/reg5_b38  (
    .a({\biu/cache_ctrl_logic/n100 [4],_al_u3947_o}),
    .b({_al_u9677_o,_al_u3950_o}),
    .c({_al_u9678_o,\biu/cache_ctrl_logic/l1i_pte [38]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u3947_o,\biu/cache_ctrl_logic/l1d_pte [38]}),
    .mi({open_n74635,\biu/cache_ctrl_logic/pte_temp [38]}),
    .sr(rst_pad),
    .f({_al_u9679_o,_al_u5776_o}),
    .q({open_n74639,\biu/cache_ctrl_logic/l1d_pte [38]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(~C*~(B*~D))"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(~C*~(B*~D))"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b0000111100000011),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b0000111100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9680|_al_u9708  (
    .b({_al_u4399_o,\biu/cache_ctrl_logic/n75_lutinv }),
    .c({\biu/cache_ctrl_logic/n204_lutinv ,\biu/cache_ctrl_logic/n204_lutinv }),
    .d({\biu/cache_ctrl_logic/n100 [4],\biu/cache_ctrl_logic/n100 [4]}),
    .f({_al_u9680_o,_al_u9708_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~(~D*~B*~A))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000011100000),
    .MODE("LOGIC"))
    \_al_u9682|_al_u9681  (
    .a({_al_u9272_o,open_n74666}),
    .b({_al_u9679_o,open_n74667}),
    .c({_al_u9680_o,\biu/cache_ctrl_logic/n97_lutinv }),
    .d({_al_u9681_o,_al_u7149_o}),
    .f({_al_u9682_o,_al_u9681_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(~D*~C)))"),
    //.LUT1("(C*A*~(D*B))"),
    .INIT_LUT0(16'b0100010001001100),
    .INIT_LUT1(16'b0010000010100000),
    .MODE("LOGIC"))
    \_al_u9685|_al_u7158  (
    .a({\biu/cache_ctrl_logic/n83 [0],_al_u7157_o}),
    .b({_al_u7157_o,\biu/cache_ctrl_logic/n75_lutinv }),
    .c({\biu/cache_ctrl_logic/n75_lutinv ,read}),
    .d({write,write}),
    .f({_al_u9685_o,_al_u7158_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*B))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000000111111),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u9686|_al_u9683  (
    .b({open_n74710,\biu/cache_ctrl_logic/n100 [4]}),
    .c({write,_al_u4834_o}),
    .d({_al_u7149_o,_al_u9682_o}),
    .f({_al_u9686_o,_al_u9683_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D*~A)))"),
    //.LUT1("(~B*~(~D*C*~A))"),
    .INIT_LUT0(16'b0000011100000011),
    .INIT_LUT1(16'b0011001100100011),
    .MODE("LOGIC"))
    \_al_u9688|_al_u9687  (
    .a({_al_u9683_o,_al_u9686_o}),
    .b({_al_u9685_o,\biu/cache_ctrl_logic/l1d_wr_sel_lutinv }),
    .c({_al_u9687_o,\biu/cache_ctrl_logic/n75_lutinv }),
    .d({_al_u2848_o,\biu/cache_ctrl_logic/n100 [4]}),
    .f({_al_u9688_o,_al_u9687_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9689|_al_u9684  (
    .b({open_n74753,read}),
    .c({_al_u7191_o,\biu/cache_ctrl_logic/n100 [4]}),
    .d({_al_u7190_o,_al_u7190_o}),
    .f({_al_u9689_o,\biu/cache_ctrl_logic/n83 [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1101000011010101),
    .MODE("LOGIC"))
    \_al_u9690|_al_u3414  (
    .a({_al_u9689_o,open_n74778}),
    .b({\biu/cache_ctrl_logic/n100 [4],open_n74779}),
    .c({_al_u7149_o,_al_u2886_o}),
    .d({_al_u2886_o,\biu/cache_ctrl_logic/n100 [4]}),
    .f({_al_u9690_o,\biu/cache_ctrl_logic/n135 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u9691|_al_u9285  (
    .c({_al_u7162_o,\biu/cache_ctrl_logic/l1d_pte [7]}),
    .d({_al_u9690_o,_al_u7193_o}),
    .f({_al_u9691_o,_al_u9285_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~D*~C*~(B*A))"),
    .INIT_LUT0(16'b1100110100001101),
    .INIT_LUT1(16'b0000000000000111),
    .MODE("LOGIC"))
    \_al_u9692|_al_u9713  (
    .a({_al_u9688_o,_al_u9712_o}),
    .b({_al_u9691_o,_al_u9286_o}),
    .c({_al_u9286_o,_al_u7193_o}),
    .d({_al_u7193_o,\biu/cache_ctrl_logic/l1d_pte [7]}),
    .f({_al_u9692_o,_al_u9713_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*B*A))"),
    //.LUT1("(~A*~(D*C*B))"),
    .INIT_LUT0(16'b0000011100001111),
    .INIT_LUT1(16'b0001010101010101),
    .MODE("LOGIC"))
    \_al_u9693|_al_u3211  (
    .a({_al_u9283_o,\exu/c_fence_lutinv }),
    .b({\exu/c_fence_lutinv ,\biu/cache_ctrl_logic/n55_lutinv }),
    .c({\biu/cache_ctrl_logic/n55_lutinv ,rst_pad}),
    .d({cache_flush,cache_flush}),
    .f({_al_u9693_o,\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~D*~(C*~B)))"),
    //.LUT1("(~D*~(C*B))"),
    .INIT_LUT0(16'b1010101000100000),
    .INIT_LUT1(16'b0000000000111111),
    .MODE("LOGIC"))
    \_al_u9695|_al_u9696  (
    .a({open_n74864,_al_u9271_o}),
    .b({_al_u9274_o,_al_u9272_o}),
    .c({\biu/cache_ctrl_logic/statu [2],_al_u9695_o}),
    .d({_al_u9273_o,_al_u4399_o}),
    .f({_al_u9695_o,_al_u9696_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*~(D*~A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*B*~(D*~A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1000000011000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1000000011000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9697|_al_u9278  (
    .a({open_n74885,\biu/cache_ctrl_logic/n100 [4]}),
    .b({open_n74886,_al_u7149_o}),
    .c({\biu/cache_ctrl_logic/n100 [4],_al_u4834_o}),
    .d({_al_u9278_o,1'b0}),
    .f({_al_u9697_o,_al_u9278_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~B*~(~C*~D))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0011001100110000),
    .MODE("LOGIC"))
    \_al_u9699|_al_u9698  (
    .b({_al_u9697_o,open_n74913}),
    .c({_al_u9698_o,_al_u3224_o}),
    .d({_al_u9696_o,_al_u7149_o}),
    .f({_al_u9699_o,_al_u9698_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(D*~B*~A))"),
    //.LUT1("(~D*~B*~(C*A))"),
    .INIT_LUT0(16'b0000111000001111),
    .INIT_LUT1(16'b0000000000010011),
    .MODE("LOGIC"))
    \_al_u9700|_al_u9281  (
    .a({_al_u9699_o,_al_u9279_o}),
    .b({_al_u9280_o,\biu/cache_ctrl_logic/n149 }),
    .c({_al_u7159_o,_al_u9280_o}),
    .d({_al_u2886_o,_al_u7159_o}),
    .f({_al_u9700_o,_al_u9281_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~D*~(~C*~A)))"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1100110000000100),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u9701|_al_u9702  (
    .a({open_n74954,_al_u9700_o}),
    .b({open_n74955,_al_u7192_o}),
    .c({_al_u2885_o,_al_u9701_o}),
    .d({_al_u7163_o,\biu/bus_unit/mmu/n19_lutinv }),
    .f({_al_u9701_o,_al_u9702_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9704|_al_u9705  (
    .b({open_n74978,_al_u9704_o}),
    .c({\biu/cache_ctrl_logic/statu [1],_al_u3947_o}),
    .d({_al_u7151_o,_al_u7149_o}),
    .f({_al_u9704_o,_al_u9705_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(C*~B*~(~D*~A))"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(C*~B*~(~D*~A))"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b0011000000100000),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b0011000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u9709|_al_u9706  (
    .a({_al_u9706_o,open_n75003}),
    .b({_al_u9707_o,_al_u9705_o}),
    .c({_al_u9708_o,_al_u3950_o}),
    .d({_al_u9681_o,\biu/cache_ctrl_logic/n100 [4]}),
    .f({_al_u9709_o,_al_u9706_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~B*~(~C*~A)))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000011001101),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u9710|_al_u9711  (
    .a({open_n75028,_al_u9709_o}),
    .b({open_n75029,_al_u9710_o}),
    .c({_al_u2885_o,_al_u7158_o}),
    .d({_al_u7163_o,\biu/bus_unit/mmu/n19_lutinv }),
    .f({_al_u9710_o,_al_u9711_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~C*~D))"),
    //.LUT1("(~B*~(~D*~C*~A))"),
    .INIT_LUT0(16'b1100110011000000),
    .INIT_LUT1(16'b0011001100110010),
    .MODE("LOGIC"))
    \_al_u9712|_al_u5116  (
    .a({_al_u9711_o,open_n75050}),
    .b({_al_u7162_o,_al_u5115_o}),
    .c({_al_u9689_o,_al_u3222_o}),
    .d({_al_u2848_o,_al_u4208_o}),
    .f({_al_u9712_o,_al_u5116_o}));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*A*~(~D*~B))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101111101111111),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u9715|biu/cache_ctrl_logic/reg8_b2  (
    .a({open_n75071,_al_u9284_o}),
    .b({_al_u9287_o,_al_u9702_o}),
    .c({\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ,_al_u9287_o}),
    .clk(clk_pad),
    .d({_al_u9284_o,_al_u7193_o}),
    .sr(\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ),
    .f({\biu/cache_ctrl_logic/mux44_b4_sel_is_2_o ,open_n75085}),
    .q({open_n75089,\biu/cache_ctrl_logic/statu [2]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add0/u0|biu/bus_unit/add0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add0/u0|biu/bus_unit/add0/ucin  (
    .a({\biu/bus_unit/addr_counter [0],1'b0}),
    .b({1'b1,open_n75090}),
    .f({\biu/bus_unit/n39 [0],open_n75110}),
    .fco(\biu/bus_unit/add0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add0/u0|biu/bus_unit/add0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add0/u2|biu/bus_unit/add0/u1  (
    .a(\biu/bus_unit/addr_counter [2:1]),
    .b(2'b00),
    .fci(\biu/bus_unit/add0/c1 ),
    .f(\biu/bus_unit/n39 [2:1]),
    .fco(\biu/bus_unit/add0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add0/u0|biu/bus_unit/add0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add0/u4|biu/bus_unit/add0/u3  (
    .a(\biu/bus_unit/addr_counter [4:3]),
    .b(2'b00),
    .fci(\biu/bus_unit/add0/c3 ),
    .f(\biu/bus_unit/n39 [4:3]),
    .fco(\biu/bus_unit/add0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add0/u0|biu/bus_unit/add0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add0/u6|biu/bus_unit/add0/u5  (
    .a(\biu/bus_unit/addr_counter [6:5]),
    .b(2'b00),
    .fci(\biu/bus_unit/add0/c5 ),
    .f(\biu/bus_unit/n39 [6:5]),
    .fco(\biu/bus_unit/add0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add0/u0|biu/bus_unit/add0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add0/u8|biu/bus_unit/add0/u7  (
    .a(\biu/bus_unit/addr_counter [8:7]),
    .b(2'b00),
    .fci(\biu/bus_unit/add0/c7 ),
    .f(\biu/bus_unit/n39 [8:7]));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin  (
    .a({\biu/bus_unit/addr_counter [0],1'b0}),
    .b({\biu/maddress [3],open_n75204}),
    .f({\biu/bus_unit/n49 [0],open_n75224}),
    .fco(\biu/bus_unit/add1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u10|biu/bus_unit/add1/u9  (
    .a(2'b00),
    .b(\biu/maddress [13:12]),
    .fci(\biu/bus_unit/add1/c9 ),
    .f(\biu/bus_unit/n49 [10:9]),
    .fco(\biu/bus_unit/add1/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u12|biu/bus_unit/add1/u11  (
    .a(2'b00),
    .b(\biu/maddress [15:14]),
    .fci(\biu/bus_unit/add1/c11 ),
    .f(\biu/bus_unit/n49 [12:11]),
    .fco(\biu/bus_unit/add1/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u14|biu/bus_unit/add1/u13  (
    .a(2'b00),
    .b(\biu/maddress [17:16]),
    .fci(\biu/bus_unit/add1/c13 ),
    .f(\biu/bus_unit/n49 [14:13]),
    .fco(\biu/bus_unit/add1/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u16|biu/bus_unit/add1/u15  (
    .a(2'b00),
    .b(\biu/maddress [19:18]),
    .fci(\biu/bus_unit/add1/c15 ),
    .f(\biu/bus_unit/n49 [16:15]),
    .fco(\biu/bus_unit/add1/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u18|biu/bus_unit/add1/u17  (
    .a(2'b00),
    .b(\biu/maddress [21:20]),
    .fci(\biu/bus_unit/add1/c17 ),
    .f(\biu/bus_unit/n49 [18:17]),
    .fco(\biu/bus_unit/add1/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u20|biu/bus_unit/add1/u19  (
    .a(2'b00),
    .b(\biu/maddress [23:22]),
    .fci(\biu/bus_unit/add1/c19 ),
    .f(\biu/bus_unit/n49 [20:19]),
    .fco(\biu/bus_unit/add1/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u22|biu/bus_unit/add1/u21  (
    .a(2'b00),
    .b(\biu/maddress [25:24]),
    .fci(\biu/bus_unit/add1/c21 ),
    .f(\biu/bus_unit/n49 [22:21]),
    .fco(\biu/bus_unit/add1/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u24|biu/bus_unit/add1/u23  (
    .a(2'b00),
    .b(\biu/maddress [27:26]),
    .fci(\biu/bus_unit/add1/c23 ),
    .f(\biu/bus_unit/n49 [24:23]),
    .fco(\biu/bus_unit/add1/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u26|biu/bus_unit/add1/u25  (
    .a(2'b00),
    .b(\biu/maddress [29:28]),
    .fci(\biu/bus_unit/add1/c25 ),
    .f(\biu/bus_unit/n49 [26:25]),
    .fco(\biu/bus_unit/add1/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u28|biu/bus_unit/add1/u27  (
    .a(2'b00),
    .b(\biu/maddress [31:30]),
    .fci(\biu/bus_unit/add1/c27 ),
    .f(\biu/bus_unit/n49 [28:27]),
    .fco(\biu/bus_unit/add1/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u2|biu/bus_unit/add1/u1  (
    .a(\biu/bus_unit/addr_counter [2:1]),
    .b(\biu/maddress [5:4]),
    .fci(\biu/bus_unit/add1/c1 ),
    .f(\biu/bus_unit/n49 [2:1]),
    .fco(\biu/bus_unit/add1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u30|biu/bus_unit/add1/u29  (
    .a(2'b00),
    .b(\biu/maddress [33:32]),
    .fci(\biu/bus_unit/add1/c29 ),
    .f(\biu/bus_unit/n49 [30:29]),
    .fco(\biu/bus_unit/add1/c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u32|biu/bus_unit/add1/u31  (
    .a(2'b00),
    .b(\biu/maddress [35:34]),
    .fci(\biu/bus_unit/add1/c31 ),
    .f(\biu/bus_unit/n49 [32:31]),
    .fco(\biu/bus_unit/add1/c33 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y8Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u34|biu/bus_unit/add1/u33  (
    .a(2'b00),
    .b(\biu/maddress [37:36]),
    .fci(\biu/bus_unit/add1/c33 ),
    .f(\biu/bus_unit/n49 [34:33]),
    .fco(\biu/bus_unit/add1/c35 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y9Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u36|biu/bus_unit/add1/u35  (
    .a(2'b00),
    .b(\biu/maddress [39:38]),
    .fci(\biu/bus_unit/add1/c35 ),
    .f(\biu/bus_unit/n49 [36:35]),
    .fco(\biu/bus_unit/add1/c37 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y9Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u38|biu/bus_unit/add1/u37  (
    .a(2'b00),
    .b(\biu/maddress [41:40]),
    .fci(\biu/bus_unit/add1/c37 ),
    .f(\biu/bus_unit/n49 [38:37]),
    .fco(\biu/bus_unit/add1/c39 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y10Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u40|biu/bus_unit/add1/u39  (
    .a(2'b00),
    .b(\biu/maddress [43:42]),
    .fci(\biu/bus_unit/add1/c39 ),
    .f(\biu/bus_unit/n49 [40:39]),
    .fco(\biu/bus_unit/add1/c41 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y10Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u42|biu/bus_unit/add1/u41  (
    .a(2'b00),
    .b(\biu/maddress [45:44]),
    .fci(\biu/bus_unit/add1/c41 ),
    .f(\biu/bus_unit/n49 [42:41]),
    .fco(\biu/bus_unit/add1/c43 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y11Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u44|biu/bus_unit/add1/u43  (
    .a(2'b00),
    .b(\biu/maddress [47:46]),
    .fci(\biu/bus_unit/add1/c43 ),
    .f(\biu/bus_unit/n49 [44:43]),
    .fco(\biu/bus_unit/add1/c45 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y11Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u46|biu/bus_unit/add1/u45  (
    .a(2'b00),
    .b(\biu/maddress [49:48]),
    .fci(\biu/bus_unit/add1/c45 ),
    .f(\biu/bus_unit/n49 [46:45]),
    .fco(\biu/bus_unit/add1/c47 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y12Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u48|biu/bus_unit/add1/u47  (
    .a(2'b00),
    .b(\biu/maddress [51:50]),
    .fci(\biu/bus_unit/add1/c47 ),
    .f(\biu/bus_unit/n49 [48:47]),
    .fco(\biu/bus_unit/add1/c49 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u4|biu/bus_unit/add1/u3  (
    .a(\biu/bus_unit/addr_counter [4:3]),
    .b(\biu/maddress [7:6]),
    .fci(\biu/bus_unit/add1/c3 ),
    .f(\biu/bus_unit/n49 [4:3]),
    .fco(\biu/bus_unit/add1/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y12Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u50|biu/bus_unit/add1/u49  (
    .a(2'b00),
    .b(\biu/maddress [53:52]),
    .fci(\biu/bus_unit/add1/c49 ),
    .f(\biu/bus_unit/n49 [50:49]),
    .fco(\biu/bus_unit/add1/c51 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y13Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u52|biu/bus_unit/add1/u51  (
    .a(2'b00),
    .b(\biu/maddress [55:54]),
    .fci(\biu/bus_unit/add1/c51 ),
    .f(\biu/bus_unit/n49 [52:51]),
    .fco(\biu/bus_unit/add1/c53 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y13Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u54|biu/bus_unit/add1/u53  (
    .a(2'b00),
    .b(\biu/maddress [57:56]),
    .fci(\biu/bus_unit/add1/c53 ),
    .f(\biu/bus_unit/n49 [54:53]),
    .fco(\biu/bus_unit/add1/c55 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y14Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u56|biu/bus_unit/add1/u55  (
    .a(2'b00),
    .b(\biu/maddress [59:58]),
    .fci(\biu/bus_unit/add1/c55 ),
    .f(\biu/bus_unit/n49 [56:55]),
    .fco(\biu/bus_unit/add1/c57 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y14Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u58|biu/bus_unit/add1/u57  (
    .a(2'b00),
    .b(\biu/maddress [61:60]),
    .fci(\biu/bus_unit/add1/c57 ),
    .f(\biu/bus_unit/n49 [58:57]),
    .fco(\biu/bus_unit/add1/c59 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y15Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u60|biu/bus_unit/add1/u59  (
    .a(2'b00),
    .b(\biu/maddress [63:62]),
    .fci(\biu/bus_unit/add1/c59 ),
    .f(\biu/bus_unit/n49 [60:59]));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u6|biu/bus_unit/add1/u5  (
    .a(\biu/bus_unit/addr_counter [6:5]),
    .b(\biu/maddress [9:8]),
    .fci(\biu/bus_unit/add1/c5 ),
    .f(\biu/bus_unit/n49 [6:5]),
    .fco(\biu/bus_unit/add1/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/add1/u0|biu/bus_unit/add1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \biu/bus_unit/add1/u8|biu/bus_unit/add1/u7  (
    .a(\biu/bus_unit/addr_counter [8:7]),
    .b(\biu/maddress [11:10]),
    .fci(\biu/bus_unit/add1/c7 ),
    .f(\biu/bus_unit/n49 [8:7]),
    .fco(\biu/bus_unit/add1/c9 ));
  // ../../RTL/CPU/BIU/mmu.v(166)
  // ../../RTL/CPU/BIU/mmu.v(166)
  EG_PHY_MSLICE #(
    //.LUT0("~(C@D)"),
    //.LUT1("(~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000001111),
    .INIT_LUT1(16'b0000000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/bus_unit/mmu/reg0_b0|biu/bus_unit/mmu/reg0_b1  (
    .c({open_n75894,\biu/bus_unit/mmu/i [1]}),
    .ce(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu/i [0],\biu/bus_unit/mmu/i [0]}),
    .sr(\biu/bus_unit/mmu/n58 ),
    .q({\biu/bus_unit/mmu/i [0],\biu/bus_unit/mmu/i [1]}));  // ../../RTL/CPU/BIU/mmu.v(166)
  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/bus_unit/mmu/reg2_b0|biu/bus_unit/mmu/reg2_b63  (
    .c({\biu/paddress [64],\biu/paddress [127]}),
    .clk(clk_pad),
    .d({_al_u3034_o,_al_u3034_o}),
    .sr(rst_pad),
    .q({\biu/paddress [64],\biu/paddress [127]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/bus_unit/mmu/reg2_b1|biu/bus_unit/mmu/reg2_b62  (
    .c({\biu/paddress [65],\biu/paddress [126]}),
    .clk(clk_pad),
    .d({_al_u3034_o,_al_u3034_o}),
    .sr(rst_pad),
    .q({\biu/paddress [65],\biu/paddress [126]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/bus_unit/mmu/reg2_b2|biu/bus_unit/mmu/reg2_b61  (
    .c({\biu/paddress [66],\biu/paddress [125]}),
    .clk(clk_pad),
    .d({_al_u3034_o,_al_u3034_o}),
    .sr(rst_pad),
    .q({\biu/paddress [66],\biu/paddress [125]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/bus_unit/mmu/reg2_b56|biu/bus_unit/mmu/reg2_b60  (
    .c({\biu/paddress [120],\biu/paddress [124]}),
    .clk(clk_pad),
    .d({_al_u3034_o,_al_u3034_o}),
    .sr(rst_pad),
    .q({\biu/paddress [120],\biu/paddress [124]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/mmu.v(200)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/bus_unit/mmu/reg2_b57|biu/bus_unit/mmu/reg2_b59  (
    .c({\biu/paddress [121],\biu/paddress [123]}),
    .clk(clk_pad),
    .d({_al_u3034_o,_al_u3034_o}),
    .sr(rst_pad),
    .q({\biu/paddress [121],\biu/paddress [123]}));  // ../../RTL/CPU/BIU/mmu.v(200)
  // ../../RTL/CPU/BIU/bus_unit.v(177)
  // ../../RTL/CPU/BIU/bus_unit.v(177)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("~(~C*~D)"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/bus_unit/reg0_b0|biu/bus_unit/reg0_b8  (
    .c({\biu/bus_unit/n39 [0],\biu/bus_unit/n39 [8]}),
    .ce(\biu/bus_unit/n39[0]_en ),
    .clk(clk_pad),
    .d({\biu/bus_unit/n15_lutinv ,\biu/bus_unit/n15_lutinv }),
    .sr(\biu/bus_unit/n37 ),
    .q({\biu/bus_unit/addr_counter [0],\biu/bus_unit/addr_counter [8]}));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  // ../../RTL/CPU/BIU/bus_unit.v(177)
  // ../../RTL/CPU/BIU/bus_unit.v(177)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/bus_unit/reg0_b1|biu/bus_unit/reg0_b7  (
    .c({\biu/bus_unit/n39 [1],\biu/bus_unit/n39 [7]}),
    .ce(\biu/bus_unit/n39[0]_en ),
    .clk(clk_pad),
    .d({\biu/bus_unit/n15_lutinv ,\biu/bus_unit/n15_lutinv }),
    .sr(\biu/bus_unit/n37 ),
    .q({\biu/bus_unit/addr_counter [1],\biu/bus_unit/addr_counter [7]}));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  // ../../RTL/CPU/BIU/bus_unit.v(177)
  // ../../RTL/CPU/BIU/bus_unit.v(177)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/bus_unit/reg0_b2|biu/bus_unit/reg0_b6  (
    .c({\biu/bus_unit/n39 [2],\biu/bus_unit/n39 [6]}),
    .ce(\biu/bus_unit/n39[0]_en ),
    .clk(clk_pad),
    .d({\biu/bus_unit/n15_lutinv ,\biu/bus_unit/n15_lutinv }),
    .sr(\biu/bus_unit/n37 ),
    .q({\biu/bus_unit/addr_counter [2],\biu/bus_unit/addr_counter [6]}));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  // ../../RTL/CPU/BIU/bus_unit.v(177)
  // ../../RTL/CPU/BIU/bus_unit.v(177)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("~(~C*~D)"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/bus_unit/reg0_b3|biu/bus_unit/reg0_b5  (
    .c({\biu/bus_unit/n39 [3],\biu/bus_unit/n39 [5]}),
    .ce(\biu/bus_unit/n39[0]_en ),
    .clk(clk_pad),
    .d({\biu/bus_unit/n15_lutinv ,\biu/bus_unit/n15_lutinv }),
    .sr(\biu/bus_unit/n37 ),
    .q({\biu/bus_unit/addr_counter [3],\biu/bus_unit/addr_counter [5]}));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/sub0/u0|biu/bus_unit/sub0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \biu/bus_unit/sub0/u0|biu/bus_unit/sub0/ucin  (
    .a({\biu/bus_unit/addr_counter [0],1'b0}),
    .b({1'b1,open_n76126}),
    .f({\biu/bus_unit/last_addr [0],open_n76146}),
    .fco(\biu/bus_unit/sub0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/sub0/u0|biu/bus_unit/sub0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \biu/bus_unit/sub0/u2|biu/bus_unit/sub0/u1  (
    .a(\biu/bus_unit/addr_counter [2:1]),
    .b(2'b00),
    .fci(\biu/bus_unit/sub0/c1 ),
    .f(\biu/bus_unit/last_addr [2:1]),
    .fco(\biu/bus_unit/sub0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/sub0/u0|biu/bus_unit/sub0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \biu/bus_unit/sub0/u4|biu/bus_unit/sub0/u3  (
    .a(\biu/bus_unit/addr_counter [4:3]),
    .b(2'b00),
    .fci(\biu/bus_unit/sub0/c3 ),
    .f(\biu/bus_unit/last_addr [4:3]),
    .fco(\biu/bus_unit/sub0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/sub0/u0|biu/bus_unit/sub0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \biu/bus_unit/sub0/u6|biu/bus_unit/sub0/u5  (
    .a(\biu/bus_unit/addr_counter [6:5]),
    .b(2'b00),
    .fci(\biu/bus_unit/sub0/c5 ),
    .f(\biu/bus_unit/last_addr [6:5]),
    .fco(\biu/bus_unit/sub0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("biu/bus_unit/sub0/u0|biu/bus_unit/sub0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \biu/bus_unit/sub0/u8|biu/bus_unit/sub0/u7  (
    .a(\biu/bus_unit/addr_counter [8:7]),
    .b(2'b00),
    .fci(\biu/bus_unit/sub0/c7 ),
    .f(\biu/bus_unit/last_addr [8:7]));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0004"),
    //.WID("0x0004"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d00_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76262,\biu/l1i_in [7:0]}),
    .wea(\biu/cache/n1 ),
    .doa({open_n76277,\biu/l1d_out [7:0]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0005"),
    //.WID("0x0005"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d10_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76309,\biu/l1i_in [15:8]}),
    .wea(\biu/cache/n3 ),
    .doa({open_n76324,\biu/l1d_out [15:8]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0006"),
    //.WID("0x0006"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d20_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76356,\biu/l1i_in [23:16]}),
    .wea(\biu/cache/n5 ),
    .doa({open_n76371,\biu/l1d_out [23:16]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0007"),
    //.WID("0x0007"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d30_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76403,\biu/l1i_in [31:24]}),
    .wea(\biu/cache/n7 ),
    .doa({open_n76418,\biu/l1d_out [31:24]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0008"),
    //.WID("0x0008"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d40_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76450,\biu/l1i_in [39:32]}),
    .wea(\biu/cache/n9 ),
    .doa({open_n76465,\biu/l1d_out [39:32]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0009"),
    //.WID("0x0009"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d50_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76497,\biu/l1i_in [47:40]}),
    .wea(\biu/cache/n11 ),
    .doa({open_n76512,\biu/l1d_out [47:40]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000A"),
    //.WID("0x000A"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d60_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76544,\biu/l1i_in [55:48]}),
    .wea(\biu/cache/n13 ),
    .doa({open_n76559,\biu/l1d_out [55:48]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000B"),
    //.WID("0x000B"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d70_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76591,\biu/l1i_in [63:56]}),
    .wea(\biu/cache/n15 ),
    .doa({open_n76606,\biu/l1d_out [63:56]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000C"),
    //.WID("0x000C"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i00_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76638,\biu/l1i_in [7:0]}),
    .wea(\biu/cache/n17 ),
    .doa({open_n76653,ins_read[7:0]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000D"),
    //.WID("0x000D"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i10_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76685,\biu/l1i_in [15:8]}),
    .wea(\biu/cache/n19 ),
    .doa({open_n76700,ins_read[15:8]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000E"),
    //.WID("0x000E"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i20_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76732,\biu/l1i_in [23:16]}),
    .wea(\biu/cache/n21 ),
    .doa({open_n76747,ins_read[23:16]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000F"),
    //.WID("0x000F"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i30_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76779,\biu/l1i_in [31:24]}),
    .wea(\biu/cache/n23 ),
    .doa({open_n76794,ins_read[31:24]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0010"),
    //.WID("0x0010"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i40_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76826,\biu/l1i_in [39:32]}),
    .wea(\biu/cache/n25 ),
    .doa({open_n76841,ins_read[39:32]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0011"),
    //.WID("0x0011"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i50_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76873,\biu/l1i_in [47:40]}),
    .wea(\biu/cache/n27 ),
    .doa({open_n76888,ins_read[47:40]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0012"),
    //.WID("0x0012"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i60_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76920,\biu/l1i_in [55:48]}),
    .wea(\biu/cache/n29 ),
    .doa({open_n76935,ins_read[55:48]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0013"),
    //.WID("0x0013"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i70_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n76967,\biu/l1i_in [63:56]}),
    .wea(\biu/cache/n31 ),
    .doa({open_n76982,ins_read[63:56]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u11_al_u9721  (
    .a({\biu/cache_ctrl_logic/pa_temp [13],\biu/cache_ctrl_logic/pa_temp [11]}),
    .b({\biu/cache_ctrl_logic/pa_temp [14],\biu/cache_ctrl_logic/pa_temp [12]}),
    .c(2'b00),
    .d({1'b0,\biu/cache_ctrl_logic/off [11]}),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c11 ),
    .f({\biu/cache_ctrl_logic/n207 [13],\biu/cache_ctrl_logic/n207 [11]}),
    .fco(\biu/cache_ctrl_logic/add0/c15 ),
    .fx({\biu/cache_ctrl_logic/n207 [14],\biu/cache_ctrl_logic/n207 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u15_al_u9722  (
    .a({\biu/cache_ctrl_logic/pa_temp [17],\biu/cache_ctrl_logic/pa_temp [15]}),
    .b({\biu/cache_ctrl_logic/pa_temp [18],\biu/cache_ctrl_logic/pa_temp [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c15 ),
    .f({\biu/cache_ctrl_logic/n207 [17],\biu/cache_ctrl_logic/n207 [15]}),
    .fco(\biu/cache_ctrl_logic/add0/c19 ),
    .fx({\biu/cache_ctrl_logic/n207 [18],\biu/cache_ctrl_logic/n207 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u19_al_u9723  (
    .a({\biu/cache_ctrl_logic/pa_temp [21],\biu/cache_ctrl_logic/pa_temp [19]}),
    .b({\biu/cache_ctrl_logic/pa_temp [22],\biu/cache_ctrl_logic/pa_temp [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c19 ),
    .f({\biu/cache_ctrl_logic/n207 [21],\biu/cache_ctrl_logic/n207 [19]}),
    .fco(\biu/cache_ctrl_logic/add0/c23 ),
    .fx({\biu/cache_ctrl_logic/n207 [22],\biu/cache_ctrl_logic/n207 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u23_al_u9724  (
    .a({\biu/cache_ctrl_logic/pa_temp [25],\biu/cache_ctrl_logic/pa_temp [23]}),
    .b({\biu/cache_ctrl_logic/pa_temp [26],\biu/cache_ctrl_logic/pa_temp [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c23 ),
    .f({\biu/cache_ctrl_logic/n207 [25],\biu/cache_ctrl_logic/n207 [23]}),
    .fco(\biu/cache_ctrl_logic/add0/c27 ),
    .fx({\biu/cache_ctrl_logic/n207 [26],\biu/cache_ctrl_logic/n207 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u27_al_u9725  (
    .a({\biu/cache_ctrl_logic/pa_temp [29],\biu/cache_ctrl_logic/pa_temp [27]}),
    .b({\biu/cache_ctrl_logic/pa_temp [30],\biu/cache_ctrl_logic/pa_temp [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c27 ),
    .f({\biu/cache_ctrl_logic/n207 [29],\biu/cache_ctrl_logic/n207 [27]}),
    .fco(\biu/cache_ctrl_logic/add0/c31 ),
    .fx({\biu/cache_ctrl_logic/n207 [30],\biu/cache_ctrl_logic/n207 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u31_al_u9726  (
    .a({\biu/cache_ctrl_logic/pa_temp [33],\biu/cache_ctrl_logic/pa_temp [31]}),
    .b({\biu/cache_ctrl_logic/pa_temp [34],\biu/cache_ctrl_logic/pa_temp [32]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c31 ),
    .f({\biu/cache_ctrl_logic/n207 [33],\biu/cache_ctrl_logic/n207 [31]}),
    .fco(\biu/cache_ctrl_logic/add0/c35 ),
    .fx({\biu/cache_ctrl_logic/n207 [34],\biu/cache_ctrl_logic/n207 [32]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u35_al_u9727  (
    .a({\biu/cache_ctrl_logic/pa_temp [37],\biu/cache_ctrl_logic/pa_temp [35]}),
    .b({\biu/cache_ctrl_logic/pa_temp [38],\biu/cache_ctrl_logic/pa_temp [36]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c35 ),
    .f({\biu/cache_ctrl_logic/n207 [37],\biu/cache_ctrl_logic/n207 [35]}),
    .fco(\biu/cache_ctrl_logic/add0/c39 ),
    .fx({\biu/cache_ctrl_logic/n207 [38],\biu/cache_ctrl_logic/n207 [36]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u39_al_u9728  (
    .a({\biu/cache_ctrl_logic/pa_temp [41],\biu/cache_ctrl_logic/pa_temp [39]}),
    .b({\biu/cache_ctrl_logic/pa_temp [42],\biu/cache_ctrl_logic/pa_temp [40]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c39 ),
    .f({\biu/cache_ctrl_logic/n207 [41],\biu/cache_ctrl_logic/n207 [39]}),
    .fco(\biu/cache_ctrl_logic/add0/c43 ),
    .fx({\biu/cache_ctrl_logic/n207 [42],\biu/cache_ctrl_logic/n207 [40]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u3_al_u9719  (
    .a({\biu/cache_ctrl_logic/pa_temp [5],\biu/cache_ctrl_logic/pa_temp [3]}),
    .b({\biu/cache_ctrl_logic/pa_temp [6],\biu/cache_ctrl_logic/pa_temp [4]}),
    .c(2'b00),
    .d({\biu/cache_ctrl_logic/off [5],\biu/cache_ctrl_logic/off [3]}),
    .e({\biu/cache_ctrl_logic/off [6],\biu/cache_ctrl_logic/off [4]}),
    .fci(\biu/cache_ctrl_logic/add0/c3 ),
    .f({\biu/cache_ctrl_logic/n207 [5],\biu/cache_ctrl_logic/n207 [3]}),
    .fco(\biu/cache_ctrl_logic/add0/c7 ),
    .fx({\biu/cache_ctrl_logic/n207 [6],\biu/cache_ctrl_logic/n207 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u43_al_u9729  (
    .a({\biu/cache_ctrl_logic/pa_temp [45],\biu/cache_ctrl_logic/pa_temp [43]}),
    .b({\biu/cache_ctrl_logic/pa_temp [46],\biu/cache_ctrl_logic/pa_temp [44]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c43 ),
    .f({\biu/cache_ctrl_logic/n207 [45],\biu/cache_ctrl_logic/n207 [43]}),
    .fco(\biu/cache_ctrl_logic/add0/c47 ),
    .fx({\biu/cache_ctrl_logic/n207 [46],\biu/cache_ctrl_logic/n207 [44]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u47_al_u9730  (
    .a({\biu/cache_ctrl_logic/pa_temp [49],\biu/cache_ctrl_logic/pa_temp [47]}),
    .b({\biu/cache_ctrl_logic/pa_temp [50],\biu/cache_ctrl_logic/pa_temp [48]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c47 ),
    .f({\biu/cache_ctrl_logic/n207 [49],\biu/cache_ctrl_logic/n207 [47]}),
    .fco(\biu/cache_ctrl_logic/add0/c51 ),
    .fx({\biu/cache_ctrl_logic/n207 [50],\biu/cache_ctrl_logic/n207 [48]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u51_al_u9731  (
    .a({\biu/cache_ctrl_logic/pa_temp [53],\biu/cache_ctrl_logic/pa_temp [51]}),
    .b({\biu/cache_ctrl_logic/pa_temp [54],\biu/cache_ctrl_logic/pa_temp [52]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c51 ),
    .f({\biu/cache_ctrl_logic/n207 [53],\biu/cache_ctrl_logic/n207 [51]}),
    .fco(\biu/cache_ctrl_logic/add0/c55 ),
    .fx({\biu/cache_ctrl_logic/n207 [54],\biu/cache_ctrl_logic/n207 [52]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u55_al_u9732  (
    .a({\biu/cache_ctrl_logic/pa_temp [57],\biu/cache_ctrl_logic/pa_temp [55]}),
    .b({\biu/cache_ctrl_logic/pa_temp [58],\biu/cache_ctrl_logic/pa_temp [56]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c55 ),
    .f({\biu/cache_ctrl_logic/n207 [57],\biu/cache_ctrl_logic/n207 [55]}),
    .fco(\biu/cache_ctrl_logic/add0/c59 ),
    .fx({\biu/cache_ctrl_logic/n207 [58],\biu/cache_ctrl_logic/n207 [56]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u59_al_u9733  (
    .a({\biu/cache_ctrl_logic/pa_temp [61],\biu/cache_ctrl_logic/pa_temp [59]}),
    .b({\biu/cache_ctrl_logic/pa_temp [62],\biu/cache_ctrl_logic/pa_temp [60]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add0/c59 ),
    .f({\biu/cache_ctrl_logic/n207 [61],\biu/cache_ctrl_logic/n207 [59]}),
    .fco(\biu/cache_ctrl_logic/add0/c63 ),
    .fx({\biu/cache_ctrl_logic/n207 [62],\biu/cache_ctrl_logic/n207 [60]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y8Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u63_al_u9734  (
    .a({open_n77244,\biu/cache_ctrl_logic/pa_temp [63]}),
    .c(2'b00),
    .d({open_n77249,1'b0}),
    .fci(\biu/cache_ctrl_logic/add0/c63 ),
    .f({open_n77266,\biu/cache_ctrl_logic/n207 [63]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add0/u7_al_u9720  (
    .a({\biu/cache_ctrl_logic/pa_temp [9],\biu/cache_ctrl_logic/pa_temp [7]}),
    .b({\biu/cache_ctrl_logic/pa_temp [10],\biu/cache_ctrl_logic/pa_temp [8]}),
    .c(2'b00),
    .d({\biu/cache_ctrl_logic/off [9],\biu/cache_ctrl_logic/off [7]}),
    .e({\biu/cache_ctrl_logic/off [10],\biu/cache_ctrl_logic/off [8]}),
    .fci(\biu/cache_ctrl_logic/add0/c7 ),
    .f({\biu/cache_ctrl_logic/n207 [9],\biu/cache_ctrl_logic/n207 [7]}),
    .fco(\biu/cache_ctrl_logic/add0/c11 ),
    .fx({\biu/cache_ctrl_logic/n207 [10],\biu/cache_ctrl_logic/n207 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add0/ucin_al_u9718"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/add0/ucin_al_u9718  (
    .a({\biu/cache_ctrl_logic/pa_temp [1],1'b0}),
    .b({\biu/cache_ctrl_logic/pa_temp [2],\biu/cache_ctrl_logic/pa_temp [0]}),
    .c(2'b00),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/off [1],1'b1}),
    .e({\biu/cache_ctrl_logic/off [2],\biu/cache_ctrl_logic/off [0]}),
    .mi(\biu/cache_ctrl_logic/pa_temp [1:0]),
    .sr(rst_pad),
    .f({\biu/cache_ctrl_logic/n207 [1],open_n77302}),
    .fco(\biu/cache_ctrl_logic/add0/c3 ),
    .fx({\biu/cache_ctrl_logic/n207 [2],\biu/cache_ctrl_logic/n207 [0]}),
    .q(\biu/cache_ctrl_logic/l1i_pa [1:0]));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u11_al_u9738  (
    .a({\biu/cache_ctrl_logic/l1i_pa [13],\biu/cache_ctrl_logic/l1i_pa [11]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [14],\biu/cache_ctrl_logic/l1i_pa [12]}),
    .c(2'b00),
    .d({1'b0,\biu/cache_ctrl_logic/off [11]}),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c11 ),
    .f({\biu/cache_ctrl_logic/n209 [13],\biu/cache_ctrl_logic/n209 [11]}),
    .fco(\biu/cache_ctrl_logic/add1/c15 ),
    .fx({\biu/cache_ctrl_logic/n209 [14],\biu/cache_ctrl_logic/n209 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u15_al_u9739  (
    .a({\biu/cache_ctrl_logic/l1i_pa [17],\biu/cache_ctrl_logic/l1i_pa [15]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [18],\biu/cache_ctrl_logic/l1i_pa [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c15 ),
    .f({\biu/cache_ctrl_logic/n209 [17],\biu/cache_ctrl_logic/n209 [15]}),
    .fco(\biu/cache_ctrl_logic/add1/c19 ),
    .fx({\biu/cache_ctrl_logic/n209 [18],\biu/cache_ctrl_logic/n209 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u19_al_u9740  (
    .a({\biu/cache_ctrl_logic/l1i_pa [21],\biu/cache_ctrl_logic/l1i_pa [19]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [22],\biu/cache_ctrl_logic/l1i_pa [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c19 ),
    .f({\biu/cache_ctrl_logic/n209 [21],\biu/cache_ctrl_logic/n209 [19]}),
    .fco(\biu/cache_ctrl_logic/add1/c23 ),
    .fx({\biu/cache_ctrl_logic/n209 [22],\biu/cache_ctrl_logic/n209 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u23_al_u9741  (
    .a({\biu/cache_ctrl_logic/l1i_pa [25],\biu/cache_ctrl_logic/l1i_pa [23]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [26],\biu/cache_ctrl_logic/l1i_pa [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c23 ),
    .f({\biu/cache_ctrl_logic/n209 [25],\biu/cache_ctrl_logic/n209 [23]}),
    .fco(\biu/cache_ctrl_logic/add1/c27 ),
    .fx({\biu/cache_ctrl_logic/n209 [26],\biu/cache_ctrl_logic/n209 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u27_al_u9742  (
    .a({\biu/cache_ctrl_logic/l1i_pa [29],\biu/cache_ctrl_logic/l1i_pa [27]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [30],\biu/cache_ctrl_logic/l1i_pa [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c27 ),
    .f({\biu/cache_ctrl_logic/n209 [29],\biu/cache_ctrl_logic/n209 [27]}),
    .fco(\biu/cache_ctrl_logic/add1/c31 ),
    .fx({\biu/cache_ctrl_logic/n209 [30],\biu/cache_ctrl_logic/n209 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u31_al_u9743  (
    .a({\biu/cache_ctrl_logic/l1i_pa [33],\biu/cache_ctrl_logic/l1i_pa [31]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [34],\biu/cache_ctrl_logic/l1i_pa [32]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c31 ),
    .f({\biu/cache_ctrl_logic/n209 [33],\biu/cache_ctrl_logic/n209 [31]}),
    .fco(\biu/cache_ctrl_logic/add1/c35 ),
    .fx({\biu/cache_ctrl_logic/n209 [34],\biu/cache_ctrl_logic/n209 [32]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u35_al_u9744  (
    .a({\biu/cache_ctrl_logic/l1i_pa [37],\biu/cache_ctrl_logic/l1i_pa [35]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [38],\biu/cache_ctrl_logic/l1i_pa [36]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c35 ),
    .f({\biu/cache_ctrl_logic/n209 [37],\biu/cache_ctrl_logic/n209 [35]}),
    .fco(\biu/cache_ctrl_logic/add1/c39 ),
    .fx({\biu/cache_ctrl_logic/n209 [38],\biu/cache_ctrl_logic/n209 [36]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u39_al_u9745  (
    .a({\biu/cache_ctrl_logic/l1i_pa [41],\biu/cache_ctrl_logic/l1i_pa [39]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [42],\biu/cache_ctrl_logic/l1i_pa [40]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c39 ),
    .f({\biu/cache_ctrl_logic/n209 [41],\biu/cache_ctrl_logic/n209 [39]}),
    .fco(\biu/cache_ctrl_logic/add1/c43 ),
    .fx({\biu/cache_ctrl_logic/n209 [42],\biu/cache_ctrl_logic/n209 [40]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u3_al_u9736  (
    .a({\biu/cache_ctrl_logic/l1i_pa [5],\biu/cache_ctrl_logic/l1i_pa [3]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [6],\biu/cache_ctrl_logic/l1i_pa [4]}),
    .c(2'b00),
    .d({\biu/cache_ctrl_logic/off [5],\biu/cache_ctrl_logic/off [3]}),
    .e({\biu/cache_ctrl_logic/off [6],\biu/cache_ctrl_logic/off [4]}),
    .fci(\biu/cache_ctrl_logic/add1/c3 ),
    .f({\biu/cache_ctrl_logic/n209 [5],\biu/cache_ctrl_logic/n209 [3]}),
    .fco(\biu/cache_ctrl_logic/add1/c7 ),
    .fx({\biu/cache_ctrl_logic/n209 [6],\biu/cache_ctrl_logic/n209 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u43_al_u9746  (
    .a({\biu/cache_ctrl_logic/l1i_pa [45],\biu/cache_ctrl_logic/l1i_pa [43]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [46],\biu/cache_ctrl_logic/l1i_pa [44]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c43 ),
    .f({\biu/cache_ctrl_logic/n209 [45],\biu/cache_ctrl_logic/n209 [43]}),
    .fco(\biu/cache_ctrl_logic/add1/c47 ),
    .fx({\biu/cache_ctrl_logic/n209 [46],\biu/cache_ctrl_logic/n209 [44]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u47_al_u9747  (
    .a({\biu/cache_ctrl_logic/l1i_pa [49],\biu/cache_ctrl_logic/l1i_pa [47]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [50],\biu/cache_ctrl_logic/l1i_pa [48]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c47 ),
    .f({\biu/cache_ctrl_logic/n209 [49],\biu/cache_ctrl_logic/n209 [47]}),
    .fco(\biu/cache_ctrl_logic/add1/c51 ),
    .fx({\biu/cache_ctrl_logic/n209 [50],\biu/cache_ctrl_logic/n209 [48]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u51_al_u9748  (
    .a({\biu/cache_ctrl_logic/l1i_pa [53],\biu/cache_ctrl_logic/l1i_pa [51]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [54],\biu/cache_ctrl_logic/l1i_pa [52]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c51 ),
    .f({\biu/cache_ctrl_logic/n209 [53],\biu/cache_ctrl_logic/n209 [51]}),
    .fco(\biu/cache_ctrl_logic/add1/c55 ),
    .fx({\biu/cache_ctrl_logic/n209 [54],\biu/cache_ctrl_logic/n209 [52]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u55_al_u9749  (
    .a({\biu/cache_ctrl_logic/l1i_pa [57],\biu/cache_ctrl_logic/l1i_pa [55]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [58],\biu/cache_ctrl_logic/l1i_pa [56]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c55 ),
    .f({\biu/cache_ctrl_logic/n209 [57],\biu/cache_ctrl_logic/n209 [55]}),
    .fco(\biu/cache_ctrl_logic/add1/c59 ),
    .fx({\biu/cache_ctrl_logic/n209 [58],\biu/cache_ctrl_logic/n209 [56]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u59_al_u9750  (
    .a({\biu/cache_ctrl_logic/l1i_pa [61],\biu/cache_ctrl_logic/l1i_pa [59]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [62],\biu/cache_ctrl_logic/l1i_pa [60]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add1/c59 ),
    .f({\biu/cache_ctrl_logic/n209 [61],\biu/cache_ctrl_logic/n209 [59]}),
    .fco(\biu/cache_ctrl_logic/add1/c63 ),
    .fx({\biu/cache_ctrl_logic/n209 [62],\biu/cache_ctrl_logic/n209 [60]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y8Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u63_al_u9751  (
    .a({open_n77555,\biu/cache_ctrl_logic/l1i_pa [63]}),
    .c(2'b00),
    .d({open_n77560,1'b0}),
    .fci(\biu/cache_ctrl_logic/add1/c63 ),
    .f({open_n77577,\biu/cache_ctrl_logic/n209 [63]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add1/u7_al_u9737  (
    .a({\biu/cache_ctrl_logic/l1i_pa [9],\biu/cache_ctrl_logic/l1i_pa [7]}),
    .b({\biu/cache_ctrl_logic/l1i_pa [10],\biu/cache_ctrl_logic/l1i_pa [8]}),
    .c(2'b00),
    .d({\biu/cache_ctrl_logic/off [9],\biu/cache_ctrl_logic/off [7]}),
    .e({\biu/cache_ctrl_logic/off [10],\biu/cache_ctrl_logic/off [8]}),
    .fci(\biu/cache_ctrl_logic/add1/c7 ),
    .f({\biu/cache_ctrl_logic/n209 [9],\biu/cache_ctrl_logic/n209 [7]}),
    .fco(\biu/cache_ctrl_logic/add1/c11 ),
    .fx({\biu/cache_ctrl_logic/n209 [10],\biu/cache_ctrl_logic/n209 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add1/ucin_al_u9735"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/add1/ucin_al_u9735  (
    .a({\biu/cache_ctrl_logic/l1i_pa [1],1'b0}),
    .b({\biu/cache_ctrl_logic/l1i_pa [2],\biu/cache_ctrl_logic/l1i_pa [0]}),
    .c(2'b00),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/off [1],1'b1}),
    .e({\biu/cache_ctrl_logic/off [2],\biu/cache_ctrl_logic/off [0]}),
    .mi({open_n77602,\biu/cache_ctrl_logic/pa_temp [2]}),
    .sr(rst_pad),
    .f({\biu/cache_ctrl_logic/n209 [1],open_n77614}),
    .fco(\biu/cache_ctrl_logic/add1/c3 ),
    .fx({\biu/cache_ctrl_logic/n209 [2],\biu/cache_ctrl_logic/n209 [0]}),
    .q({open_n77615,\biu/cache_ctrl_logic/l1i_pa [2]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u11_al_u9755  (
    .a({\biu/cache_ctrl_logic/l1d_pa [13],\biu/cache_ctrl_logic/l1d_pa [11]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [14],\biu/cache_ctrl_logic/l1d_pa [12]}),
    .c(2'b00),
    .d({1'b0,\biu/cache_ctrl_logic/off [11]}),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c11 ),
    .f({\biu/cache_ctrl_logic/n212 [13],\biu/cache_ctrl_logic/n212 [11]}),
    .fco(\biu/cache_ctrl_logic/add2/c15 ),
    .fx({\biu/cache_ctrl_logic/n212 [14],\biu/cache_ctrl_logic/n212 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u15_al_u9756  (
    .a({\biu/cache_ctrl_logic/l1d_pa [17],\biu/cache_ctrl_logic/l1d_pa [15]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [18],\biu/cache_ctrl_logic/l1d_pa [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c15 ),
    .f({\biu/cache_ctrl_logic/n212 [17],\biu/cache_ctrl_logic/n212 [15]}),
    .fco(\biu/cache_ctrl_logic/add2/c19 ),
    .fx({\biu/cache_ctrl_logic/n212 [18],\biu/cache_ctrl_logic/n212 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u19_al_u9757  (
    .a({\biu/cache_ctrl_logic/l1d_pa [21],\biu/cache_ctrl_logic/l1d_pa [19]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [22],\biu/cache_ctrl_logic/l1d_pa [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c19 ),
    .f({\biu/cache_ctrl_logic/n212 [21],\biu/cache_ctrl_logic/n212 [19]}),
    .fco(\biu/cache_ctrl_logic/add2/c23 ),
    .fx({\biu/cache_ctrl_logic/n212 [22],\biu/cache_ctrl_logic/n212 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u23_al_u9758  (
    .a({\biu/cache_ctrl_logic/l1d_pa [25],\biu/cache_ctrl_logic/l1d_pa [23]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [26],\biu/cache_ctrl_logic/l1d_pa [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c23 ),
    .f({\biu/cache_ctrl_logic/n212 [25],\biu/cache_ctrl_logic/n212 [23]}),
    .fco(\biu/cache_ctrl_logic/add2/c27 ),
    .fx({\biu/cache_ctrl_logic/n212 [26],\biu/cache_ctrl_logic/n212 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u27_al_u9759  (
    .a({\biu/cache_ctrl_logic/l1d_pa [29],\biu/cache_ctrl_logic/l1d_pa [27]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [30],\biu/cache_ctrl_logic/l1d_pa [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c27 ),
    .f({\biu/cache_ctrl_logic/n212 [29],\biu/cache_ctrl_logic/n212 [27]}),
    .fco(\biu/cache_ctrl_logic/add2/c31 ),
    .fx({\biu/cache_ctrl_logic/n212 [30],\biu/cache_ctrl_logic/n212 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u31_al_u9760  (
    .a({\biu/cache_ctrl_logic/l1d_pa [33],\biu/cache_ctrl_logic/l1d_pa [31]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [34],\biu/cache_ctrl_logic/l1d_pa [32]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c31 ),
    .f({\biu/cache_ctrl_logic/n212 [33],\biu/cache_ctrl_logic/n212 [31]}),
    .fco(\biu/cache_ctrl_logic/add2/c35 ),
    .fx({\biu/cache_ctrl_logic/n212 [34],\biu/cache_ctrl_logic/n212 [32]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u35_al_u9761  (
    .a({\biu/cache_ctrl_logic/l1d_pa [37],\biu/cache_ctrl_logic/l1d_pa [35]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [38],\biu/cache_ctrl_logic/l1d_pa [36]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c35 ),
    .f({\biu/cache_ctrl_logic/n212 [37],\biu/cache_ctrl_logic/n212 [35]}),
    .fco(\biu/cache_ctrl_logic/add2/c39 ),
    .fx({\biu/cache_ctrl_logic/n212 [38],\biu/cache_ctrl_logic/n212 [36]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u39_al_u9762  (
    .a({\biu/cache_ctrl_logic/l1d_pa [41],\biu/cache_ctrl_logic/l1d_pa [39]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [42],\biu/cache_ctrl_logic/l1d_pa [40]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c39 ),
    .f({\biu/cache_ctrl_logic/n212 [41],\biu/cache_ctrl_logic/n212 [39]}),
    .fco(\biu/cache_ctrl_logic/add2/c43 ),
    .fx({\biu/cache_ctrl_logic/n212 [42],\biu/cache_ctrl_logic/n212 [40]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u3_al_u9753  (
    .a({\biu/cache_ctrl_logic/l1d_pa [5],\biu/cache_ctrl_logic/l1d_pa [3]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [6],\biu/cache_ctrl_logic/l1d_pa [4]}),
    .c(2'b00),
    .d({\biu/cache_ctrl_logic/off [5],\biu/cache_ctrl_logic/off [3]}),
    .e({\biu/cache_ctrl_logic/off [6],\biu/cache_ctrl_logic/off [4]}),
    .fci(\biu/cache_ctrl_logic/add2/c3 ),
    .f({\biu/cache_ctrl_logic/n212 [5],\biu/cache_ctrl_logic/n212 [3]}),
    .fco(\biu/cache_ctrl_logic/add2/c7 ),
    .fx({\biu/cache_ctrl_logic/n212 [6],\biu/cache_ctrl_logic/n212 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u43_al_u9763  (
    .a({\biu/cache_ctrl_logic/l1d_pa [45],\biu/cache_ctrl_logic/l1d_pa [43]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [46],\biu/cache_ctrl_logic/l1d_pa [44]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c43 ),
    .f({\biu/cache_ctrl_logic/n212 [45],\biu/cache_ctrl_logic/n212 [43]}),
    .fco(\biu/cache_ctrl_logic/add2/c47 ),
    .fx({\biu/cache_ctrl_logic/n212 [46],\biu/cache_ctrl_logic/n212 [44]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u47_al_u9764  (
    .a({\biu/cache_ctrl_logic/l1d_pa [49],\biu/cache_ctrl_logic/l1d_pa [47]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [50],\biu/cache_ctrl_logic/l1d_pa [48]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c47 ),
    .f({\biu/cache_ctrl_logic/n212 [49],\biu/cache_ctrl_logic/n212 [47]}),
    .fco(\biu/cache_ctrl_logic/add2/c51 ),
    .fx({\biu/cache_ctrl_logic/n212 [50],\biu/cache_ctrl_logic/n212 [48]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u51_al_u9765  (
    .a({\biu/cache_ctrl_logic/l1d_pa [53],\biu/cache_ctrl_logic/l1d_pa [51]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [54],\biu/cache_ctrl_logic/l1d_pa [52]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c51 ),
    .f({\biu/cache_ctrl_logic/n212 [53],\biu/cache_ctrl_logic/n212 [51]}),
    .fco(\biu/cache_ctrl_logic/add2/c55 ),
    .fx({\biu/cache_ctrl_logic/n212 [54],\biu/cache_ctrl_logic/n212 [52]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u55_al_u9766  (
    .a({\biu/cache_ctrl_logic/l1d_pa [57],\biu/cache_ctrl_logic/l1d_pa [55]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [58],\biu/cache_ctrl_logic/l1d_pa [56]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c55 ),
    .f({\biu/cache_ctrl_logic/n212 [57],\biu/cache_ctrl_logic/n212 [55]}),
    .fco(\biu/cache_ctrl_logic/add2/c59 ),
    .fx({\biu/cache_ctrl_logic/n212 [58],\biu/cache_ctrl_logic/n212 [56]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u59_al_u9767  (
    .a({\biu/cache_ctrl_logic/l1d_pa [61],\biu/cache_ctrl_logic/l1d_pa [59]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [62],\biu/cache_ctrl_logic/l1d_pa [60]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\biu/cache_ctrl_logic/add2/c59 ),
    .f({\biu/cache_ctrl_logic/n212 [61],\biu/cache_ctrl_logic/n212 [59]}),
    .fco(\biu/cache_ctrl_logic/add2/c63 ),
    .fx({\biu/cache_ctrl_logic/n212 [62],\biu/cache_ctrl_logic/n212 [60]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y8Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u63_al_u9768  (
    .a({open_n77868,\biu/cache_ctrl_logic/l1d_pa [63]}),
    .c(2'b00),
    .d({open_n77873,1'b0}),
    .fci(\biu/cache_ctrl_logic/add2/c63 ),
    .f({open_n77890,\biu/cache_ctrl_logic/n212 [63]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \biu/cache_ctrl_logic/add2/u7_al_u9754  (
    .a({\biu/cache_ctrl_logic/l1d_pa [9],\biu/cache_ctrl_logic/l1d_pa [7]}),
    .b({\biu/cache_ctrl_logic/l1d_pa [10],\biu/cache_ctrl_logic/l1d_pa [8]}),
    .c(2'b00),
    .d({\biu/cache_ctrl_logic/off [9],\biu/cache_ctrl_logic/off [7]}),
    .e({\biu/cache_ctrl_logic/off [10],\biu/cache_ctrl_logic/off [8]}),
    .fci(\biu/cache_ctrl_logic/add2/c7 ),
    .f({\biu/cache_ctrl_logic/n212 [9],\biu/cache_ctrl_logic/n212 [7]}),
    .fco(\biu/cache_ctrl_logic/add2/c11 ),
    .fx({\biu/cache_ctrl_logic/n212 [10],\biu/cache_ctrl_logic/n212 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("biu/cache_ctrl_logic/add2/ucin_al_u9752"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/add2/ucin_al_u9752  (
    .a({\biu/cache_ctrl_logic/l1d_pa [1],1'b0}),
    .b({\biu/cache_ctrl_logic/l1d_pa [2],\biu/cache_ctrl_logic/l1d_pa [0]}),
    .c(2'b00),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/off [1],1'b1}),
    .e({\biu/cache_ctrl_logic/off [2],\biu/cache_ctrl_logic/off [0]}),
    .mi(\biu/cache_ctrl_logic/pa_temp [1:0]),
    .sr(rst_pad),
    .f({\biu/cache_ctrl_logic/n212 [1],open_n77926}),
    .fco(\biu/cache_ctrl_logic/add2/c3 ),
    .fx({\biu/cache_ctrl_logic/n212 [2],\biu/cache_ctrl_logic/n212 [0]}),
    .q(\biu/cache_ctrl_logic/l1d_pa [1:0]));
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(394)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(347)
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \biu/cache_ctrl_logic/l1i_value_reg|biu/cache_ctrl_logic/l1d_value_reg  (
    .c({\biu/cache_ctrl_logic/l1i_value ,\biu/cache_ctrl_logic/l1d_value }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/n135 ,\biu/cache_ctrl_logic/n149 }),
    .sr(\biu/cache_ctrl_logic/u128_sel_is_0_o ),
    .q({\biu/cache_ctrl_logic/l1i_value ,\biu/cache_ctrl_logic/l1d_value }));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(394)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0000001000010011),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0000001000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b12|biu/cache_ctrl_logic/reg2_b36  (
    .a({\ins_fetch/n27 ,_al_u3945_o}),
    .b({pip_flush,_al_u3950_o}),
    .c({\ins_fetch/n1 [10],\biu/cache_ctrl_logic/l1i_pte [36]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[12],\biu/cache_ctrl_logic/pte_temp [36]}),
    .mi({addr_if[12],\biu/cache_ctrl_logic/pte_temp [36]}),
    .sr(rst_pad),
    .f({_al_u9664_o,_al_u5784_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [12],\biu/cache_ctrl_logic/l1i_pte [36]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b13|biu/cache_ctrl_logic/reg0_b63  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [11],\ins_fetch/n1 [61]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[13],addr_if[63]}),
    .mi({addr_if[13],addr_if[63]}),
    .sr(rst_pad),
    .f({_al_u9657_o,_al_u9311_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [13],\biu/cache_ctrl_logic/l1i_va [63]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000100100000),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b14|biu/cache_ctrl_logic/reg0_b62  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [12],\ins_fetch/n1 [60]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[14],addr_if[62]}),
    .mi({addr_if[14],addr_if[62]}),
    .sr(rst_pad),
    .f({_al_u9650_o,_al_u9317_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [14],\biu/cache_ctrl_logic/l1i_va [62]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000001000010011),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000001000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b15|biu/cache_ctrl_logic/reg0_b58  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [13],\ins_fetch/n1 [56]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[15],addr_if[58]}),
    .mi({addr_if[15],addr_if[58]}),
    .sr(rst_pad),
    .f({_al_u9645_o,_al_u9340_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [15],\biu/cache_ctrl_logic/l1i_va [58]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000001000010011),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000001000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b16|biu/cache_ctrl_logic/reg0_b54  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [14],\ins_fetch/n1 [52]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[16],addr_if[54]}),
    .mi({addr_if[16],addr_if[54]}),
    .sr(rst_pad),
    .f({_al_u9638_o,_al_u9366_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [16],\biu/cache_ctrl_logic/l1i_va [54]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b17|biu/cache_ctrl_logic/reg0_b50  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [15],\ins_fetch/n1 [48]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[17],addr_if[50]}),
    .mi({addr_if[17],addr_if[50]}),
    .sr(rst_pad),
    .f({_al_u9631_o,_al_u9399_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [17],\biu/cache_ctrl_logic/l1i_va [50]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b18|biu/cache_ctrl_logic/reg0_b38  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [16],\ins_fetch/n1 [36]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[18],addr_if[38]}),
    .mi({addr_if[18],addr_if[38]}),
    .sr(rst_pad),
    .f({_al_u9624_o,_al_u9480_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [18],\biu/cache_ctrl_logic/l1i_va [38]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000001000010011),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000001000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b19|biu/cache_ctrl_logic/reg0_b34  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [17],\ins_fetch/n1 [32]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[19],addr_if[34]}),
    .mi({addr_if[19],addr_if[34]}),
    .sr(rst_pad),
    .f({_al_u9619_o,_al_u9506_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [19],\biu/cache_ctrl_logic/l1i_va [34]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000001000010011),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000001000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b20|biu/cache_ctrl_logic/reg0_b26  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [18],\ins_fetch/n1 [24]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[20],addr_if[26]}),
    .mi({addr_if[20],addr_if[26]}),
    .sr(rst_pad),
    .f({_al_u9612_o,_al_u9565_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [20],\biu/cache_ctrl_logic/l1i_va [26]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b21|biu/cache_ctrl_logic/reg0_b60  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [19],\ins_fetch/n1 [58]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[21],addr_if[60]}),
    .mi({addr_if[21],addr_if[60]}),
    .sr(rst_pad),
    .f({_al_u9605_o,_al_u9330_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [21],\biu/cache_ctrl_logic/l1i_va [60]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000001000010011),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000001000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b22|biu/cache_ctrl_logic/reg0_b49  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [20],\ins_fetch/n1 [47]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[22],addr_if[49]}),
    .mi({addr_if[22],addr_if[49]}),
    .sr(rst_pad),
    .f({_al_u9591_o,_al_u9404_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [22],\biu/cache_ctrl_logic/l1i_va [49]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b23|biu/cache_ctrl_logic/reg0_b48  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [21],\ins_fetch/n1 [46]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[23],addr_if[48]}),
    .mi({addr_if[23],addr_if[48]}),
    .sr(rst_pad),
    .f({_al_u9586_o,_al_u9411_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [23],\biu/cache_ctrl_logic/l1i_va [48]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b25|biu/cache_ctrl_logic/reg0_b39  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [23],\ins_fetch/n1 [37]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[25],addr_if[39]}),
    .mi({addr_if[25],addr_if[39]}),
    .sr(rst_pad),
    .f({_al_u9572_o,_al_u9473_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [25],\biu/cache_ctrl_logic/l1i_va [39]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b27|biu/cache_ctrl_logic/reg0_b56  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [25],\ins_fetch/n1 [54]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[27],addr_if[56]}),
    .mi({addr_if[27],addr_if[56]}),
    .sr(rst_pad),
    .f({_al_u9558_o,_al_u9352_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [27],\biu/cache_ctrl_logic/l1i_va [56]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000001000010011),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000001000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b29|biu/cache_ctrl_logic/reg0_b45  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [27],\ins_fetch/n1 [43]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[29],addr_if[45]}),
    .mi({addr_if[29],addr_if[45]}),
    .sr(rst_pad),
    .f({_al_u9544_o,_al_u9430_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [29],\biu/cache_ctrl_logic/l1i_va [45]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b31|biu/cache_ctrl_logic/reg0_b57  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [29],\ins_fetch/n1 [55]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[31],addr_if[57]}),
    .mi({addr_if[31],addr_if[57]}),
    .sr(rst_pad),
    .f({_al_u9530_o,_al_u9345_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [31],\biu/cache_ctrl_logic/l1i_va [57]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b33|biu/cache_ctrl_logic/reg0_b55  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [31],\ins_fetch/n1 [53]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[33],addr_if[55]}),
    .mi({addr_if[33],addr_if[55]}),
    .sr(rst_pad),
    .f({_al_u9513_o,_al_u9359_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [33],\biu/cache_ctrl_logic/l1i_va [55]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b0000001000010011),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b0000001000010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b35|biu/cache_ctrl_logic/reg0_b51  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [33],\ins_fetch/n1 [49]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[35],addr_if[51]}),
    .mi({addr_if[35],addr_if[51]}),
    .sr(rst_pad),
    .f({_al_u9499_o,_al_u9392_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [35],\biu/cache_ctrl_logic/l1i_va [51]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg0_b41|biu/cache_ctrl_logic/reg0_b47  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [39],\ins_fetch/n1 [45]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({addr_if[41],addr_if[47]}),
    .mi({addr_if[41],addr_if[47]}),
    .sr(rst_pad),
    .f({_al_u9461_o,_al_u9418_o}),
    .q({\biu/cache_ctrl_logic/l1i_va [41],\biu/cache_ctrl_logic/l1i_va [47]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b100|biu/cache_ctrl_logic/reg1_b96  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [100],\biu/cache_ctrl_logic/l1i_pa [96]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pa_temp [100],\biu/cache_ctrl_logic/pa_temp [96]}),
    .mi({\biu/cache_ctrl_logic/pa_temp [100],\biu/cache_ctrl_logic/pa_temp [96]}),
    .sr(rst_pad),
    .f({_al_u4600_o,_al_u4624_o}),
    .q({\biu/cache_ctrl_logic/l1i_pa [100],\biu/cache_ctrl_logic/l1i_pa [96]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b101|biu/cache_ctrl_logic/reg1_b68  (
    .a({\biu/cache_ctrl_logic/n75_lutinv ,_al_u3945_o}),
    .b({_al_u3945_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [101],\biu/cache_ctrl_logic/l1i_pa [68]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({addr_ex[37],\biu/cache_ctrl_logic/pa_temp [68]}),
    .mi({\biu/cache_ctrl_logic/pa_temp [101],\biu/cache_ctrl_logic/pa_temp [68]}),
    .sr(rst_pad),
    .f({_al_u4594_o,_al_u4576_o}),
    .q({\biu/cache_ctrl_logic/l1i_pa [101],\biu/cache_ctrl_logic/l1i_pa [68]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b106|biu/cache_ctrl_logic/reg1_b94  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [106],\biu/cache_ctrl_logic/l1i_pa [94]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pa_temp [106],\biu/cache_ctrl_logic/pa_temp [94]}),
    .mi({\biu/cache_ctrl_logic/pa_temp [106],\biu/cache_ctrl_logic/pa_temp [94]}),
    .sr(rst_pad),
    .f({_al_u4558_o,_al_u4636_o}),
    .q({\biu/cache_ctrl_logic/l1i_pa [106],\biu/cache_ctrl_logic/l1i_pa [94]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b10|biu/cache_ctrl_logic/reg1_b9  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi(\biu/cache_ctrl_logic/pa_temp [10:9]),
    .sr(rst_pad),
    .q(\biu/cache_ctrl_logic/l1i_pa [10:9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b116|biu/cache_ctrl_logic/reg1_b93  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [116],\biu/cache_ctrl_logic/l1i_pa [93]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pa_temp [116],\biu/cache_ctrl_logic/pa_temp [93]}),
    .mi({\biu/cache_ctrl_logic/pa_temp [116],\biu/cache_ctrl_logic/pa_temp [93]}),
    .sr(rst_pad),
    .f({_al_u4492_o,_al_u4648_o}),
    .q({\biu/cache_ctrl_logic/l1i_pa [116],\biu/cache_ctrl_logic/l1i_pa [93]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b117|biu/cache_ctrl_logic/reg1_b83  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [117],\biu/cache_ctrl_logic/l1i_pa [83]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pa_temp [117],\biu/cache_ctrl_logic/pa_temp [83]}),
    .mi({\biu/cache_ctrl_logic/pa_temp [117],\biu/cache_ctrl_logic/pa_temp [83]}),
    .sr(rst_pad),
    .f({_al_u4486_o,_al_u4708_o}),
    .q({\biu/cache_ctrl_logic/l1i_pa [117],\biu/cache_ctrl_logic/l1i_pa [83]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b11|biu/cache_ctrl_logic/reg1_b8  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [11],\biu/cache_ctrl_logic/pa_temp [8]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [11],\biu/cache_ctrl_logic/l1i_pa [8]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b124|biu/cache_ctrl_logic/reg1_b76  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [124],\biu/cache_ctrl_logic/l1i_pa [76]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pa_temp [124],\biu/cache_ctrl_logic/pa_temp [76]}),
    .mi({\biu/cache_ctrl_logic/pa_temp [124],\biu/cache_ctrl_logic/pa_temp [76]}),
    .sr(rst_pad),
    .f({_al_u4438_o,_al_u4750_o}),
    .q({\biu/cache_ctrl_logic/l1i_pa [124],\biu/cache_ctrl_logic/l1i_pa [76]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b12|biu/cache_ctrl_logic/reg1_b7  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [12],\biu/cache_ctrl_logic/pa_temp [7]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [12],\biu/cache_ctrl_logic/l1i_pa [7]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b13|biu/cache_ctrl_logic/reg1_b63  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [13],\biu/cache_ctrl_logic/pa_temp [63]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [13],\biu/cache_ctrl_logic/l1i_pa [63]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b14|biu/cache_ctrl_logic/reg1_b62  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [14],\biu/cache_ctrl_logic/pa_temp [62]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [14],\biu/cache_ctrl_logic/l1i_pa [62]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b15|biu/cache_ctrl_logic/reg1_b61  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [15],\biu/cache_ctrl_logic/pa_temp [61]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [15],\biu/cache_ctrl_logic/l1i_pa [61]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b16|biu/cache_ctrl_logic/reg1_b60  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [16],\biu/cache_ctrl_logic/pa_temp [60]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [16],\biu/cache_ctrl_logic/l1i_pa [60]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b17|biu/cache_ctrl_logic/reg1_b6  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [17],\biu/cache_ctrl_logic/pa_temp [6]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [17],\biu/cache_ctrl_logic/l1i_pa [6]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b18|biu/cache_ctrl_logic/reg1_b59  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [18],\biu/cache_ctrl_logic/pa_temp [59]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [18],\biu/cache_ctrl_logic/l1i_pa [59]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b19|biu/cache_ctrl_logic/reg1_b58  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [19],\biu/cache_ctrl_logic/pa_temp [58]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [19],\biu/cache_ctrl_logic/l1i_pa [58]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b20|biu/cache_ctrl_logic/reg1_b57  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [20],\biu/cache_ctrl_logic/pa_temp [57]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [20],\biu/cache_ctrl_logic/l1i_pa [57]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b21|biu/cache_ctrl_logic/reg1_b56  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [21],\biu/cache_ctrl_logic/pa_temp [56]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [21],\biu/cache_ctrl_logic/l1i_pa [56]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b22|biu/cache_ctrl_logic/reg1_b55  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [22],\biu/cache_ctrl_logic/pa_temp [55]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [22],\biu/cache_ctrl_logic/l1i_pa [55]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b23|biu/cache_ctrl_logic/reg1_b54  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [23],\biu/cache_ctrl_logic/pa_temp [54]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [23],\biu/cache_ctrl_logic/l1i_pa [54]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b24|biu/cache_ctrl_logic/reg1_b53  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [24],\biu/cache_ctrl_logic/pa_temp [53]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [24],\biu/cache_ctrl_logic/l1i_pa [53]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b25|biu/cache_ctrl_logic/reg1_b52  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [25],\biu/cache_ctrl_logic/pa_temp [52]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [25],\biu/cache_ctrl_logic/l1i_pa [52]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b26|biu/cache_ctrl_logic/reg1_b51  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [26],\biu/cache_ctrl_logic/pa_temp [51]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [26],\biu/cache_ctrl_logic/l1i_pa [51]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b27|biu/cache_ctrl_logic/reg1_b50  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [27],\biu/cache_ctrl_logic/pa_temp [50]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [27],\biu/cache_ctrl_logic/l1i_pa [50]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b28|biu/cache_ctrl_logic/reg1_b5  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [28],\biu/cache_ctrl_logic/pa_temp [5]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [28],\biu/cache_ctrl_logic/l1i_pa [5]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b29|biu/cache_ctrl_logic/reg1_b49  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [29],\biu/cache_ctrl_logic/pa_temp [49]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [29],\biu/cache_ctrl_logic/l1i_pa [49]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b3  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({open_n78836,\biu/cache_ctrl_logic/pa_temp [3]}),
    .sr(rst_pad),
    .q({open_n78842,\biu/cache_ctrl_logic/l1i_pa [3]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b30|biu/cache_ctrl_logic/reg1_b48  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [30],\biu/cache_ctrl_logic/pa_temp [48]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [30],\biu/cache_ctrl_logic/l1i_pa [48]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b31|biu/cache_ctrl_logic/reg1_b47  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [31],\biu/cache_ctrl_logic/pa_temp [47]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [31],\biu/cache_ctrl_logic/l1i_pa [47]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b32|biu/cache_ctrl_logic/reg1_b46  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [32],\biu/cache_ctrl_logic/pa_temp [46]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [32],\biu/cache_ctrl_logic/l1i_pa [46]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b33|biu/cache_ctrl_logic/reg1_b45  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [33],\biu/cache_ctrl_logic/pa_temp [45]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [33],\biu/cache_ctrl_logic/l1i_pa [45]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b34|biu/cache_ctrl_logic/reg1_b44  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [34],\biu/cache_ctrl_logic/pa_temp [44]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [34],\biu/cache_ctrl_logic/l1i_pa [44]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b35|biu/cache_ctrl_logic/reg1_b43  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [35],\biu/cache_ctrl_logic/pa_temp [43]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [35],\biu/cache_ctrl_logic/l1i_pa [43]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b36|biu/cache_ctrl_logic/reg1_b42  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [36],\biu/cache_ctrl_logic/pa_temp [42]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [36],\biu/cache_ctrl_logic/l1i_pa [42]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b37|biu/cache_ctrl_logic/reg1_b41  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [37],\biu/cache_ctrl_logic/pa_temp [41]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [37],\biu/cache_ctrl_logic/l1i_pa [41]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b38|biu/cache_ctrl_logic/reg1_b40  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [38],\biu/cache_ctrl_logic/pa_temp [40]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [38],\biu/cache_ctrl_logic/l1i_pa [40]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b39|biu/cache_ctrl_logic/reg1_b4  (
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [39],\biu/cache_ctrl_logic/pa_temp [4]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1i_pa [39],\biu/cache_ctrl_logic/l1i_pa [4]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg1_b67|biu/cache_ctrl_logic/reg1_b70  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pa [67],\biu/cache_ctrl_logic/l1i_pa [70]}),
    .ce(\biu/cache_ctrl_logic/n140 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pa_temp [67],\biu/cache_ctrl_logic/pa_temp [70]}),
    .mi({\biu/cache_ctrl_logic/pa_temp [67],\biu/cache_ctrl_logic/pa_temp [70]}),
    .sr(rst_pad),
    .f({_al_u4642_o,_al_u4444_o}),
    .q({\biu/cache_ctrl_logic/l1i_pa [67],\biu/cache_ctrl_logic/l1i_pa [70]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg2_b0|biu/cache_ctrl_logic/reg2_b61  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [0],\biu/cache_ctrl_logic/l1i_pte [61]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pte_temp [0],\biu/cache_ctrl_logic/pte_temp [61]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [0],\biu/cache_ctrl_logic/pte_temp [61]}),
    .sr(rst_pad),
    .f({_al_u4796_o,_al_u5684_o}),
    .q({\biu/cache_ctrl_logic/l1i_pte [0],\biu/cache_ctrl_logic/l1i_pte [61]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg2_b23|biu/cache_ctrl_logic/reg2_b54  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [23],\biu/cache_ctrl_logic/l1i_pte [54]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pte_temp [23],\biu/cache_ctrl_logic/pte_temp [54]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [23],\biu/cache_ctrl_logic/pte_temp [54]}),
    .sr(rst_pad),
    .f({_al_u5118_o,_al_u5712_o}),
    .q({\biu/cache_ctrl_logic/l1i_pte [23],\biu/cache_ctrl_logic/l1i_pte [54]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg2_b25|biu/cache_ctrl_logic/reg2_b53  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [25],\biu/cache_ctrl_logic/l1i_pte [53]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pte_temp [25],\biu/cache_ctrl_logic/pte_temp [53]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [25],\biu/cache_ctrl_logic/pte_temp [53]}),
    .sr(rst_pad),
    .f({_al_u5828_o,_al_u5716_o}),
    .q({\biu/cache_ctrl_logic/l1i_pte [25],\biu/cache_ctrl_logic/l1i_pte [53]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg2_b26|biu/cache_ctrl_logic/reg2_b51  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [26],\biu/cache_ctrl_logic/l1i_pte [51]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pte_temp [26],\biu/cache_ctrl_logic/pte_temp [51]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [26],\biu/cache_ctrl_logic/pte_temp [51]}),
    .sr(rst_pad),
    .f({_al_u5824_o,_al_u5724_o}),
    .q({\biu/cache_ctrl_logic/l1i_pte [26],\biu/cache_ctrl_logic/l1i_pte [51]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg2_b32|biu/cache_ctrl_logic/reg2_b44  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [32],\biu/cache_ctrl_logic/l1i_pte [44]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pte_temp [32],\biu/cache_ctrl_logic/pte_temp [44]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [32],\biu/cache_ctrl_logic/pte_temp [44]}),
    .sr(rst_pad),
    .f({_al_u5800_o,_al_u5752_o}),
    .q({\biu/cache_ctrl_logic/l1i_pte [32],\biu/cache_ctrl_logic/l1i_pte [44]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg2_b35|biu/cache_ctrl_logic/reg2_b40  (
    .a({_al_u3945_o,_al_u3945_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [35],\biu/cache_ctrl_logic/l1i_pte [40]}),
    .ce(\biu/cache_ctrl_logic/n135 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/pte_temp [35],\biu/cache_ctrl_logic/pte_temp [40]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [35],\biu/cache_ctrl_logic/pte_temp [40]}),
    .sr(rst_pad),
    .f({_al_u5788_o,_al_u5768_o}),
    .q({\biu/cache_ctrl_logic/l1i_pte [35],\biu/cache_ctrl_logic/l1i_pte [40]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b15|biu/cache_ctrl_logic/reg3_b25  (
    .a({\biu/cache_ctrl_logic/l1i_va [15],\biu/cache_ctrl_logic/l1i_va [13]}),
    .b({\biu/cache_ctrl_logic/l1i_va [25],\biu/cache_ctrl_logic/l1i_va [25]}),
    .c({addr_ex[15],addr_ex[13]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[25],addr_ex[25]}),
    .mi({addr_ex[15],addr_ex[25]}),
    .sr(rst_pad),
    .f({_al_u6374_o,_al_u6367_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [15],\biu/cache_ctrl_logic/l1d_va [25]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1100010011110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b18|biu/cache_ctrl_logic/reg3_b24  (
    .a({\biu/cache_ctrl_logic/l1i_va [18],\biu/cache_ctrl_logic/l1i_va [18]}),
    .b({\biu/cache_ctrl_logic/l1i_va [32],\biu/cache_ctrl_logic/l1i_va [24]}),
    .c({addr_ex[18],addr_ex[18]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[32],addr_ex[24]}),
    .mi({addr_ex[18],addr_ex[24]}),
    .sr(rst_pad),
    .f({_al_u6407_o,_al_u6368_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [18],\biu/cache_ctrl_logic/l1d_va [24]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100110001),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b33|biu/cache_ctrl_logic/reg3_b13  (
    .a({open_n79222,\biu/cache_ctrl_logic/l1i_va [13]}),
    .b({\biu/cache_ctrl_logic/l1i_va [33],\biu/cache_ctrl_logic/l1i_va [15]}),
    .c({addr_ex[33],addr_ex[13]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6372_o,addr_ex[15]}),
    .mi({addr_ex[33],addr_ex[13]}),
    .sr(rst_pad),
    .f({_al_u6373_o,_al_u6372_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [33],\biu/cache_ctrl_logic/l1d_va [13]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b35|biu/cache_ctrl_logic/reg3_b23  (
    .a({\biu/cache_ctrl_logic/l1d_va [23],\biu/cache_ctrl_logic/l1i_va [23]}),
    .b({\biu/cache_ctrl_logic/l1d_va [35],\biu/cache_ctrl_logic/l1i_va [53]}),
    .c({addr_ex[23],addr_ex[23]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[35],addr_ex[53]}),
    .mi({addr_ex[35],addr_ex[23]}),
    .sr(rst_pad),
    .f({_al_u6279_o,_al_u6376_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [35],\biu/cache_ctrl_logic/l1d_va [23]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b36|biu/cache_ctrl_logic/reg3_b26  (
    .a({\biu/cache_ctrl_logic/l1i_va [36],\biu/cache_ctrl_logic/l1i_va [26]}),
    .b({\biu/cache_ctrl_logic/l1i_va [40],\biu/cache_ctrl_logic/l1i_va [36]}),
    .c({addr_ex[36],addr_ex[26]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[40],addr_ex[36]}),
    .mi({addr_ex[36],addr_ex[26]}),
    .sr(rst_pad),
    .f({_al_u6406_o,_al_u6413_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [36],\biu/cache_ctrl_logic/l1d_va [26]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b39|biu/cache_ctrl_logic/reg3_b31  (
    .a({\biu/cache_ctrl_logic/l1d_va [31],\biu/cache_ctrl_logic/l1i_va [31]}),
    .b({\biu/cache_ctrl_logic/l1d_va [39],\biu/cache_ctrl_logic/l1i_va [55]}),
    .c({addr_ex[31],addr_ex[31]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[39],addr_ex[55]}),
    .mi({addr_ex[39],addr_ex[31]}),
    .sr(rst_pad),
    .f({_al_u6267_o,_al_u6398_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [39],\biu/cache_ctrl_logic/l1d_va [31]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b43|biu/cache_ctrl_logic/reg3_b45  (
    .a({\biu/cache_ctrl_logic/l1i_va [43],\biu/cache_ctrl_logic/l1i_va [45]}),
    .b({\biu/cache_ctrl_logic/l1i_va [45],\biu/cache_ctrl_logic/l1i_va [58]}),
    .c({addr_ex[43],addr_ex[45]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[45],addr_ex[58]}),
    .mi({addr_ex[43],addr_ex[45]}),
    .sr(rst_pad),
    .f({_al_u6381_o,_al_u6385_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [43],\biu/cache_ctrl_logic/l1d_va [45]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C@A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010010100101),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b47|biu/cache_ctrl_logic/reg3_b53  (
    .a({open_n79304,\biu/cache_ctrl_logic/l1d_va [47]}),
    .b({\biu/cache_ctrl_logic/l1i_va [47],\biu/cache_ctrl_logic/l1d_va [53]}),
    .c({addr_ex[47],addr_ex[47]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6374_o,addr_ex[53]}),
    .mi({addr_ex[47],addr_ex[53]}),
    .sr(rst_pad),
    .f({_al_u6375_o,_al_u6295_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [47],\biu/cache_ctrl_logic/l1d_va [53]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b56|biu/cache_ctrl_logic/reg3_b54  (
    .a({\biu/cache_ctrl_logic/l1i_va [29],\biu/cache_ctrl_logic/l1i_va [54]}),
    .b({\biu/cache_ctrl_logic/l1i_va [56],\biu/cache_ctrl_logic/l1i_va [56]}),
    .c({addr_ex[29],addr_ex[54]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[56],addr_ex[56]}),
    .mi({addr_ex[56],addr_ex[54]}),
    .sr(rst_pad),
    .f({_al_u6401_o,_al_u6386_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [56],\biu/cache_ctrl_logic/l1d_va [54]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b57|biu/cache_ctrl_logic/reg3_b42  (
    .a({open_n79335,\biu/cache_ctrl_logic/l1i_va [42]}),
    .b({\biu/cache_ctrl_logic/l1i_va [57],\biu/cache_ctrl_logic/l1i_va [43]}),
    .c({addr_ex[57],addr_ex[42]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({_al_u6379_o,addr_ex[43]}),
    .mi({addr_ex[57],addr_ex[42]}),
    .sr(rst_pad),
    .f({_al_u6380_o,_al_u6379_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [57],\biu/cache_ctrl_logic/l1d_va [42]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b61|biu/cache_ctrl_logic/reg3_b21  (
    .a({\biu/cache_ctrl_logic/l1d_va [21],\biu/cache_ctrl_logic/l1i_va [21]}),
    .b({\biu/cache_ctrl_logic/l1d_va [61],\biu/cache_ctrl_logic/l1i_va [39]}),
    .c({addr_ex[21],addr_ex[21]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[61],addr_ex[39]}),
    .mi({addr_ex[61],addr_ex[21]}),
    .sr(rst_pad),
    .f({_al_u6269_o,_al_u6390_o}),
    .q({\biu/cache_ctrl_logic/l1d_va [61],\biu/cache_ctrl_logic/l1d_va [21]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b1100010011110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg3_b63|biu/cache_ctrl_logic/reg3_b62  (
    .a({\biu/cache_ctrl_logic/l1d_va [62],\biu/cache_ctrl_logic/l1i_va [62]}),
    .b({\biu/cache_ctrl_logic/l1d_va [63],\biu/cache_ctrl_logic/l1i_va [63]}),
    .c({addr_ex[62],addr_ex[62]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({addr_ex[63],addr_ex[63]}),
    .mi(addr_ex[63:62]),
    .sr(rst_pad),
    .f({_al_u6262_o,_al_u6370_o}),
    .q(\biu/cache_ctrl_logic/l1d_va [63:62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b102|biu/cache_ctrl_logic/reg4_b33  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [102],\biu/cache_ctrl_logic/pa_temp [33]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [102],\biu/cache_ctrl_logic/l1d_pa [33]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b103|biu/cache_ctrl_logic/reg4_b31  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [103],\biu/cache_ctrl_logic/pa_temp [31]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [103],\biu/cache_ctrl_logic/l1d_pa [31]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b107|biu/cache_ctrl_logic/reg4_b30  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [107],\biu/cache_ctrl_logic/pa_temp [30]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [107],\biu/cache_ctrl_logic/l1d_pa [30]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b108|biu/cache_ctrl_logic/reg4_b29  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [108],\biu/cache_ctrl_logic/pa_temp [29]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [108],\biu/cache_ctrl_logic/l1d_pa [29]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b10|biu/cache_ctrl_logic/reg4_b7  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [10],\biu/cache_ctrl_logic/pa_temp [7]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [10],\biu/cache_ctrl_logic/l1d_pa [7]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b110|biu/cache_ctrl_logic/reg4_b28  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [110],\biu/cache_ctrl_logic/pa_temp [28]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [110],\biu/cache_ctrl_logic/l1d_pa [28]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b111|biu/cache_ctrl_logic/reg4_b27  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [111],\biu/cache_ctrl_logic/pa_temp [27]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [111],\biu/cache_ctrl_logic/l1d_pa [27]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b112|biu/cache_ctrl_logic/reg4_b26  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [112],\biu/cache_ctrl_logic/pa_temp [26]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [112],\biu/cache_ctrl_logic/l1d_pa [26]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b113|biu/cache_ctrl_logic/reg4_b25  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [113],\biu/cache_ctrl_logic/pa_temp [25]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [113],\biu/cache_ctrl_logic/l1d_pa [25]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b115|biu/cache_ctrl_logic/reg4_b24  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [115],\biu/cache_ctrl_logic/pa_temp [24]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [115],\biu/cache_ctrl_logic/l1d_pa [24]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b118|biu/cache_ctrl_logic/reg4_b23  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [118],\biu/cache_ctrl_logic/pa_temp [23]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [118],\biu/cache_ctrl_logic/l1d_pa [23]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b119|biu/cache_ctrl_logic/reg4_b22  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [119],\biu/cache_ctrl_logic/pa_temp [22]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [119],\biu/cache_ctrl_logic/l1d_pa [22]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b11|biu/cache_ctrl_logic/reg4_b21  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [11],\biu/cache_ctrl_logic/pa_temp [21]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [11],\biu/cache_ctrl_logic/l1d_pa [21]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b120|biu/cache_ctrl_logic/reg4_b20  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [120],\biu/cache_ctrl_logic/pa_temp [20]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [120],\biu/cache_ctrl_logic/l1d_pa [20]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b121|biu/cache_ctrl_logic/reg4_b2  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [121],\biu/cache_ctrl_logic/pa_temp [2]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [121],\biu/cache_ctrl_logic/l1d_pa [2]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b122|biu/cache_ctrl_logic/reg4_b19  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [122],\biu/cache_ctrl_logic/pa_temp [19]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [122],\biu/cache_ctrl_logic/l1d_pa [19]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b123|biu/cache_ctrl_logic/reg4_b18  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [123],\biu/cache_ctrl_logic/pa_temp [18]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [123],\biu/cache_ctrl_logic/l1d_pa [18]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b125|biu/cache_ctrl_logic/reg4_b17  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [125],\biu/cache_ctrl_logic/pa_temp [17]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [125],\biu/cache_ctrl_logic/l1d_pa [17]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b126|biu/cache_ctrl_logic/reg4_b16  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [126],\biu/cache_ctrl_logic/pa_temp [16]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [126],\biu/cache_ctrl_logic/l1d_pa [16]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b127|biu/cache_ctrl_logic/reg4_b15  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [127],\biu/cache_ctrl_logic/pa_temp [15]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [127],\biu/cache_ctrl_logic/l1d_pa [15]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b12|biu/cache_ctrl_logic/reg4_b14  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [12],\biu/cache_ctrl_logic/pa_temp [14]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [12],\biu/cache_ctrl_logic/l1d_pa [14]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b32|biu/cache_ctrl_logic/reg4_b34  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [32],\biu/cache_ctrl_logic/pa_temp [34]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [32],\biu/cache_ctrl_logic/l1d_pa [34]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b35|biu/cache_ctrl_logic/reg4_b37  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [35],\biu/cache_ctrl_logic/pa_temp [37]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [35],\biu/cache_ctrl_logic/l1d_pa [37]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b36|biu/cache_ctrl_logic/reg4_b38  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [36],\biu/cache_ctrl_logic/pa_temp [38]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [36],\biu/cache_ctrl_logic/l1d_pa [38]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b39|biu/cache_ctrl_logic/reg4_b41  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [39],\biu/cache_ctrl_logic/pa_temp [41]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [39],\biu/cache_ctrl_logic/l1d_pa [41]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b3|biu/cache_ctrl_logic/reg4_b5  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [3],\biu/cache_ctrl_logic/pa_temp [5]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [3],\biu/cache_ctrl_logic/l1d_pa [5]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b40|biu/cache_ctrl_logic/reg4_b42  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [40],\biu/cache_ctrl_logic/pa_temp [42]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [40],\biu/cache_ctrl_logic/l1d_pa [42]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b43|biu/cache_ctrl_logic/reg4_b45  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [43],\biu/cache_ctrl_logic/pa_temp [45]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [43],\biu/cache_ctrl_logic/l1d_pa [45]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b44|biu/cache_ctrl_logic/reg4_b46  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [44],\biu/cache_ctrl_logic/pa_temp [46]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [44],\biu/cache_ctrl_logic/l1d_pa [46]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b47|biu/cache_ctrl_logic/reg4_b49  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [47],\biu/cache_ctrl_logic/pa_temp [49]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [47],\biu/cache_ctrl_logic/l1d_pa [49]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b48|biu/cache_ctrl_logic/reg4_b50  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [48],\biu/cache_ctrl_logic/pa_temp [50]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [48],\biu/cache_ctrl_logic/l1d_pa [50]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b4|biu/cache_ctrl_logic/reg4_b6  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [4],\biu/cache_ctrl_logic/pa_temp [6]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [4],\biu/cache_ctrl_logic/l1d_pa [6]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b51|biu/cache_ctrl_logic/reg4_b53  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [51],\biu/cache_ctrl_logic/pa_temp [53]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [51],\biu/cache_ctrl_logic/l1d_pa [53]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b52|biu/cache_ctrl_logic/reg4_b54  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [52],\biu/cache_ctrl_logic/pa_temp [54]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [52],\biu/cache_ctrl_logic/l1d_pa [54]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b55|biu/cache_ctrl_logic/reg4_b57  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [55],\biu/cache_ctrl_logic/pa_temp [57]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [55],\biu/cache_ctrl_logic/l1d_pa [57]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b56|biu/cache_ctrl_logic/reg4_b58  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [56],\biu/cache_ctrl_logic/pa_temp [58]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [56],\biu/cache_ctrl_logic/l1d_pa [58]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b59|biu/cache_ctrl_logic/reg4_b61  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [59],\biu/cache_ctrl_logic/pa_temp [61]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [59],\biu/cache_ctrl_logic/l1d_pa [61]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b60|biu/cache_ctrl_logic/reg4_b62  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [60],\biu/cache_ctrl_logic/pa_temp [62]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [60],\biu/cache_ctrl_logic/l1d_pa [62]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b63  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({open_n80343,\biu/cache_ctrl_logic/pa_temp [63]}),
    .sr(rst_pad),
    .q({open_n80349,\biu/cache_ctrl_logic/l1d_pa [63]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b65|biu/cache_ctrl_logic/reg4_b13  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [65],\biu/cache_ctrl_logic/pa_temp [13]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [65],\biu/cache_ctrl_logic/l1d_pa [13]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b66|biu/cache_ctrl_logic/reg5_b9  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [66],\biu/cache_ctrl_logic/pte_temp [9]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [66],\biu/cache_ctrl_logic/l1d_pte [9]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b69|biu/cache_ctrl_logic/reg5_b8  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [69],\biu/cache_ctrl_logic/pte_temp [8]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [69],\biu/cache_ctrl_logic/l1d_pte [8]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b71|biu/cache_ctrl_logic/reg5_b57  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [71],\biu/cache_ctrl_logic/pte_temp [57]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [71],\biu/cache_ctrl_logic/l1d_pte [57]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b72|biu/cache_ctrl_logic/reg5_b55  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [72],\biu/cache_ctrl_logic/pte_temp [55]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [72],\biu/cache_ctrl_logic/l1d_pte [55]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b74|biu/cache_ctrl_logic/reg5_b50  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [74],\biu/cache_ctrl_logic/pte_temp [50]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [74],\biu/cache_ctrl_logic/l1d_pte [50]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b78|biu/cache_ctrl_logic/reg5_b47  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [78],\biu/cache_ctrl_logic/pte_temp [47]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [78],\biu/cache_ctrl_logic/l1d_pte [47]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b79|biu/cache_ctrl_logic/reg5_b45  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [79],\biu/cache_ctrl_logic/pte_temp [45]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [79],\biu/cache_ctrl_logic/l1d_pte [45]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b82|biu/cache_ctrl_logic/reg5_b31  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [82],\biu/cache_ctrl_logic/pte_temp [31]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [82],\biu/cache_ctrl_logic/l1d_pte [31]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b84|biu/cache_ctrl_logic/reg5_b28  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [84],\biu/cache_ctrl_logic/pte_temp [28]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [84],\biu/cache_ctrl_logic/l1d_pte [28]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b86|biu/cache_ctrl_logic/reg5_b21  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [86],\biu/cache_ctrl_logic/pte_temp [21]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [86],\biu/cache_ctrl_logic/l1d_pte [21]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b87|biu/cache_ctrl_logic/reg5_b18  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [87],\biu/cache_ctrl_logic/pte_temp [18]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [87],\biu/cache_ctrl_logic/l1d_pte [18]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b89|biu/cache_ctrl_logic/reg5_b16  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [89],\biu/cache_ctrl_logic/pte_temp [16]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [89],\biu/cache_ctrl_logic/l1d_pte [16]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b8|biu/cache_ctrl_logic/reg4_b9  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [8],\biu/cache_ctrl_logic/pa_temp [9]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [8],\biu/cache_ctrl_logic/l1d_pa [9]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b90|biu/cache_ctrl_logic/reg5_b14  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [90],\biu/cache_ctrl_logic/pte_temp [14]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [90],\biu/cache_ctrl_logic/l1d_pte [14]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b91|biu/cache_ctrl_logic/reg5_b11  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [91],\biu/cache_ctrl_logic/pte_temp [11]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [91],\biu/cache_ctrl_logic/l1d_pte [11]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b92|biu/cache_ctrl_logic/reg4_b99  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [92],\biu/cache_ctrl_logic/pa_temp [99]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [92],\biu/cache_ctrl_logic/l1d_pa [99]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b95|biu/cache_ctrl_logic/reg4_b98  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({\biu/cache_ctrl_logic/pa_temp [95],\biu/cache_ctrl_logic/pa_temp [98]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/l1d_pa [95],\biu/cache_ctrl_logic/l1d_pa [98]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg4_b97  (
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .mi({open_n80815,\biu/cache_ctrl_logic/pa_temp [97]}),
    .sr(rst_pad),
    .q({open_n80832,\biu/cache_ctrl_logic/l1d_pa [97]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b10|biu/cache_ctrl_logic/reg5_b62  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [10],\biu/cache_ctrl_logic/l1i_pte [62]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [10],\biu/cache_ctrl_logic/l1d_pte [62]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [10],\biu/cache_ctrl_logic/pte_temp [62]}),
    .sr(rst_pad),
    .f({_al_u4860_o,_al_u5680_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [10],\biu/cache_ctrl_logic/l1d_pte [62]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b12|biu/cache_ctrl_logic/reg5_b60  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [12],\biu/cache_ctrl_logic/l1i_pte [60]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [12],\biu/cache_ctrl_logic/l1d_pte [60]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [12],\biu/cache_ctrl_logic/pte_temp [60]}),
    .sr(rst_pad),
    .f({_al_u4852_o,_al_u5688_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [12],\biu/cache_ctrl_logic/l1d_pte [60]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b13|biu/cache_ctrl_logic/reg5_b6  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [13],\biu/cache_ctrl_logic/l1i_pte [6]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [13],\biu/cache_ctrl_logic/l1d_pte [6]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [13],\biu/cache_ctrl_logic/pte_temp [6]}),
    .sr(rst_pad),
    .f({_al_u4848_o,_al_u4772_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [13],\biu/cache_ctrl_logic/l1d_pte [6]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b15|biu/cache_ctrl_logic/reg5_b59  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [15],\biu/cache_ctrl_logic/l1i_pte [59]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [15],\biu/cache_ctrl_logic/l1d_pte [59]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [15],\biu/cache_ctrl_logic/pte_temp [59]}),
    .sr(rst_pad),
    .f({_al_u4840_o,_al_u5692_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [15],\biu/cache_ctrl_logic/l1d_pte [59]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b17|biu/cache_ctrl_logic/reg5_b58  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [17],\biu/cache_ctrl_logic/l1i_pte [58]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [17],\biu/cache_ctrl_logic/l1d_pte [58]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [17],\biu/cache_ctrl_logic/pte_temp [58]}),
    .sr(rst_pad),
    .f({_al_u5110_o,_al_u5696_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [17],\biu/cache_ctrl_logic/l1d_pte [58]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b19|biu/cache_ctrl_logic/reg5_b56  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [19],\biu/cache_ctrl_logic/l1i_pte [56]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [19],\biu/cache_ctrl_logic/l1d_pte [56]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [19],\biu/cache_ctrl_logic/pte_temp [56]}),
    .sr(rst_pad),
    .f({_al_u5134_o,_al_u5704_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [19],\biu/cache_ctrl_logic/l1d_pte [56]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~B*~(D*C)))"),
    //.LUTF1("(A*~(~B*~(D*C)))"),
    //.LUTG0("(A*~(~B*~(D*C)))"),
    //.LUTG1("(A*~(~B*~(D*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010100010001000),
    .INIT_LUTF1(16'b1010100010001000),
    .INIT_LUTG0(16'b1010100010001000),
    .INIT_LUTG1(16'b1010100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b1|biu/cache_ctrl_logic/reg5_b3  (
    .a({read,read}),
    .b({\biu/cache_ctrl_logic/l1d_pte [1],\biu/cache_ctrl_logic/l1i_pte [1]}),
    .c({\biu/cache_ctrl_logic/l1d_pte [3],\biu/cache_ctrl_logic/l1d_pte [3]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({mxr,mxr}),
    .mi({\biu/cache_ctrl_logic/pte_temp [1],\biu/cache_ctrl_logic/pte_temp [3]}),
    .sr(rst_pad),
    .f({\biu/cache_ctrl_logic/n34 ,\biu/cache_ctrl_logic/n42 }),
    .q({\biu/cache_ctrl_logic/l1d_pte [1],\biu/cache_ctrl_logic/l1d_pte [3]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b20|biu/cache_ctrl_logic/reg5_b52  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [20],\biu/cache_ctrl_logic/l1i_pte [52]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [20],\biu/cache_ctrl_logic/l1d_pte [52]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [20],\biu/cache_ctrl_logic/pte_temp [52]}),
    .sr(rst_pad),
    .f({_al_u5130_o,_al_u5720_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [20],\biu/cache_ctrl_logic/l1d_pte [52]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b22|biu/cache_ctrl_logic/reg5_b5  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [22],\biu/cache_ctrl_logic/l1i_pte [5]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [22],\biu/cache_ctrl_logic/l1d_pte [5]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [22],\biu/cache_ctrl_logic/pte_temp [5]}),
    .sr(rst_pad),
    .f({_al_u5122_o,_al_u4776_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [22],\biu/cache_ctrl_logic/l1d_pte [5]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b24|biu/cache_ctrl_logic/reg5_b49  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [24],\biu/cache_ctrl_logic/l1i_pte [49]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [24],\biu/cache_ctrl_logic/l1d_pte [49]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [24],\biu/cache_ctrl_logic/pte_temp [49]}),
    .sr(rst_pad),
    .f({_al_u5832_o,_al_u5732_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [24],\biu/cache_ctrl_logic/l1d_pte [49]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b27|biu/cache_ctrl_logic/reg5_b48  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [27],\biu/cache_ctrl_logic/l1i_pte [48]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [27],\biu/cache_ctrl_logic/l1d_pte [48]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [27],\biu/cache_ctrl_logic/pte_temp [48]}),
    .sr(rst_pad),
    .f({_al_u5820_o,_al_u5736_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [27],\biu/cache_ctrl_logic/l1d_pte [48]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b29|biu/cache_ctrl_logic/reg5_b46  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [29],\biu/cache_ctrl_logic/l1i_pte [46]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [29],\biu/cache_ctrl_logic/l1d_pte [46]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [29],\biu/cache_ctrl_logic/pte_temp [46]}),
    .sr(rst_pad),
    .f({_al_u5812_o,_al_u5744_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [29],\biu/cache_ctrl_logic/l1d_pte [46]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b30|biu/cache_ctrl_logic/reg5_b43  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [30],\biu/cache_ctrl_logic/l1i_pte [43]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [30],\biu/cache_ctrl_logic/l1d_pte [43]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [30],\biu/cache_ctrl_logic/pte_temp [43]}),
    .sr(rst_pad),
    .f({_al_u5808_o,_al_u5756_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [30],\biu/cache_ctrl_logic/l1d_pte [43]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b33|biu/cache_ctrl_logic/reg5_b42  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [33],\biu/cache_ctrl_logic/l1i_pte [42]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [33],\biu/cache_ctrl_logic/l1d_pte [42]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [33],\biu/cache_ctrl_logic/pte_temp [42]}),
    .sr(rst_pad),
    .f({_al_u5796_o,_al_u5760_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [33],\biu/cache_ctrl_logic/l1d_pte [42]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*B)*~(D*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(C*B)*~(D*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001010100111111),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b0001010100111111),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b34|biu/cache_ctrl_logic/reg5_b41  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [34],\biu/cache_ctrl_logic/l1i_pte [41]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [34],\biu/cache_ctrl_logic/l1d_pte [41]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [34],\biu/cache_ctrl_logic/pte_temp [41]}),
    .sr(rst_pad),
    .f({_al_u5792_o,_al_u5764_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [34],\biu/cache_ctrl_logic/l1d_pte [41]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg5_b37|biu/cache_ctrl_logic/reg5_b39  (
    .a({_al_u3947_o,_al_u3947_o}),
    .b({_al_u3950_o,_al_u3950_o}),
    .c({\biu/cache_ctrl_logic/l1i_pte [37],\biu/cache_ctrl_logic/l1i_pte [39]}),
    .ce(\biu/cache_ctrl_logic/n149 ),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_pte [37],\biu/cache_ctrl_logic/l1d_pte [39]}),
    .mi({\biu/cache_ctrl_logic/pte_temp [37],\biu/cache_ctrl_logic/pte_temp [39]}),
    .sr(rst_pad),
    .f({_al_u5780_o,_al_u5772_o}),
    .q({\biu/cache_ctrl_logic/l1d_pte [37],\biu/cache_ctrl_logic/l1d_pte [39]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000101100000000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1000101100000000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b0|biu/bus_unit/mmu/reg1_b0  (
    .a({open_n81077,_al_u2914_o}),
    .b({\biu/paddress [0],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [0],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [0]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [0],\biu/paddress [0]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b100|biu/cache_ctrl_logic/reg6_b75  (
    .a({_al_u2698_o,open_n81100}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [8]}),
    .c({\biu/paddress [100],\biu/paddress [75]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [34],_al_u2705_o}),
    .mi({\biu/paddress [100],\biu/paddress [75]}),
    .sr(rst_pad),
    .f({_al_u3101_o,haddr_pad[11]}),
    .q({\biu/cache_ctrl_logic/pa_temp [100],\biu/cache_ctrl_logic/pa_temp [75]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b101|biu/cache_ctrl_logic/reg6_b74  (
    .a({_al_u2698_o,open_n81114}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [7]}),
    .c({\biu/paddress [101],\biu/paddress [74]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [35],_al_u2705_o}),
    .mi({\biu/paddress [101],\biu/paddress [74]}),
    .sr(rst_pad),
    .f({_al_u3098_o,haddr_pad[10]}),
    .q({\biu/cache_ctrl_logic/pa_temp [101],\biu/cache_ctrl_logic/pa_temp [74]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b102|biu/cache_ctrl_logic/reg6_b73  (
    .a({_al_u2698_o,open_n81128}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [6]}),
    .c({\biu/paddress [102],\biu/paddress [73]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [36],_al_u2705_o}),
    .mi({\biu/paddress [102],\biu/paddress [73]}),
    .sr(rst_pad),
    .f({_al_u3095_o,haddr_pad[9]}),
    .q({\biu/cache_ctrl_logic/pa_temp [102],\biu/cache_ctrl_logic/pa_temp [73]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b103|biu/cache_ctrl_logic/reg6_b72  (
    .a({_al_u2698_o,open_n81146}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [5]}),
    .c({\biu/paddress [103],\biu/paddress [72]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [37],_al_u2705_o}),
    .mi({\biu/paddress [103],\biu/paddress [72]}),
    .sr(rst_pad),
    .f({_al_u3092_o,haddr_pad[8]}),
    .q({\biu/cache_ctrl_logic/pa_temp [103],\biu/cache_ctrl_logic/pa_temp [72]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b104|biu/cache_ctrl_logic/reg6_b71  (
    .a({_al_u2698_o,open_n81164}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [4]}),
    .c({\biu/paddress [104],\biu/paddress [71]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [38],_al_u2705_o}),
    .mi({\biu/paddress [104],\biu/paddress [71]}),
    .sr(rst_pad),
    .f({_al_u3089_o,haddr_pad[7]}),
    .q({\biu/cache_ctrl_logic/pa_temp [104],\biu/cache_ctrl_logic/pa_temp [71]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b105|biu/cache_ctrl_logic/reg6_b70  (
    .a({_al_u2698_o,open_n81178}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [3]}),
    .c({\biu/paddress [105],\biu/paddress [70]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [39],_al_u2705_o}),
    .mi({\biu/paddress [105],\biu/paddress [70]}),
    .sr(rst_pad),
    .f({_al_u3086_o,haddr_pad[6]}),
    .q({\biu/cache_ctrl_logic/pa_temp [105],\biu/cache_ctrl_logic/pa_temp [70]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b106|biu/cache_ctrl_logic/reg6_b69  (
    .a({_al_u2698_o,open_n81192}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [2]}),
    .c({\biu/paddress [106],\biu/paddress [69]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [40],_al_u2705_o}),
    .mi({\biu/paddress [106],\biu/paddress [69]}),
    .sr(rst_pad),
    .f({_al_u3083_o,haddr_pad[5]}),
    .q({\biu/cache_ctrl_logic/pa_temp [106],\biu/cache_ctrl_logic/pa_temp [69]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b107|biu/cache_ctrl_logic/reg6_b68  (
    .a({_al_u2698_o,open_n81210}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [1]}),
    .c({\biu/paddress [107],\biu/paddress [68]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [41],_al_u2705_o}),
    .mi({\biu/paddress [107],\biu/paddress [68]}),
    .sr(rst_pad),
    .f({_al_u3080_o,haddr_pad[4]}),
    .q({\biu/cache_ctrl_logic/pa_temp [107],\biu/cache_ctrl_logic/pa_temp [68]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b108|biu/cache_ctrl_logic/reg6_b67  (
    .a({_al_u2698_o,open_n81228}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [0]}),
    .c({\biu/paddress [108],\biu/paddress [67]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [42],_al_u2705_o}),
    .mi({\biu/paddress [108],\biu/paddress [67]}),
    .sr(rst_pad),
    .f({_al_u3077_o,haddr_pad[3]}),
    .q({\biu/cache_ctrl_logic/pa_temp [108],\biu/cache_ctrl_logic/pa_temp [67]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b109|biu/cache_ctrl_logic/reg6_b127  (
    .a({_al_u2698_o,open_n81242}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [60]}),
    .c({\biu/paddress [109],\biu/paddress [127]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [43],_al_u2705_o}),
    .mi({\biu/paddress [109],\biu/paddress [127]}),
    .sr(rst_pad),
    .f({_al_u3074_o,haddr_pad[63]}),
    .q({\biu/cache_ctrl_logic/pa_temp [109],\biu/cache_ctrl_logic/pa_temp [127]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000101100000000),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b10|biu/bus_unit/mmu/reg1_b10  (
    .a({open_n81256,_al_u2914_o}),
    .b({\biu/paddress [10],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [10],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [10]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [10],\biu/paddress [10]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b110|biu/cache_ctrl_logic/reg6_b126  (
    .a({_al_u2698_o,open_n81275}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [59]}),
    .c({\biu/paddress [110],\biu/paddress [126]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [44],_al_u2705_o}),
    .mi({\biu/paddress [110],\biu/paddress [126]}),
    .sr(rst_pad),
    .f({_al_u3071_o,haddr_pad[62]}),
    .q({\biu/cache_ctrl_logic/pa_temp [110],\biu/cache_ctrl_logic/pa_temp [126]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b111|biu/cache_ctrl_logic/reg6_b125  (
    .a({_al_u2698_o,open_n81289}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [58]}),
    .c({\biu/paddress [111],\biu/paddress [125]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [45],_al_u2705_o}),
    .mi({\biu/paddress [111],\biu/paddress [125]}),
    .sr(rst_pad),
    .f({_al_u3068_o,haddr_pad[61]}),
    .q({\biu/cache_ctrl_logic/pa_temp [111],\biu/cache_ctrl_logic/pa_temp [125]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b112|biu/cache_ctrl_logic/reg6_b124  (
    .a({_al_u2698_o,open_n81307}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [57]}),
    .c({\biu/paddress [112],\biu/paddress [124]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [46],_al_u2705_o}),
    .mi({\biu/paddress [112],\biu/paddress [124]}),
    .sr(rst_pad),
    .f({_al_u3065_o,haddr_pad[60]}),
    .q({\biu/cache_ctrl_logic/pa_temp [112],\biu/cache_ctrl_logic/pa_temp [124]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b113|biu/cache_ctrl_logic/reg6_b123  (
    .a({_al_u2698_o,open_n81325}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [56]}),
    .c({\biu/paddress [113],\biu/paddress [123]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [47],_al_u2705_o}),
    .mi({\biu/paddress [113],\biu/paddress [123]}),
    .sr(rst_pad),
    .f({_al_u3062_o,haddr_pad[59]}),
    .q({\biu/cache_ctrl_logic/pa_temp [113],\biu/cache_ctrl_logic/pa_temp [123]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b114|biu/cache_ctrl_logic/reg6_b122  (
    .a({_al_u2698_o,open_n81339}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [55]}),
    .c({\biu/paddress [114],\biu/paddress [122]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [48],_al_u2705_o}),
    .mi({\biu/paddress [114],\biu/paddress [122]}),
    .sr(rst_pad),
    .f({_al_u3059_o,haddr_pad[58]}),
    .q({\biu/cache_ctrl_logic/pa_temp [114],\biu/cache_ctrl_logic/pa_temp [122]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b115|biu/cache_ctrl_logic/reg6_b121  (
    .a({_al_u2698_o,open_n81353}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [54]}),
    .c({\biu/paddress [115],\biu/paddress [121]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [49],_al_u2705_o}),
    .mi({\biu/paddress [115],\biu/paddress [121]}),
    .sr(rst_pad),
    .f({_al_u3056_o,haddr_pad[57]}),
    .q({\biu/cache_ctrl_logic/pa_temp [115],\biu/cache_ctrl_logic/pa_temp [121]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000101000101),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000101000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b116|biu/cache_ctrl_logic/reg6_b120  (
    .a({_al_u2698_o,open_n81371}),
    .b({\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ,\biu/bus_unit/n49 [53]}),
    .c({\biu/paddress [116],\biu/paddress [120]}),
    .ce(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .clk(clk_pad),
    .d({\biu/bus_unit/mmu_hwdata [50],_al_u2705_o}),
    .mi({\biu/paddress [116],\biu/paddress [120]}),
    .sr(rst_pad),
    .f({_al_u3053_o,haddr_pad[56]}),
    .q({\biu/cache_ctrl_logic/pa_temp [116],\biu/cache_ctrl_logic/pa_temp [120]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000101100000000),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b11|biu/bus_unit/mmu/reg1_b11  (
    .a({open_n81389,_al_u2914_o}),
    .b({\biu/paddress [11],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [11],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [11]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [11],\biu/paddress [11]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000101100000000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1000101100000000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b1|biu/bus_unit/mmu/reg1_b1  (
    .a({open_n81408,_al_u2914_o}),
    .b({\biu/paddress [1],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [1],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [1]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [1],\biu/paddress [1]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000101100000000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1000101100000000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b2|biu/bus_unit/mmu/reg1_b2  (
    .a({open_n81431,_al_u2914_o}),
    .b({\biu/paddress [2],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [2],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [2]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [2],\biu/paddress [2]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b30|biu/cache_ctrl_logic/reg6_b60  (
    .b({\biu/paddress [30],\biu/paddress [60]}),
    .c({\biu/cache_ctrl_logic/pa_temp [30],\biu/cache_ctrl_logic/pa_temp [60]}),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o }),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [30],\biu/cache_ctrl_logic/pa_temp [60]}));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000101100000000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1000101100000000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b3|biu/bus_unit/mmu/reg1_b3  (
    .a({open_n81478,_al_u2914_o}),
    .b({\biu/paddress [3],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [3],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [3]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [3],\biu/paddress [3]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000101100000000),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b4|biu/bus_unit/mmu/reg1_b4  (
    .a({open_n81501,_al_u2914_o}),
    .b({\biu/paddress [4],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [4],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [4]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [4],\biu/paddress [4]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000101100000000),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b5|biu/bus_unit/mmu/reg1_b5  (
    .a({open_n81520,_al_u2914_o}),
    .b({\biu/paddress [5],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [5],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [5]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [5],\biu/paddress [5]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000101100000000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1000101100000000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b6|biu/bus_unit/mmu/reg1_b6  (
    .a({open_n81539,_al_u2914_o}),
    .b({\biu/paddress [6],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [6],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [6]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [6],\biu/paddress [6]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000101100000000),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b1000101100000000),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b7|biu/bus_unit/mmu/reg1_b7  (
    .a({open_n81562,_al_u2914_o}),
    .b({\biu/paddress [7],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [7],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [7]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [7],\biu/paddress [7]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000101100000000),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b8|biu/bus_unit/mmu/reg1_b8  (
    .a({open_n81585,_al_u2914_o}),
    .b({\biu/paddress [8],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [8],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [8]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [8],\biu/paddress [8]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  EG_PHY_MSLICE #(
    //.LUT0("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000101100000000),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg6_b9|biu/bus_unit/mmu/reg1_b9  (
    .a({open_n81604,_al_u2914_o}),
    .b({\biu/paddress [9],_al_u2698_o}),
    .c({\biu/cache_ctrl_logic/pa_temp [9],\biu/bus_unit/mmu/mux24_b0_sel_is_1_o }),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ,\biu/paddress [9]}),
    .sr(rst_pad),
    .q({\biu/cache_ctrl_logic/pa_temp [9],\biu/paddress [9]}));  // ../../RTL/CPU/BIU/mmu.v(183)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(~A*~(~C*~B)))"),
    //.LUTF1("~(C*~(B*~D))"),
    //.LUTG0("~(D*~(~A*~(~C*~B)))"),
    //.LUTG1("~(C*~(B*~D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010011111111),
    .INIT_LUTF1(16'b0000111111001111),
    .INIT_LUTG0(16'b0101010011111111),
    .INIT_LUTG1(16'b0000111111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \biu/cache_ctrl_logic/reg8_b1|biu/cache_ctrl_logic/reg8_b0  (
    .a({open_n81623,_al_u9676_o}),
    .b({_al_u9713_o,_al_u9692_o}),
    .c({_al_u9693_o,_al_u9285_o}),
    .clk(clk_pad),
    .d({_al_u9676_o,_al_u9693_o}),
    .sr(rst_pad),
    .q(\biu/cache_ctrl_logic/statu [1:0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("DISABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u0|cu_ru/add0_2/ucin  (
    .a({\cu_ru/tvec [4],1'b0}),
    .b({\cu_ru/trap_cause [0],open_n81693}),
    .f({\cu_ru/n43 [0],open_n81713}),
    .fco(\cu_ru/add0_2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u10|cu_ru/add0_2/u9  (
    .a(\cu_ru/tvec [14:13]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c9 ),
    .f(\cu_ru/n43 [10:9]),
    .fco(\cu_ru/add0_2/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u12|cu_ru/add0_2/u11  (
    .a(\cu_ru/tvec [16:15]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c11 ),
    .f(\cu_ru/n43 [12:11]),
    .fco(\cu_ru/add0_2/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u14|cu_ru/add0_2/u13  (
    .a(\cu_ru/tvec [18:17]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c13 ),
    .f(\cu_ru/n43 [14:13]),
    .fco(\cu_ru/add0_2/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u16|cu_ru/add0_2/u15  (
    .a(\cu_ru/tvec [20:19]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c15 ),
    .f(\cu_ru/n43 [16:15]),
    .fco(\cu_ru/add0_2/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u18|cu_ru/add0_2/u17  (
    .a(\cu_ru/tvec [22:21]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c17 ),
    .f(\cu_ru/n43 [18:17]),
    .fco(\cu_ru/add0_2/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u20|cu_ru/add0_2/u19  (
    .a(\cu_ru/tvec [24:23]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c19 ),
    .f(\cu_ru/n43 [20:19]),
    .fco(\cu_ru/add0_2/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u22|cu_ru/add0_2/u21  (
    .a(\cu_ru/tvec [26:25]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c21 ),
    .f(\cu_ru/n43 [22:21]),
    .fco(\cu_ru/add0_2/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u24|cu_ru/add0_2/u23  (
    .a(\cu_ru/tvec [28:27]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c23 ),
    .f(\cu_ru/n43 [24:23]),
    .fco(\cu_ru/add0_2/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u26|cu_ru/add0_2/u25  (
    .a(\cu_ru/tvec [30:29]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c25 ),
    .f(\cu_ru/n43 [26:25]),
    .fco(\cu_ru/add0_2/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u28|cu_ru/add0_2/u27  (
    .a(\cu_ru/tvec [32:31]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c27 ),
    .f(\cu_ru/n43 [28:27]),
    .fco(\cu_ru/add0_2/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u2|cu_ru/add0_2/u1  (
    .a(\cu_ru/tvec [6:5]),
    .b(\cu_ru/trap_cause [2:1]),
    .fci(\cu_ru/add0_2/c1 ),
    .f(\cu_ru/n43 [2:1]),
    .fco(\cu_ru/add0_2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u30|cu_ru/add0_2/u29  (
    .a(\cu_ru/tvec [34:33]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c29 ),
    .f(\cu_ru/n43 [30:29]),
    .fco(\cu_ru/add0_2/c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u32|cu_ru/add0_2/u31  (
    .a(\cu_ru/tvec [36:35]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c31 ),
    .f(\cu_ru/n43 [32:31]),
    .fco(\cu_ru/add0_2/c33 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y8Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u34|cu_ru/add0_2/u33  (
    .a(\cu_ru/tvec [38:37]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c33 ),
    .f(\cu_ru/n43 [34:33]),
    .fco(\cu_ru/add0_2/c35 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y9Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u36|cu_ru/add0_2/u35  (
    .a(\cu_ru/tvec [40:39]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c35 ),
    .f(\cu_ru/n43 [36:35]),
    .fco(\cu_ru/add0_2/c37 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y9Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u38|cu_ru/add0_2/u37  (
    .a(\cu_ru/tvec [42:41]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c37 ),
    .f(\cu_ru/n43 [38:37]),
    .fco(\cu_ru/add0_2/c39 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y10Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u40|cu_ru/add0_2/u39  (
    .a(\cu_ru/tvec [44:43]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c39 ),
    .f(\cu_ru/n43 [40:39]),
    .fco(\cu_ru/add0_2/c41 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y10Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u42|cu_ru/add0_2/u41  (
    .a(\cu_ru/tvec [46:45]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c41 ),
    .f(\cu_ru/n43 [42:41]),
    .fco(\cu_ru/add0_2/c43 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y11Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u44|cu_ru/add0_2/u43  (
    .a(\cu_ru/tvec [48:47]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c43 ),
    .f(\cu_ru/n43 [44:43]),
    .fco(\cu_ru/add0_2/c45 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y11Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u46|cu_ru/add0_2/u45  (
    .a(\cu_ru/tvec [50:49]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c45 ),
    .f(\cu_ru/n43 [46:45]),
    .fco(\cu_ru/add0_2/c47 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y12Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u48|cu_ru/add0_2/u47  (
    .a(\cu_ru/tvec [52:51]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c47 ),
    .f(\cu_ru/n43 [48:47]),
    .fco(\cu_ru/add0_2/c49 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u4|cu_ru/add0_2/u3  (
    .a(\cu_ru/tvec [8:7]),
    .b({1'b0,\cu_ru/trap_cause [3]}),
    .fci(\cu_ru/add0_2/c3 ),
    .f(\cu_ru/n43 [4:3]),
    .fco(\cu_ru/add0_2/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y12Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u50|cu_ru/add0_2/u49  (
    .a(\cu_ru/tvec [54:53]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c49 ),
    .f(\cu_ru/n43 [50:49]),
    .fco(\cu_ru/add0_2/c51 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y13Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u52|cu_ru/add0_2/u51  (
    .a(\cu_ru/tvec [56:55]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c51 ),
    .f(\cu_ru/n43 [52:51]),
    .fco(\cu_ru/add0_2/c53 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y13Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u54|cu_ru/add0_2/u53  (
    .a(\cu_ru/tvec [58:57]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c53 ),
    .f(\cu_ru/n43 [54:53]),
    .fco(\cu_ru/add0_2/c55 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y14Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u56|cu_ru/add0_2/u55  (
    .a(\cu_ru/tvec [60:59]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c55 ),
    .f(\cu_ru/n43 [56:55]),
    .fco(\cu_ru/add0_2/c57 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y14Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u58|cu_ru/add0_2/u57  (
    .a(\cu_ru/tvec [62:61]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c57 ),
    .f(\cu_ru/n43 [58:57]),
    .fco(\cu_ru/add0_2/c59 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u6|cu_ru/add0_2/u5  (
    .a(\cu_ru/tvec [10:9]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c5 ),
    .f(\cu_ru/n43 [6:5]),
    .fco(\cu_ru/add0_2/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/u8|cu_ru/add0_2/u7  (
    .a(\cu_ru/tvec [12:11]),
    .b(2'b00),
    .fci(\cu_ru/add0_2/c7 ),
    .f(\cu_ru/n43 [8:7]),
    .fco(\cu_ru/add0_2/c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/add0_2/u0|cu_ru/add0_2/ucin"),
    //.R_POSITION("X0Y15Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \cu_ru/add0_2/ucout|cu_ru/add0_2/u59  (
    .a({open_n82356,\cu_ru/tvec [63]}),
    .b({open_n82357,1'b0}),
    .fci(\cu_ru/add0_2/c59 ),
    .f({\cu_ru/add0_2_co ,\cu_ru/n43 [59]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c0_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c0_l  (
    .a({data_rd[0],\cu_ru/n52 [0]}),
    .b({data_rd[1],\cu_ru/n52 [1]}),
    .c({data_rd[2],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[3],\cu_ru/n52 [3]}),
    .e({open_n82382,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c0_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c0_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c0_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c0_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c0_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_001 ,\cu_ru/al_ram_gpr_al_u0_do_i0_000 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c0_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c0_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c0_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c0_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_003 ,\cu_ru/al_ram_gpr_al_u0_do_i0_002 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c10_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c10_l  (
    .a({data_rd[40],\cu_ru/n52 [0]}),
    .b({data_rd[41],\cu_ru/n52 [1]}),
    .c({data_rd[42],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[43],\cu_ru/n52 [3]}),
    .e({open_n82417,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c10_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c10_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c10_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c10_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c10_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c10_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_041 ,\cu_ru/al_ram_gpr_al_u0_do_i0_040 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c10_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c10_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c10_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c10_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_043 ,\cu_ru/al_ram_gpr_al_u0_do_i0_042 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c11_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c11_l  (
    .a({data_rd[44],\cu_ru/n52 [0]}),
    .b({data_rd[45],\cu_ru/n52 [1]}),
    .c({data_rd[46],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[47],\cu_ru/n52 [3]}),
    .e({open_n82452,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c11_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c11_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c11_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c11_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c11_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c11_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_045 ,\cu_ru/al_ram_gpr_al_u0_do_i0_044 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c11_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c11_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c11_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c11_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_047 ,\cu_ru/al_ram_gpr_al_u0_do_i0_046 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c12_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c12_l  (
    .a({data_rd[48],\cu_ru/n52 [0]}),
    .b({data_rd[49],\cu_ru/n52 [1]}),
    .c({data_rd[50],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[51],\cu_ru/n52 [3]}),
    .e({open_n82487,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c12_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c12_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c12_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c12_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c12_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c12_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_049 ,\cu_ru/al_ram_gpr_al_u0_do_i0_048 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c12_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c12_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c12_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c12_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_051 ,\cu_ru/al_ram_gpr_al_u0_do_i0_050 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c13_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c13_l  (
    .a({data_rd[52],\cu_ru/n52 [0]}),
    .b({data_rd[53],\cu_ru/n52 [1]}),
    .c({data_rd[54],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[55],\cu_ru/n52 [3]}),
    .e({open_n82522,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c13_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c13_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c13_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c13_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c13_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c13_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_053 ,\cu_ru/al_ram_gpr_al_u0_do_i0_052 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c13_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c13_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c13_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c13_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_055 ,\cu_ru/al_ram_gpr_al_u0_do_i0_054 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c14_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c14_l  (
    .a({data_rd[56],\cu_ru/n52 [0]}),
    .b({data_rd[57],\cu_ru/n52 [1]}),
    .c({data_rd[58],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[59],\cu_ru/n52 [3]}),
    .e({open_n82557,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c14_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c14_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c14_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c14_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c14_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c14_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_057 ,\cu_ru/al_ram_gpr_al_u0_do_i0_056 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c14_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c14_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c14_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c14_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_059 ,\cu_ru/al_ram_gpr_al_u0_do_i0_058 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c15_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c15_l  (
    .a({data_rd[60],\cu_ru/n52 [0]}),
    .b({data_rd[61],\cu_ru/n52 [1]}),
    .c({data_rd[62],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[63],\cu_ru/n52 [3]}),
    .e({open_n82592,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c15_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c15_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c15_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c15_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c15_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c15_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_061 ,\cu_ru/al_ram_gpr_al_u0_do_i0_060 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c15_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c15_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c15_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c15_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_063 ,\cu_ru/al_ram_gpr_al_u0_do_i0_062 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c1_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c1_l  (
    .a({data_rd[4],\cu_ru/n52 [0]}),
    .b({data_rd[5],\cu_ru/n52 [1]}),
    .c({data_rd[6],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[7],\cu_ru/n52 [3]}),
    .e({open_n82627,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c1_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c1_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c1_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c1_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c1_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_005 ,\cu_ru/al_ram_gpr_al_u0_do_i0_004 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c1_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c1_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c1_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c1_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_007 ,\cu_ru/al_ram_gpr_al_u0_do_i0_006 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c2_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c2_l  (
    .a({data_rd[8],\cu_ru/n52 [0]}),
    .b({data_rd[9],\cu_ru/n52 [1]}),
    .c({data_rd[10],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[11],\cu_ru/n52 [3]}),
    .e({open_n82662,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c2_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c2_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c2_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c2_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c2_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_009 ,\cu_ru/al_ram_gpr_al_u0_do_i0_008 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c2_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c2_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c2_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c2_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_011 ,\cu_ru/al_ram_gpr_al_u0_do_i0_010 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c3_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c3_l  (
    .a({data_rd[12],\cu_ru/n52 [0]}),
    .b({data_rd[13],\cu_ru/n52 [1]}),
    .c({data_rd[14],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[15],\cu_ru/n52 [3]}),
    .e({open_n82697,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c3_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c3_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c3_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c3_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c3_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_013 ,\cu_ru/al_ram_gpr_al_u0_do_i0_012 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c3_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c3_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c3_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c3_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_015 ,\cu_ru/al_ram_gpr_al_u0_do_i0_014 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c4_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c4_l  (
    .a({data_rd[16],\cu_ru/n52 [0]}),
    .b({data_rd[17],\cu_ru/n52 [1]}),
    .c({data_rd[18],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[19],\cu_ru/n52 [3]}),
    .e({open_n82732,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c4_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c4_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c4_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c4_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c4_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_017 ,\cu_ru/al_ram_gpr_al_u0_do_i0_016 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c4_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c4_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c4_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c4_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_019 ,\cu_ru/al_ram_gpr_al_u0_do_i0_018 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c5_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c5_l  (
    .a({data_rd[20],\cu_ru/n52 [0]}),
    .b({data_rd[21],\cu_ru/n52 [1]}),
    .c({data_rd[22],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[23],\cu_ru/n52 [3]}),
    .e({open_n82767,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c5_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c5_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c5_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c5_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c5_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_021 ,\cu_ru/al_ram_gpr_al_u0_do_i0_020 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c5_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c5_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c5_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c5_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_023 ,\cu_ru/al_ram_gpr_al_u0_do_i0_022 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c6_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c6_l  (
    .a({data_rd[24],\cu_ru/n52 [0]}),
    .b({data_rd[25],\cu_ru/n52 [1]}),
    .c({data_rd[26],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[27],\cu_ru/n52 [3]}),
    .e({open_n82802,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c6_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c6_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c6_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c6_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c6_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_025 ,\cu_ru/al_ram_gpr_al_u0_do_i0_024 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c6_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c6_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c6_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c6_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_027 ,\cu_ru/al_ram_gpr_al_u0_do_i0_026 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c7_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c7_l  (
    .a({data_rd[28],\cu_ru/n52 [0]}),
    .b({data_rd[29],\cu_ru/n52 [1]}),
    .c({data_rd[30],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[31],\cu_ru/n52 [3]}),
    .e({open_n82837,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c7_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c7_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c7_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c7_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c7_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_029 ,\cu_ru/al_ram_gpr_al_u0_do_i0_028 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c7_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c7_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c7_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c7_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_031 ,\cu_ru/al_ram_gpr_al_u0_do_i0_030 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c8_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c8_l  (
    .a({data_rd[32],\cu_ru/n52 [0]}),
    .b({data_rd[33],\cu_ru/n52 [1]}),
    .c({data_rd[34],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[35],\cu_ru/n52 [3]}),
    .e({open_n82872,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c8_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c8_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c8_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c8_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c8_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c8_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_033 ,\cu_ru/al_ram_gpr_al_u0_do_i0_032 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c8_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c8_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c8_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c8_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_035 ,\cu_ru/al_ram_gpr_al_u0_do_i0_034 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c9_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r0_c9_l  (
    .a({data_rd[36],\cu_ru/n52 [0]}),
    .b({data_rd[37],\cu_ru/n52 [1]}),
    .c({data_rd[38],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[39],\cu_ru/n52 [3]}),
    .e({open_n82907,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c9_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c9_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c9_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c9_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c9_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c9_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_037 ,\cu_ru/al_ram_gpr_al_u0_do_i0_036 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r0_c9_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r0_c9_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r0_c9_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r0_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r0_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r0_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r0_c9_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i0_039 ,\cu_ru/al_ram_gpr_al_u0_do_i0_038 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c0_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c0_l  (
    .a({data_rd[0],\cu_ru/n52 [0]}),
    .b({data_rd[1],\cu_ru/n52 [1]}),
    .c({data_rd[2],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[3],\cu_ru/n52 [3]}),
    .e({open_n82942,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c0_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c0_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c0_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c0_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c0_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_001 ,\cu_ru/al_ram_gpr_al_u0_do_i1_000 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c0_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c0_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c0_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c0_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_003 ,\cu_ru/al_ram_gpr_al_u0_do_i1_002 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c10_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c10_l  (
    .a({data_rd[40],\cu_ru/n52 [0]}),
    .b({data_rd[41],\cu_ru/n52 [1]}),
    .c({data_rd[42],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[43],\cu_ru/n52 [3]}),
    .e({open_n82977,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c10_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c10_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c10_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c10_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c10_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c10_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_041 ,\cu_ru/al_ram_gpr_al_u0_do_i1_040 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c10_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c10_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c10_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c10_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_043 ,\cu_ru/al_ram_gpr_al_u0_do_i1_042 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c11_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c11_l  (
    .a({data_rd[44],\cu_ru/n52 [0]}),
    .b({data_rd[45],\cu_ru/n52 [1]}),
    .c({data_rd[46],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[47],\cu_ru/n52 [3]}),
    .e({open_n83012,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c11_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c11_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c11_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c11_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c11_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c11_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_045 ,\cu_ru/al_ram_gpr_al_u0_do_i1_044 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c11_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c11_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c11_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c11_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_047 ,\cu_ru/al_ram_gpr_al_u0_do_i1_046 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c12_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c12_l  (
    .a({data_rd[48],\cu_ru/n52 [0]}),
    .b({data_rd[49],\cu_ru/n52 [1]}),
    .c({data_rd[50],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[51],\cu_ru/n52 [3]}),
    .e({open_n83047,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c12_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c12_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c12_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c12_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c12_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c12_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_049 ,\cu_ru/al_ram_gpr_al_u0_do_i1_048 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c12_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c12_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c12_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c12_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_051 ,\cu_ru/al_ram_gpr_al_u0_do_i1_050 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c13_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c13_l  (
    .a({data_rd[52],\cu_ru/n52 [0]}),
    .b({data_rd[53],\cu_ru/n52 [1]}),
    .c({data_rd[54],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[55],\cu_ru/n52 [3]}),
    .e({open_n83082,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c13_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c13_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c13_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c13_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c13_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c13_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_053 ,\cu_ru/al_ram_gpr_al_u0_do_i1_052 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c13_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c13_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c13_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c13_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_055 ,\cu_ru/al_ram_gpr_al_u0_do_i1_054 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c14_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c14_l  (
    .a({data_rd[56],\cu_ru/n52 [0]}),
    .b({data_rd[57],\cu_ru/n52 [1]}),
    .c({data_rd[58],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[59],\cu_ru/n52 [3]}),
    .e({open_n83117,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c14_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c14_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c14_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c14_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c14_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c14_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_057 ,\cu_ru/al_ram_gpr_al_u0_do_i1_056 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c14_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c14_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c14_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c14_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_059 ,\cu_ru/al_ram_gpr_al_u0_do_i1_058 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c15_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c15_l  (
    .a({data_rd[60],\cu_ru/n52 [0]}),
    .b({data_rd[61],\cu_ru/n52 [1]}),
    .c({data_rd[62],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[63],\cu_ru/n52 [3]}),
    .e({open_n83152,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c15_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c15_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c15_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c15_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c15_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c15_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_061 ,\cu_ru/al_ram_gpr_al_u0_do_i1_060 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c15_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c15_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c15_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c15_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_063 ,\cu_ru/al_ram_gpr_al_u0_do_i1_062 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c1_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c1_l  (
    .a({data_rd[4],\cu_ru/n52 [0]}),
    .b({data_rd[5],\cu_ru/n52 [1]}),
    .c({data_rd[6],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[7],\cu_ru/n52 [3]}),
    .e({open_n83187,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c1_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c1_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c1_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c1_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c1_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_005 ,\cu_ru/al_ram_gpr_al_u0_do_i1_004 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c1_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c1_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c1_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c1_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_007 ,\cu_ru/al_ram_gpr_al_u0_do_i1_006 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c2_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c2_l  (
    .a({data_rd[8],\cu_ru/n52 [0]}),
    .b({data_rd[9],\cu_ru/n52 [1]}),
    .c({data_rd[10],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[11],\cu_ru/n52 [3]}),
    .e({open_n83222,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c2_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c2_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c2_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c2_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c2_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_009 ,\cu_ru/al_ram_gpr_al_u0_do_i1_008 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c2_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c2_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c2_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c2_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_011 ,\cu_ru/al_ram_gpr_al_u0_do_i1_010 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c3_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c3_l  (
    .a({data_rd[12],\cu_ru/n52 [0]}),
    .b({data_rd[13],\cu_ru/n52 [1]}),
    .c({data_rd[14],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[15],\cu_ru/n52 [3]}),
    .e({open_n83257,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c3_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c3_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c3_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c3_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c3_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_013 ,\cu_ru/al_ram_gpr_al_u0_do_i1_012 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c3_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c3_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c3_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c3_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_015 ,\cu_ru/al_ram_gpr_al_u0_do_i1_014 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c4_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c4_l  (
    .a({data_rd[16],\cu_ru/n52 [0]}),
    .b({data_rd[17],\cu_ru/n52 [1]}),
    .c({data_rd[18],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[19],\cu_ru/n52 [3]}),
    .e({open_n83292,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c4_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c4_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c4_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c4_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c4_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_017 ,\cu_ru/al_ram_gpr_al_u0_do_i1_016 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c4_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c4_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c4_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c4_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_019 ,\cu_ru/al_ram_gpr_al_u0_do_i1_018 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c5_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c5_l  (
    .a({data_rd[20],\cu_ru/n52 [0]}),
    .b({data_rd[21],\cu_ru/n52 [1]}),
    .c({data_rd[22],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[23],\cu_ru/n52 [3]}),
    .e({open_n83327,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c5_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c5_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c5_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c5_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c5_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_021 ,\cu_ru/al_ram_gpr_al_u0_do_i1_020 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c5_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c5_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c5_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c5_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_023 ,\cu_ru/al_ram_gpr_al_u0_do_i1_022 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c6_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c6_l  (
    .a({data_rd[24],\cu_ru/n52 [0]}),
    .b({data_rd[25],\cu_ru/n52 [1]}),
    .c({data_rd[26],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[27],\cu_ru/n52 [3]}),
    .e({open_n83362,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c6_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c6_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c6_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c6_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c6_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_025 ,\cu_ru/al_ram_gpr_al_u0_do_i1_024 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c6_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c6_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c6_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c6_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_027 ,\cu_ru/al_ram_gpr_al_u0_do_i1_026 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c7_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c7_l  (
    .a({data_rd[28],\cu_ru/n52 [0]}),
    .b({data_rd[29],\cu_ru/n52 [1]}),
    .c({data_rd[30],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[31],\cu_ru/n52 [3]}),
    .e({open_n83397,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c7_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c7_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c7_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c7_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c7_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_029 ,\cu_ru/al_ram_gpr_al_u0_do_i1_028 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c7_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c7_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c7_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c7_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_031 ,\cu_ru/al_ram_gpr_al_u0_do_i1_030 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c8_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c8_l  (
    .a({data_rd[32],\cu_ru/n52 [0]}),
    .b({data_rd[33],\cu_ru/n52 [1]}),
    .c({data_rd[34],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[35],\cu_ru/n52 [3]}),
    .e({open_n83432,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c8_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c8_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c8_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c8_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c8_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c8_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_033 ,\cu_ru/al_ram_gpr_al_u0_do_i1_032 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c8_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c8_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c8_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c8_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_035 ,\cu_ru/al_ram_gpr_al_u0_do_i1_034 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c9_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_al_u0_r1_c9_l  (
    .a({data_rd[36],\cu_ru/n52 [0]}),
    .b({data_rd[37],\cu_ru/n52 [1]}),
    .c({data_rd[38],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[39],\cu_ru/n52 [3]}),
    .e({open_n83467,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c9_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c9_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c9_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c9_m0  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c9_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c9_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_037 ,\cu_ru/al_ram_gpr_al_u0_do_i1_036 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_al_u0_r1_c9_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_al_u0_r1_c9_m1  (
    .a({\cu_ru/n49 [0],\cu_ru/n49 [0]}),
    .b({\cu_ru/n49 [1],\cu_ru/n49 [1]}),
    .c({\cu_ru/n49 [2],\cu_ru/n49 [2]}),
    .d({\cu_ru/n49 [3],\cu_ru/n49 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_al_u0_r1_c9_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_al_u0_r1_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_al_u0_r1_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_al_u0_r1_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_al_u0_r1_c9_we ),
    .f({\cu_ru/al_ram_gpr_al_u0_do_i1_039 ,\cu_ru/al_ram_gpr_al_u0_do_i1_038 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c0_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c0_l  (
    .a({data_rd[0],\cu_ru/n52 [0]}),
    .b({data_rd[1],\cu_ru/n52 [1]}),
    .c({data_rd[2],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[3],\cu_ru/n52 [3]}),
    .e({open_n83502,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c0_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c0_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c0_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c0_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c0_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_001 ,\cu_ru/al_ram_gpr_do_i0_000 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c0_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c0_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c0_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c0_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_003 ,\cu_ru/al_ram_gpr_do_i0_002 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c10_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c10_l  (
    .a({data_rd[40],\cu_ru/n52 [0]}),
    .b({data_rd[41],\cu_ru/n52 [1]}),
    .c({data_rd[42],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[43],\cu_ru/n52 [3]}),
    .e({open_n83537,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c10_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c10_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c10_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c10_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c10_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c10_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_041 ,\cu_ru/al_ram_gpr_do_i0_040 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c10_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c10_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c10_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c10_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_043 ,\cu_ru/al_ram_gpr_do_i0_042 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c11_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c11_l  (
    .a({data_rd[44],\cu_ru/n52 [0]}),
    .b({data_rd[45],\cu_ru/n52 [1]}),
    .c({data_rd[46],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[47],\cu_ru/n52 [3]}),
    .e({open_n83572,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c11_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c11_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c11_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c11_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c11_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c11_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_045 ,\cu_ru/al_ram_gpr_do_i0_044 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c11_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c11_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c11_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c11_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_047 ,\cu_ru/al_ram_gpr_do_i0_046 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c12_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c12_l  (
    .a({data_rd[48],\cu_ru/n52 [0]}),
    .b({data_rd[49],\cu_ru/n52 [1]}),
    .c({data_rd[50],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[51],\cu_ru/n52 [3]}),
    .e({open_n83607,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c12_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c12_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c12_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c12_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c12_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c12_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_049 ,\cu_ru/al_ram_gpr_do_i0_048 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c12_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c12_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c12_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c12_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_051 ,\cu_ru/al_ram_gpr_do_i0_050 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c13_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c13_l  (
    .a({data_rd[52],\cu_ru/n52 [0]}),
    .b({data_rd[53],\cu_ru/n52 [1]}),
    .c({data_rd[54],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[55],\cu_ru/n52 [3]}),
    .e({open_n83642,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c13_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c13_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c13_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c13_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c13_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c13_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_053 ,\cu_ru/al_ram_gpr_do_i0_052 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c13_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c13_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c13_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c13_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_055 ,\cu_ru/al_ram_gpr_do_i0_054 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c14_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c14_l  (
    .a({data_rd[56],\cu_ru/n52 [0]}),
    .b({data_rd[57],\cu_ru/n52 [1]}),
    .c({data_rd[58],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[59],\cu_ru/n52 [3]}),
    .e({open_n83677,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c14_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c14_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c14_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c14_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c14_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c14_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_057 ,\cu_ru/al_ram_gpr_do_i0_056 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c14_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c14_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c14_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c14_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_059 ,\cu_ru/al_ram_gpr_do_i0_058 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c15_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c15_l  (
    .a({data_rd[60],\cu_ru/n52 [0]}),
    .b({data_rd[61],\cu_ru/n52 [1]}),
    .c({data_rd[62],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[63],\cu_ru/n52 [3]}),
    .e({open_n83712,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c15_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c15_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c15_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c15_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c15_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c15_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_061 ,\cu_ru/al_ram_gpr_do_i0_060 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c15_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c15_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c15_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c15_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_063 ,\cu_ru/al_ram_gpr_do_i0_062 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c1_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c1_l  (
    .a({data_rd[4],\cu_ru/n52 [0]}),
    .b({data_rd[5],\cu_ru/n52 [1]}),
    .c({data_rd[6],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[7],\cu_ru/n52 [3]}),
    .e({open_n83747,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c1_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c1_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c1_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c1_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c1_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_005 ,\cu_ru/al_ram_gpr_do_i0_004 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c1_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c1_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c1_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c1_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_007 ,\cu_ru/al_ram_gpr_do_i0_006 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c2_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c2_l  (
    .a({data_rd[8],\cu_ru/n52 [0]}),
    .b({data_rd[9],\cu_ru/n52 [1]}),
    .c({data_rd[10],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[11],\cu_ru/n52 [3]}),
    .e({open_n83782,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c2_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c2_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c2_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c2_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c2_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_009 ,\cu_ru/al_ram_gpr_do_i0_008 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c2_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c2_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c2_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c2_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_011 ,\cu_ru/al_ram_gpr_do_i0_010 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c3_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c3_l  (
    .a({data_rd[12],\cu_ru/n52 [0]}),
    .b({data_rd[13],\cu_ru/n52 [1]}),
    .c({data_rd[14],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[15],\cu_ru/n52 [3]}),
    .e({open_n83817,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c3_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c3_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c3_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c3_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c3_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_013 ,\cu_ru/al_ram_gpr_do_i0_012 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c3_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c3_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c3_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c3_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_015 ,\cu_ru/al_ram_gpr_do_i0_014 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c4_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c4_l  (
    .a({data_rd[16],\cu_ru/n52 [0]}),
    .b({data_rd[17],\cu_ru/n52 [1]}),
    .c({data_rd[18],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[19],\cu_ru/n52 [3]}),
    .e({open_n83852,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c4_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c4_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c4_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c4_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c4_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_017 ,\cu_ru/al_ram_gpr_do_i0_016 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c4_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c4_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c4_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c4_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_019 ,\cu_ru/al_ram_gpr_do_i0_018 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c5_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c5_l  (
    .a({data_rd[20],\cu_ru/n52 [0]}),
    .b({data_rd[21],\cu_ru/n52 [1]}),
    .c({data_rd[22],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[23],\cu_ru/n52 [3]}),
    .e({open_n83887,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c5_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c5_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c5_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c5_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c5_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_021 ,\cu_ru/al_ram_gpr_do_i0_020 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c5_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c5_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c5_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c5_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_023 ,\cu_ru/al_ram_gpr_do_i0_022 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c6_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c6_l  (
    .a({data_rd[24],\cu_ru/n52 [0]}),
    .b({data_rd[25],\cu_ru/n52 [1]}),
    .c({data_rd[26],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[27],\cu_ru/n52 [3]}),
    .e({open_n83922,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c6_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c6_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c6_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c6_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c6_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_025 ,\cu_ru/al_ram_gpr_do_i0_024 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c6_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c6_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c6_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c6_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_027 ,\cu_ru/al_ram_gpr_do_i0_026 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c7_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c7_l  (
    .a({data_rd[28],\cu_ru/n52 [0]}),
    .b({data_rd[29],\cu_ru/n52 [1]}),
    .c({data_rd[30],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[31],\cu_ru/n52 [3]}),
    .e({open_n83957,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c7_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c7_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c7_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c7_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c7_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_029 ,\cu_ru/al_ram_gpr_do_i0_028 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c7_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c7_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c7_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c7_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_031 ,\cu_ru/al_ram_gpr_do_i0_030 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c8_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c8_l  (
    .a({data_rd[32],\cu_ru/n52 [0]}),
    .b({data_rd[33],\cu_ru/n52 [1]}),
    .c({data_rd[34],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[35],\cu_ru/n52 [3]}),
    .e({open_n83992,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c8_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c8_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c8_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c8_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c8_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c8_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_033 ,\cu_ru/al_ram_gpr_do_i0_032 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c8_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c8_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c8_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c8_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_035 ,\cu_ru/al_ram_gpr_do_i0_034 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c9_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r0_c9_l  (
    .a({data_rd[36],\cu_ru/n52 [0]}),
    .b({data_rd[37],\cu_ru/n52 [1]}),
    .c({data_rd[38],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[39],\cu_ru/n52 [3]}),
    .e({open_n84027,\cu_ru/n53_0_al_n1985 }),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c9_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c9_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c9_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c9_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c9_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c9_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_037 ,\cu_ru/al_ram_gpr_do_i0_036 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r0_c9_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r0_c9_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r0_c9_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r0_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r0_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r0_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r0_c9_we ),
    .f({\cu_ru/al_ram_gpr_do_i0_039 ,\cu_ru/al_ram_gpr_do_i0_038 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c0_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c0_l  (
    .a({data_rd[0],\cu_ru/n52 [0]}),
    .b({data_rd[1],\cu_ru/n52 [1]}),
    .c({data_rd[2],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[3],\cu_ru/n52 [3]}),
    .e({open_n84062,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c0_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c0_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c0_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c0_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c0_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_001 ,\cu_ru/al_ram_gpr_do_i1_000 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c0_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c0_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c0_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c0_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c0_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c0_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c0_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_003 ,\cu_ru/al_ram_gpr_do_i1_002 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c10_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c10_l  (
    .a({data_rd[40],\cu_ru/n52 [0]}),
    .b({data_rd[41],\cu_ru/n52 [1]}),
    .c({data_rd[42],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[43],\cu_ru/n52 [3]}),
    .e({open_n84097,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c10_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c10_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c10_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c10_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c10_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c10_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_041 ,\cu_ru/al_ram_gpr_do_i1_040 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c10_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c10_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c10_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c10_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c10_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c10_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c10_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_043 ,\cu_ru/al_ram_gpr_do_i1_042 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c11_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c11_l  (
    .a({data_rd[44],\cu_ru/n52 [0]}),
    .b({data_rd[45],\cu_ru/n52 [1]}),
    .c({data_rd[46],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[47],\cu_ru/n52 [3]}),
    .e({open_n84132,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c11_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c11_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c11_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c11_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c11_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c11_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_045 ,\cu_ru/al_ram_gpr_do_i1_044 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c11_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c11_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c11_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c11_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c11_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c11_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c11_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_047 ,\cu_ru/al_ram_gpr_do_i1_046 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c12_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c12_l  (
    .a({data_rd[48],\cu_ru/n52 [0]}),
    .b({data_rd[49],\cu_ru/n52 [1]}),
    .c({data_rd[50],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[51],\cu_ru/n52 [3]}),
    .e({open_n84167,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c12_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c12_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c12_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c12_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c12_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c12_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_049 ,\cu_ru/al_ram_gpr_do_i1_048 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c12_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c12_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c12_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c12_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c12_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c12_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c12_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_051 ,\cu_ru/al_ram_gpr_do_i1_050 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c13_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c13_l  (
    .a({data_rd[52],\cu_ru/n52 [0]}),
    .b({data_rd[53],\cu_ru/n52 [1]}),
    .c({data_rd[54],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[55],\cu_ru/n52 [3]}),
    .e({open_n84202,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c13_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c13_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c13_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c13_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c13_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c13_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_053 ,\cu_ru/al_ram_gpr_do_i1_052 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c13_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c13_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c13_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c13_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c13_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c13_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c13_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_055 ,\cu_ru/al_ram_gpr_do_i1_054 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c14_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c14_l  (
    .a({data_rd[56],\cu_ru/n52 [0]}),
    .b({data_rd[57],\cu_ru/n52 [1]}),
    .c({data_rd[58],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[59],\cu_ru/n52 [3]}),
    .e({open_n84237,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c14_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c14_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c14_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c14_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c14_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c14_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_057 ,\cu_ru/al_ram_gpr_do_i1_056 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c14_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c14_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c14_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c14_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c14_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c14_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c14_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_059 ,\cu_ru/al_ram_gpr_do_i1_058 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c15_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c15_l  (
    .a({data_rd[60],\cu_ru/n52 [0]}),
    .b({data_rd[61],\cu_ru/n52 [1]}),
    .c({data_rd[62],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[63],\cu_ru/n52 [3]}),
    .e({open_n84272,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c15_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c15_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c15_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c15_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c15_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c15_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_061 ,\cu_ru/al_ram_gpr_do_i1_060 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c15_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c15_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c15_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c15_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c15_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c15_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c15_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_063 ,\cu_ru/al_ram_gpr_do_i1_062 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c1_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c1_l  (
    .a({data_rd[4],\cu_ru/n52 [0]}),
    .b({data_rd[5],\cu_ru/n52 [1]}),
    .c({data_rd[6],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[7],\cu_ru/n52 [3]}),
    .e({open_n84307,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c1_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c1_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c1_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c1_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c1_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_005 ,\cu_ru/al_ram_gpr_do_i1_004 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c1_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c1_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c1_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c1_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c1_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c1_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c1_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_007 ,\cu_ru/al_ram_gpr_do_i1_006 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c2_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c2_l  (
    .a({data_rd[8],\cu_ru/n52 [0]}),
    .b({data_rd[9],\cu_ru/n52 [1]}),
    .c({data_rd[10],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[11],\cu_ru/n52 [3]}),
    .e({open_n84342,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c2_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c2_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c2_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c2_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c2_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_009 ,\cu_ru/al_ram_gpr_do_i1_008 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c2_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c2_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c2_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c2_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c2_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c2_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c2_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_011 ,\cu_ru/al_ram_gpr_do_i1_010 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c3_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c3_l  (
    .a({data_rd[12],\cu_ru/n52 [0]}),
    .b({data_rd[13],\cu_ru/n52 [1]}),
    .c({data_rd[14],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[15],\cu_ru/n52 [3]}),
    .e({open_n84377,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c3_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c3_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c3_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c3_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c3_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_013 ,\cu_ru/al_ram_gpr_do_i1_012 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c3_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c3_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c3_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c3_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c3_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c3_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c3_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_015 ,\cu_ru/al_ram_gpr_do_i1_014 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c4_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c4_l  (
    .a({data_rd[16],\cu_ru/n52 [0]}),
    .b({data_rd[17],\cu_ru/n52 [1]}),
    .c({data_rd[18],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[19],\cu_ru/n52 [3]}),
    .e({open_n84412,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c4_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c4_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c4_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c4_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c4_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_017 ,\cu_ru/al_ram_gpr_do_i1_016 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c4_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c4_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c4_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c4_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c4_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c4_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c4_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_019 ,\cu_ru/al_ram_gpr_do_i1_018 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c5_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c5_l  (
    .a({data_rd[20],\cu_ru/n52 [0]}),
    .b({data_rd[21],\cu_ru/n52 [1]}),
    .c({data_rd[22],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[23],\cu_ru/n52 [3]}),
    .e({open_n84447,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c5_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c5_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c5_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c5_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c5_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_021 ,\cu_ru/al_ram_gpr_do_i1_020 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c5_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c5_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c5_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c5_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c5_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c5_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c5_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_023 ,\cu_ru/al_ram_gpr_do_i1_022 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c6_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c6_l  (
    .a({data_rd[24],\cu_ru/n52 [0]}),
    .b({data_rd[25],\cu_ru/n52 [1]}),
    .c({data_rd[26],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[27],\cu_ru/n52 [3]}),
    .e({open_n84482,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c6_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c6_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c6_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c6_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c6_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_025 ,\cu_ru/al_ram_gpr_do_i1_024 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c6_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c6_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c6_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c6_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c6_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c6_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c6_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_027 ,\cu_ru/al_ram_gpr_do_i1_026 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c7_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c7_l  (
    .a({data_rd[28],\cu_ru/n52 [0]}),
    .b({data_rd[29],\cu_ru/n52 [1]}),
    .c({data_rd[30],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[31],\cu_ru/n52 [3]}),
    .e({open_n84517,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c7_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c7_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c7_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c7_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c7_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_029 ,\cu_ru/al_ram_gpr_do_i1_028 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c7_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c7_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c7_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c7_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c7_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c7_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c7_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_031 ,\cu_ru/al_ram_gpr_do_i1_030 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c8_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c8_l  (
    .a({data_rd[32],\cu_ru/n52 [0]}),
    .b({data_rd[33],\cu_ru/n52 [1]}),
    .c({data_rd[34],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[35],\cu_ru/n52 [3]}),
    .e({open_n84552,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c8_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c8_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c8_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c8_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c8_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c8_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_033 ,\cu_ru/al_ram_gpr_do_i1_032 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c8_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c8_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c8_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c8_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c8_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c8_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c8_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_035 ,\cu_ru/al_ram_gpr_do_i1_034 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c9_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \cu_ru/al_ram_gpr_r1_c9_l  (
    .a({data_rd[36],\cu_ru/n52 [0]}),
    .b({data_rd[37],\cu_ru/n52 [1]}),
    .c({data_rd[38],\cu_ru/n52 [2]}),
    .clk(clk_pad),
    .d({data_rd[39],\cu_ru/n52 [3]}),
    .e({open_n84587,\cu_ru/n53_1_al_n1986 }),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c9_di ),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c9_we ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c9_l"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c9_m0  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c9_di [1:0]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c9_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_037 ,\cu_ru/al_ram_gpr_do_i1_036 }));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/al_ram_gpr_r1_c9_l"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \cu_ru/al_ram_gpr_r1_c9_m1  (
    .a({\cu_ru/n46 [0],\cu_ru/n46 [0]}),
    .b({\cu_ru/n46 [1],\cu_ru/n46 [1]}),
    .c({\cu_ru/n46 [2],\cu_ru/n46 [2]}),
    .d({\cu_ru/n46 [3],\cu_ru/n46 [3]}),
    .dpram_di(\cu_ru/al_ram_gpr_r1_c9_di [3:2]),
    .dpram_mode(\cu_ru/al_ram_gpr_r1_c9_mode ),
    .dpram_waddr(\cu_ru/al_ram_gpr_r1_c9_waddr ),
    .dpram_wclk(\cu_ru/al_ram_gpr_r1_c9_wclk ),
    .dpram_we(\cu_ru/al_ram_gpr_r1_c9_we ),
    .f({\cu_ru/al_ram_gpr_do_i1_039 ,\cu_ru/al_ram_gpr_do_i1_038 }));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u11_al_u9772  (
    .a({\cu_ru/mcycle [13],\cu_ru/mcycle [11]}),
    .b({\cu_ru/mcycle [14],\cu_ru/mcycle [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c11 ),
    .f({\cu_ru/m_cycle_event/n2 [13],\cu_ru/m_cycle_event/n2 [11]}),
    .fco(\cu_ru/m_cycle_event/add0/c15 ),
    .fx({\cu_ru/m_cycle_event/n2 [14],\cu_ru/m_cycle_event/n2 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u15_al_u9773  (
    .a({\cu_ru/mcycle [17],\cu_ru/mcycle [15]}),
    .b({\cu_ru/mcycle [18],\cu_ru/mcycle [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c15 ),
    .f({\cu_ru/m_cycle_event/n2 [17],\cu_ru/m_cycle_event/n2 [15]}),
    .fco(\cu_ru/m_cycle_event/add0/c19 ),
    .fx({\cu_ru/m_cycle_event/n2 [18],\cu_ru/m_cycle_event/n2 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u19_al_u9774  (
    .a({\cu_ru/mcycle [21],\cu_ru/mcycle [19]}),
    .b({\cu_ru/mcycle [22],\cu_ru/mcycle [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c19 ),
    .f({\cu_ru/m_cycle_event/n2 [21],\cu_ru/m_cycle_event/n2 [19]}),
    .fco(\cu_ru/m_cycle_event/add0/c23 ),
    .fx({\cu_ru/m_cycle_event/n2 [22],\cu_ru/m_cycle_event/n2 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u23_al_u9775  (
    .a({\cu_ru/mcycle [25],\cu_ru/mcycle [23]}),
    .b({\cu_ru/mcycle [26],\cu_ru/mcycle [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c23 ),
    .f({\cu_ru/m_cycle_event/n2 [25],\cu_ru/m_cycle_event/n2 [23]}),
    .fco(\cu_ru/m_cycle_event/add0/c27 ),
    .fx({\cu_ru/m_cycle_event/n2 [26],\cu_ru/m_cycle_event/n2 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u27_al_u9776  (
    .a({\cu_ru/mcycle [29],\cu_ru/mcycle [27]}),
    .b({\cu_ru/mcycle [30],\cu_ru/mcycle [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c27 ),
    .f({\cu_ru/m_cycle_event/n2 [29],\cu_ru/m_cycle_event/n2 [27]}),
    .fco(\cu_ru/m_cycle_event/add0/c31 ),
    .fx({\cu_ru/m_cycle_event/n2 [30],\cu_ru/m_cycle_event/n2 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u31_al_u9777  (
    .a({\cu_ru/mcycle [33],\cu_ru/mcycle [31]}),
    .b({\cu_ru/mcycle [34],\cu_ru/mcycle [32]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c31 ),
    .f({\cu_ru/m_cycle_event/n2 [33],\cu_ru/m_cycle_event/n2 [31]}),
    .fco(\cu_ru/m_cycle_event/add0/c35 ),
    .fx({\cu_ru/m_cycle_event/n2 [34],\cu_ru/m_cycle_event/n2 [32]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u35_al_u9778  (
    .a({\cu_ru/mcycle [37],\cu_ru/mcycle [35]}),
    .b({\cu_ru/mcycle [38],\cu_ru/mcycle [36]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c35 ),
    .f({\cu_ru/m_cycle_event/n2 [37],\cu_ru/m_cycle_event/n2 [35]}),
    .fco(\cu_ru/m_cycle_event/add0/c39 ),
    .fx({\cu_ru/m_cycle_event/n2 [38],\cu_ru/m_cycle_event/n2 [36]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u39_al_u9779  (
    .a({\cu_ru/mcycle [41],\cu_ru/mcycle [39]}),
    .b({\cu_ru/mcycle [42],\cu_ru/mcycle [40]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c39 ),
    .f({\cu_ru/m_cycle_event/n2 [41],\cu_ru/m_cycle_event/n2 [39]}),
    .fco(\cu_ru/m_cycle_event/add0/c43 ),
    .fx({\cu_ru/m_cycle_event/n2 [42],\cu_ru/m_cycle_event/n2 [40]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u3_al_u9770  (
    .a({\cu_ru/mcycle [5],\cu_ru/mcycle [3]}),
    .b({\cu_ru/mcycle [6],\cu_ru/mcycle [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c3 ),
    .f({\cu_ru/m_cycle_event/n2 [5],\cu_ru/m_cycle_event/n2 [3]}),
    .fco(\cu_ru/m_cycle_event/add0/c7 ),
    .fx({\cu_ru/m_cycle_event/n2 [6],\cu_ru/m_cycle_event/n2 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u43_al_u9780  (
    .a({\cu_ru/mcycle [45],\cu_ru/mcycle [43]}),
    .b({\cu_ru/mcycle [46],\cu_ru/mcycle [44]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c43 ),
    .f({\cu_ru/m_cycle_event/n2 [45],\cu_ru/m_cycle_event/n2 [43]}),
    .fco(\cu_ru/m_cycle_event/add0/c47 ),
    .fx({\cu_ru/m_cycle_event/n2 [46],\cu_ru/m_cycle_event/n2 [44]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u47_al_u9781  (
    .a({\cu_ru/mcycle [49],\cu_ru/mcycle [47]}),
    .b({\cu_ru/mcycle [50],\cu_ru/mcycle [48]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c47 ),
    .f({\cu_ru/m_cycle_event/n2 [49],\cu_ru/m_cycle_event/n2 [47]}),
    .fco(\cu_ru/m_cycle_event/add0/c51 ),
    .fx({\cu_ru/m_cycle_event/n2 [50],\cu_ru/m_cycle_event/n2 [48]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u51_al_u9782  (
    .a({\cu_ru/mcycle [53],\cu_ru/mcycle [51]}),
    .b({\cu_ru/mcycle [54],\cu_ru/mcycle [52]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c51 ),
    .f({\cu_ru/m_cycle_event/n2 [53],\cu_ru/m_cycle_event/n2 [51]}),
    .fco(\cu_ru/m_cycle_event/add0/c55 ),
    .fx({\cu_ru/m_cycle_event/n2 [54],\cu_ru/m_cycle_event/n2 [52]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u55_al_u9783  (
    .a({\cu_ru/mcycle [57],\cu_ru/mcycle [55]}),
    .b({\cu_ru/mcycle [58],\cu_ru/mcycle [56]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c55 ),
    .f({\cu_ru/m_cycle_event/n2 [57],\cu_ru/m_cycle_event/n2 [55]}),
    .fco(\cu_ru/m_cycle_event/add0/c59 ),
    .fx({\cu_ru/m_cycle_event/n2 [58],\cu_ru/m_cycle_event/n2 [56]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u59_al_u9784  (
    .a({\cu_ru/mcycle [61],\cu_ru/mcycle [59]}),
    .b({\cu_ru/mcycle [62],\cu_ru/mcycle [60]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c59 ),
    .f({\cu_ru/m_cycle_event/n2 [61],\cu_ru/m_cycle_event/n2 [59]}),
    .fco(\cu_ru/m_cycle_event/add0/c63 ),
    .fx({\cu_ru/m_cycle_event/n2 [62],\cu_ru/m_cycle_event/n2 [60]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y8Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u63_al_u9785  (
    .a({open_n84873,\cu_ru/mcycle [63]}),
    .c(2'b00),
    .d({open_n84878,1'b0}),
    .fci(\cu_ru/m_cycle_event/add0/c63 ),
    .f({open_n84895,\cu_ru/m_cycle_event/n2 [63]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/u7_al_u9771  (
    .a({\cu_ru/mcycle [9],\cu_ru/mcycle [7]}),
    .b({\cu_ru/mcycle [10],\cu_ru/mcycle [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add0/c7 ),
    .f({\cu_ru/m_cycle_event/n2 [9],\cu_ru/m_cycle_event/n2 [7]}),
    .fco(\cu_ru/m_cycle_event/add0/c11 ),
    .fx({\cu_ru/m_cycle_event/n2 [10],\cu_ru/m_cycle_event/n2 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add0/ucin_al_u9769"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add0/ucin_al_u9769  (
    .a({\cu_ru/mcycle [1],1'b0}),
    .b({\cu_ru/mcycle [2],\cu_ru/mcycle [0]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\cu_ru/m_cycle_event/n2 [1],open_n84936}),
    .fco(\cu_ru/m_cycle_event/add0/c3 ),
    .fx({\cu_ru/m_cycle_event/n2 [2],\cu_ru/m_cycle_event/n2 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u11_al_u9789  (
    .a({\cu_ru/minstret [13],\cu_ru/minstret [11]}),
    .b({\cu_ru/minstret [14],\cu_ru/minstret [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c11 ),
    .f({\cu_ru/m_cycle_event/n4 [13],\cu_ru/m_cycle_event/n4 [11]}),
    .fco(\cu_ru/m_cycle_event/add1/c15 ),
    .fx({\cu_ru/m_cycle_event/n4 [14],\cu_ru/m_cycle_event/n4 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u15_al_u9790  (
    .a({\cu_ru/minstret [17],\cu_ru/minstret [15]}),
    .b({\cu_ru/minstret [18],\cu_ru/minstret [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c15 ),
    .f({\cu_ru/m_cycle_event/n4 [17],\cu_ru/m_cycle_event/n4 [15]}),
    .fco(\cu_ru/m_cycle_event/add1/c19 ),
    .fx({\cu_ru/m_cycle_event/n4 [18],\cu_ru/m_cycle_event/n4 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u19_al_u9791  (
    .a({\cu_ru/minstret [21],\cu_ru/minstret [19]}),
    .b({\cu_ru/minstret [22],\cu_ru/minstret [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c19 ),
    .f({\cu_ru/m_cycle_event/n4 [21],\cu_ru/m_cycle_event/n4 [19]}),
    .fco(\cu_ru/m_cycle_event/add1/c23 ),
    .fx({\cu_ru/m_cycle_event/n4 [22],\cu_ru/m_cycle_event/n4 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u23_al_u9792  (
    .a({\cu_ru/minstret [25],\cu_ru/minstret [23]}),
    .b({\cu_ru/minstret [26],\cu_ru/minstret [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c23 ),
    .f({\cu_ru/m_cycle_event/n4 [25],\cu_ru/m_cycle_event/n4 [23]}),
    .fco(\cu_ru/m_cycle_event/add1/c27 ),
    .fx({\cu_ru/m_cycle_event/n4 [26],\cu_ru/m_cycle_event/n4 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u27_al_u9793  (
    .a({\cu_ru/minstret [29],\cu_ru/minstret [27]}),
    .b({\cu_ru/minstret [30],\cu_ru/minstret [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c27 ),
    .f({\cu_ru/m_cycle_event/n4 [29],\cu_ru/m_cycle_event/n4 [27]}),
    .fco(\cu_ru/m_cycle_event/add1/c31 ),
    .fx({\cu_ru/m_cycle_event/n4 [30],\cu_ru/m_cycle_event/n4 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u31_al_u9794  (
    .a({\cu_ru/minstret [33],\cu_ru/minstret [31]}),
    .b({\cu_ru/minstret [34],\cu_ru/minstret [32]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c31 ),
    .f({\cu_ru/m_cycle_event/n4 [33],\cu_ru/m_cycle_event/n4 [31]}),
    .fco(\cu_ru/m_cycle_event/add1/c35 ),
    .fx({\cu_ru/m_cycle_event/n4 [34],\cu_ru/m_cycle_event/n4 [32]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u35_al_u9795  (
    .a({\cu_ru/minstret [37],\cu_ru/minstret [35]}),
    .b({\cu_ru/minstret [38],\cu_ru/minstret [36]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c35 ),
    .f({\cu_ru/m_cycle_event/n4 [37],\cu_ru/m_cycle_event/n4 [35]}),
    .fco(\cu_ru/m_cycle_event/add1/c39 ),
    .fx({\cu_ru/m_cycle_event/n4 [38],\cu_ru/m_cycle_event/n4 [36]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u39_al_u9796  (
    .a({\cu_ru/minstret [41],\cu_ru/minstret [39]}),
    .b({\cu_ru/minstret [42],\cu_ru/minstret [40]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c39 ),
    .f({\cu_ru/m_cycle_event/n4 [41],\cu_ru/m_cycle_event/n4 [39]}),
    .fco(\cu_ru/m_cycle_event/add1/c43 ),
    .fx({\cu_ru/m_cycle_event/n4 [42],\cu_ru/m_cycle_event/n4 [40]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u3_al_u9787  (
    .a({\cu_ru/minstret [5],\cu_ru/minstret [3]}),
    .b({\cu_ru/minstret [6],\cu_ru/minstret [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c3 ),
    .f({\cu_ru/m_cycle_event/n4 [5],\cu_ru/m_cycle_event/n4 [3]}),
    .fco(\cu_ru/m_cycle_event/add1/c7 ),
    .fx({\cu_ru/m_cycle_event/n4 [6],\cu_ru/m_cycle_event/n4 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u43_al_u9797  (
    .a({\cu_ru/minstret [45],\cu_ru/minstret [43]}),
    .b({\cu_ru/minstret [46],\cu_ru/minstret [44]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c43 ),
    .f({\cu_ru/m_cycle_event/n4 [45],\cu_ru/m_cycle_event/n4 [43]}),
    .fco(\cu_ru/m_cycle_event/add1/c47 ),
    .fx({\cu_ru/m_cycle_event/n4 [46],\cu_ru/m_cycle_event/n4 [44]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u47_al_u9798  (
    .a({\cu_ru/minstret [49],\cu_ru/minstret [47]}),
    .b({\cu_ru/minstret [50],\cu_ru/minstret [48]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c47 ),
    .f({\cu_ru/m_cycle_event/n4 [49],\cu_ru/m_cycle_event/n4 [47]}),
    .fco(\cu_ru/m_cycle_event/add1/c51 ),
    .fx({\cu_ru/m_cycle_event/n4 [50],\cu_ru/m_cycle_event/n4 [48]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u51_al_u9799  (
    .a({\cu_ru/minstret [53],\cu_ru/minstret [51]}),
    .b({\cu_ru/minstret [54],\cu_ru/minstret [52]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c51 ),
    .f({\cu_ru/m_cycle_event/n4 [53],\cu_ru/m_cycle_event/n4 [51]}),
    .fco(\cu_ru/m_cycle_event/add1/c55 ),
    .fx({\cu_ru/m_cycle_event/n4 [54],\cu_ru/m_cycle_event/n4 [52]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u55_al_u9800  (
    .a({\cu_ru/minstret [57],\cu_ru/minstret [55]}),
    .b({\cu_ru/minstret [58],\cu_ru/minstret [56]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c55 ),
    .f({\cu_ru/m_cycle_event/n4 [57],\cu_ru/m_cycle_event/n4 [55]}),
    .fco(\cu_ru/m_cycle_event/add1/c59 ),
    .fx({\cu_ru/m_cycle_event/n4 [58],\cu_ru/m_cycle_event/n4 [56]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u59_al_u9801  (
    .a({\cu_ru/minstret [61],\cu_ru/minstret [59]}),
    .b({\cu_ru/minstret [62],\cu_ru/minstret [60]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c59 ),
    .f({\cu_ru/m_cycle_event/n4 [61],\cu_ru/m_cycle_event/n4 [59]}),
    .fco(\cu_ru/m_cycle_event/add1/c63 ),
    .fx({\cu_ru/m_cycle_event/n4 [62],\cu_ru/m_cycle_event/n4 [60]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y8Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u63_al_u9802  (
    .a({open_n85191,\cu_ru/minstret [63]}),
    .c(2'b00),
    .d({open_n85196,1'b0}),
    .fci(\cu_ru/m_cycle_event/add1/c63 ),
    .f({open_n85213,\cu_ru/m_cycle_event/n4 [63]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_cycle_event/add1/u7_al_u9788  (
    .a({\cu_ru/minstret [9],\cu_ru/minstret [7]}),
    .b({\cu_ru/minstret [10],\cu_ru/minstret [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_cycle_event/add1/c7 ),
    .f({\cu_ru/m_cycle_event/n4 [9],\cu_ru/m_cycle_event/n4 [7]}),
    .fco(\cu_ru/m_cycle_event/add1/c11 ),
    .fx({\cu_ru/m_cycle_event/n4 [10],\cu_ru/m_cycle_event/n4 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_cycle_event/add1/ucin_al_u9786"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/add1/ucin_al_u9786  (
    .a({\cu_ru/minstret [1],1'b0}),
    .b({\cu_ru/minstret [2],\cu_ru/minstret [0]}),
    .c(2'b00),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d(2'b01),
    .e(2'b01),
    .mi(\cu_ru/m_cycle_event/n4 [2:1]),
    .sr(rst_pad),
    .f({\cu_ru/m_cycle_event/n4 [1],open_n85249}),
    .fco(\cu_ru/m_cycle_event/add1/c3 ),
    .fx({\cu_ru/m_cycle_event/n4 [2],\cu_ru/m_cycle_event/n4 [0]}),
    .q(\cu_ru/minstret [2:1]));
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(51)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(51)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/cy_reg|cu_ru/m_cycle_event/ir_reg  (
    .a({open_n85250,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({_al_u3198_o,\cu_ru/trap_target_m }),
    .c({_al_u3184_o,\cu_ru/mepc [2]}),
    .ce(\cu_ru/m_cycle_event/n13 ),
    .clk(clk_pad),
    .d({_al_u3195_o,data_csr[2]}),
    .mi({data_csr[0],data_csr[2]}),
    .sr(rst_pad),
    .f({\cu_ru/m_cycle_event/n13 ,_al_u6652_o}),
    .q({\cu_ru/mcountinhibit ,\cu_ru/m_cycle_event/mcountinhibit[2] }));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(51)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(B*~(C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/reg0_b16|cu_ru/m_cycle_event/reg0_b55  (
    .a({open_n85264,_al_u6763_o}),
    .b({_al_u7131_o,\cu_ru/read_stval_sel_lutinv }),
    .c({\cu_ru/minstret [16],\cu_ru/minstret [55]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u6763_o,\cu_ru/stval [55]}),
    .mi({\cu_ru/m_cycle_event/n4 [16],\cu_ru/m_cycle_event/n4 [55]}),
    .sr(rst_pad),
    .f({_al_u7132_o,_al_u6829_o}),
    .q({\cu_ru/minstret [16],\cu_ru/minstret [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/reg0_b18|cu_ru/m_cycle_event/reg0_b34  (
    .a({_al_u6763_o,_al_u6763_o}),
    .b({\cu_ru/read_sepc_sel_lutinv ,\cu_ru/read_sepc_sel_lutinv }),
    .c({\cu_ru/minstret [18],\cu_ru/minstret [34]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/sepc [18],\cu_ru/sepc [34]}),
    .mi({\cu_ru/m_cycle_event/n4 [18],\cu_ru/m_cycle_event/n4 [34]}),
    .sr(rst_pad),
    .f({_al_u7631_o,_al_u7234_o}),
    .q({\cu_ru/minstret [18],\cu_ru/minstret [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/reg0_b19|cu_ru/m_cycle_event/reg0_b22  (
    .a({\cu_ru/read_instret_sel_lutinv ,\cu_ru/read_instret_sel_lutinv }),
    .b({\cu_ru/n64 [32],\cu_ru/read_mscratch_sel_lutinv }),
    .c({\cu_ru/minstret [19],\cu_ru/minstret [22]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({mxr,\cu_ru/mscratch [22]}),
    .mi({\cu_ru/m_cycle_event/n4 [19],\cu_ru/m_cycle_event/n4 [22]}),
    .sr(rst_pad),
    .f({_al_u7452_o,_al_u7609_o}),
    .q({\cu_ru/minstret [19],\cu_ru/minstret [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~D))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(B*~(C*~D))"),
    //.LUTG1("(B*~(C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110000001100),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b1100110000001100),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/reg0_b27|cu_ru/m_cycle_event/reg0_b58  (
    .b({_al_u7088_o,_al_u6794_o}),
    .c({\cu_ru/minstret [27],\cu_ru/minstret [58]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u6763_o,_al_u6763_o}),
    .mi({\cu_ru/m_cycle_event/n4 [27],\cu_ru/m_cycle_event/n4 [58]}),
    .sr(rst_pad),
    .f({_al_u7089_o,_al_u6795_o}),
    .q({\cu_ru/minstret [27],\cu_ru/minstret [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/reg0_b28|cu_ru/m_cycle_event/reg0_b45  (
    .a({_al_u6763_o,_al_u6763_o}),
    .b({\cu_ru/read_mtval_sel_lutinv ,\cu_ru/read_mtval_sel_lutinv }),
    .c({\cu_ru/minstret [28],\cu_ru/minstret [45]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtval [28],\cu_ru/mtval [45]}),
    .mi({\cu_ru/m_cycle_event/n4 [28],\cu_ru/m_cycle_event/n4 [45]}),
    .sr(rst_pad),
    .f({_al_u7444_o,_al_u6919_o}),
    .q({\cu_ru/minstret [28],\cu_ru/minstret [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(B*~(C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/reg0_b29|cu_ru/m_cycle_event/reg0_b44  (
    .b({_al_u7078_o,_al_u6926_o}),
    .c({\cu_ru/minstret [29],\cu_ru/minstret [44]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u6763_o,_al_u6763_o}),
    .mi({\cu_ru/m_cycle_event/n4 [29],\cu_ru/m_cycle_event/n4 [44]}),
    .sr(rst_pad),
    .f({_al_u7079_o,_al_u6927_o}),
    .q({\cu_ru/minstret [29],\cu_ru/minstret [44]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~D))"),
    //.LUT1("(B*~(C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110000001100),
    .INIT_LUT1(16'b1100110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/reg0_b31|cu_ru/m_cycle_event/reg0_b37  (
    .b({_al_u7068_o,_al_u7048_o}),
    .c({\cu_ru/minstret [31],\cu_ru/minstret [37]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u6763_o,_al_u6763_o}),
    .mi({\cu_ru/m_cycle_event/n4 [31],\cu_ru/m_cycle_event/n4 [37]}),
    .sr(rst_pad),
    .f({_al_u7069_o,_al_u7049_o}),
    .q({\cu_ru/minstret [31],\cu_ru/minstret [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*B)*~(C*~A))"),
    //.LUTF1("(~(D*B)*~(C*~A))"),
    //.LUTG0("(~(D*B)*~(C*~A))"),
    //.LUTG1("(~(D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001110101111),
    .INIT_LUTF1(16'b0010001110101111),
    .INIT_LUTG0(16'b0010001110101111),
    .INIT_LUTG1(16'b0010001110101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/reg0_b48|cu_ru/m_cycle_event/reg0_b57  (
    .a({_al_u6763_o,_al_u6763_o}),
    .b({\cu_ru/read_stval_sel_lutinv ,\cu_ru/read_stval_sel_lutinv }),
    .c({\cu_ru/minstret [48],\cu_ru/minstret [57]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/stval [48],\cu_ru/stval [57]}),
    .mi({\cu_ru/m_cycle_event/n4 [48],\cu_ru/m_cycle_event/n4 [57]}),
    .sr(rst_pad),
    .f({_al_u6897_o,_al_u6810_o}),
    .q({\cu_ru/minstret [48],\cu_ru/minstret [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/reg0_b50|cu_ru/m_cycle_event/reg0_b56  (
    .a({_al_u6763_o,_al_u6763_o}),
    .b({\cu_ru/read_stval_sel_lutinv ,\cu_ru/read_stval_sel_lutinv }),
    .c({\cu_ru/minstret [50],\cu_ru/minstret [56]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/stval [50],\cu_ru/stval [56]}),
    .mi({\cu_ru/m_cycle_event/n4 [50],\cu_ru/m_cycle_event/n4 [56]}),
    .sr(rst_pad),
    .f({_al_u6870_o,_al_u6812_o}),
    .q({\cu_ru/minstret [50],\cu_ru/minstret [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*~A))"),
    //.LUT1("(~(D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001110101111),
    .INIT_LUT1(16'b0010001110101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_cycle_event/reg0_b6|cu_ru/m_cycle_event/reg0_b9  (
    .a({_al_u6763_o,_al_u6763_o}),
    .b({\cu_ru/read_mtvec_sel_lutinv ,\cu_ru/read_mtvec_sel_lutinv }),
    .c({\cu_ru/minstret [6],\cu_ru/minstret [9]}),
    .ce(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/mtvec [6],\cu_ru/mtvec [9]}),
    .mi({\cu_ru/m_cycle_event/n4 [6],\cu_ru/m_cycle_event/n4 [9]}),
    .sr(rst_pad),
    .f({_al_u7348_o,_al_u7812_o}),
    .q({\cu_ru/minstret [6],\cu_ru/minstret [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b10|cu_ru/m_s_cause/reg1_b6  (
    .a({open_n85409,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({open_n85410,\cu_ru/trap_target_m }),
    .c({_al_u3206_o,\cu_ru/mtval [6]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u5992_o,data_csr[6]}),
    .mi({data_csr[10],data_csr[6]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ,_al_u6447_o}),
    .q({\cu_ru/mcause [10],\cu_ru/mcause [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b11|cu_ru/m_s_cause/reg1_b9  (
    .a({open_n85424,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/mcause [1],\cu_ru/trap_target_m }),
    .c({data_csr[1],\cu_ru/mtval [9]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ,data_csr[9]}),
    .mi({data_csr[11],data_csr[9]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u7335_o,_al_u6441_o}),
    .q({\cu_ru/mcause [11],\cu_ru/mcause [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b12|cu_ru/m_s_cause/reg1_b7  (
    .a({open_n85442,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/mcause [3],\cu_ru/trap_target_m }),
    .c({data_csr[3],\cu_ru/mtval [7]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ,data_csr[7]}),
    .mi({data_csr[12],data_csr[7]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6727_o,_al_u6445_o}),
    .q({\cu_ru/mcause [12],\cu_ru/mcause [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b13|cu_ru/m_s_cause/reg1_b8  (
    .a({\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mcause [0],\cu_ru/mtval [8]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[0],data_csr[8]}),
    .mi({data_csr[13],data_csr[8]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6702_o,_al_u6443_o}),
    .q({\cu_ru/mcause [13],\cu_ru/mcause [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b14|cu_ru/m_s_cause/reg1_b4  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [14],\cu_ru/mtval [4]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[14],data_csr[4]}),
    .mi({data_csr[14],data_csr[4]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6557_o,_al_u6479_o}),
    .q({\cu_ru/mcause [14],\cu_ru/mcause [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b15|cu_ru/m_s_cause/reg1_b21  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [15],\cu_ru/mtval [21]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[15],data_csr[21]}),
    .mi({data_csr[15],data_csr[21]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6555_o,_al_u6541_o}),
    .q({\cu_ru/mcause [15],\cu_ru/mcause [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b16|cu_ru/m_s_cause/reg1_b20  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [16],\cu_ru/mtval [20]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[16],data_csr[20]}),
    .mi({data_csr[16],data_csr[20]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6553_o,_al_u6543_o}),
    .q({\cu_ru/mcause [16],\cu_ru/mcause [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b17|cu_ru/m_s_cause/reg1_b19  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [17],\cu_ru/mtval [19]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[17],data_csr[19]}),
    .mi({data_csr[17],data_csr[19]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6551_o,_al_u6547_o}),
    .q({\cu_ru/mcause [17],\cu_ru/mcause [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b23|cu_ru/m_s_cause/reg1_b62  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [23],\cu_ru/mtval [62]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[23],data_csr[62]}),
    .mi({data_csr[23],data_csr[62]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6537_o,_al_u6451_o}),
    .q({\cu_ru/mcause [23],\cu_ru/mcause [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b24|cu_ru/m_s_cause/reg1_b60  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [24],\cu_ru/mtval [60]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[24],data_csr[60]}),
    .mi({data_csr[24],data_csr[60]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6535_o,_al_u6455_o}),
    .q({\cu_ru/mcause [24],\cu_ru/mcause [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b25|cu_ru/m_s_cause/reg1_b42  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [25],\cu_ru/mtval [42]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[25],data_csr[42]}),
    .mi({data_csr[25],data_csr[42]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6533_o,_al_u6495_o}),
    .q({\cu_ru/mcause [25],\cu_ru/mcause [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b26|cu_ru/m_s_cause/reg1_b41  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [26],\cu_ru/mtval [41]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[26],data_csr[41]}),
    .mi({data_csr[26],data_csr[41]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6531_o,_al_u6497_o}),
    .q({\cu_ru/mcause [26],\cu_ru/mcause [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b27|cu_ru/m_s_cause/reg1_b40  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [27],\cu_ru/mtval [40]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[27],data_csr[40]}),
    .mi({data_csr[27],data_csr[40]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6529_o,_al_u6499_o}),
    .q({\cu_ru/mcause [27],\cu_ru/mcause [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b28|cu_ru/m_s_cause/reg1_b39  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [28],\cu_ru/mtval [39]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[28],data_csr[39]}),
    .mi({data_csr[28],data_csr[39]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6527_o,_al_u6503_o}),
    .q({\cu_ru/mcause [28],\cu_ru/mcause [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b29|cu_ru/m_s_cause/reg1_b38  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [29],\cu_ru/mtval [38]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[29],data_csr[38]}),
    .mi({data_csr[29],data_csr[38]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6525_o,_al_u6505_o}),
    .q({\cu_ru/mcause [29],\cu_ru/mcause [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b30|cu_ru/m_s_cause/reg1_b37  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [30],\cu_ru/mtval [37]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[30],data_csr[37]}),
    .mi({data_csr[30],data_csr[37]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6521_o,_al_u6507_o}),
    .q({\cu_ru/mcause [30],\cu_ru/mcause [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b31|cu_ru/m_s_cause/reg1_b36  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [31],\cu_ru/mtval [36]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[31],data_csr[36]}),
    .mi({data_csr[31],data_csr[36]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6519_o,_al_u6509_o}),
    .q({\cu_ru/mcause [31],\cu_ru/mcause [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b32|cu_ru/m_s_cause/reg1_b35  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [32],\cu_ru/mtval [35]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[32],data_csr[35]}),
    .mi({data_csr[32],data_csr[35]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6517_o,_al_u6511_o}),
    .q({\cu_ru/mcause [32],\cu_ru/mcause [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b44|cu_ru/m_s_cause/reg1_b33  (
    .a({\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [44],\cu_ru/mtval [33]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[44],data_csr[33]}),
    .mi({data_csr[44],data_csr[33]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6620_o,_al_u6515_o}),
    .q({\cu_ru/mcause [44],\cu_ru/mcause [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \cu_ru/m_s_cause/reg1_b45|cu_ru/m_s_cause/reg1_b58  (
    .a({\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ,\cu_ru/m_s_epc/mux6_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mepc [45],\cu_ru/mepc [58]}),
    .ce(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({data_csr[45],data_csr[58]}),
    .mi({data_csr[45],data_csr[58]}),
    .sr(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .f({_al_u6618_o,_al_u6590_o}),
    .q({\cu_ru/mcause [45],\cu_ru/mcause [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u11_al_u9840  (
    .a({wb_ins_pc[15],wb_ins_pc[13]}),
    .b({wb_ins_pc[16],wb_ins_pc[14]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c11 ),
    .f({\cu_ru/m_s_epc/n0 [13],\cu_ru/m_s_epc/n0 [11]}),
    .fco(\cu_ru/m_s_epc/add0/c15 ),
    .fx({\cu_ru/m_s_epc/n0 [14],\cu_ru/m_s_epc/n0 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u15_al_u9841  (
    .a({wb_ins_pc[19],wb_ins_pc[17]}),
    .b({wb_ins_pc[20],wb_ins_pc[18]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c15 ),
    .f({\cu_ru/m_s_epc/n0 [17],\cu_ru/m_s_epc/n0 [15]}),
    .fco(\cu_ru/m_s_epc/add0/c19 ),
    .fx({\cu_ru/m_s_epc/n0 [18],\cu_ru/m_s_epc/n0 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u19_al_u9842  (
    .a({wb_ins_pc[23],wb_ins_pc[21]}),
    .b({wb_ins_pc[24],wb_ins_pc[22]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c19 ),
    .f({\cu_ru/m_s_epc/n0 [21],\cu_ru/m_s_epc/n0 [19]}),
    .fco(\cu_ru/m_s_epc/add0/c23 ),
    .fx({\cu_ru/m_s_epc/n0 [22],\cu_ru/m_s_epc/n0 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u23_al_u9843  (
    .a({wb_ins_pc[27],wb_ins_pc[25]}),
    .b({wb_ins_pc[28],wb_ins_pc[26]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c23 ),
    .f({\cu_ru/m_s_epc/n0 [25],\cu_ru/m_s_epc/n0 [23]}),
    .fco(\cu_ru/m_s_epc/add0/c27 ),
    .fx({\cu_ru/m_s_epc/n0 [26],\cu_ru/m_s_epc/n0 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u27_al_u9844  (
    .a({wb_ins_pc[31],wb_ins_pc[29]}),
    .b({wb_ins_pc[32],wb_ins_pc[30]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c27 ),
    .f({\cu_ru/m_s_epc/n0 [29],\cu_ru/m_s_epc/n0 [27]}),
    .fco(\cu_ru/m_s_epc/add0/c31 ),
    .fx({\cu_ru/m_s_epc/n0 [30],\cu_ru/m_s_epc/n0 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u31_al_u9845  (
    .a({wb_ins_pc[35],wb_ins_pc[33]}),
    .b({wb_ins_pc[36],wb_ins_pc[34]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c31 ),
    .f({\cu_ru/m_s_epc/n0 [33],\cu_ru/m_s_epc/n0 [31]}),
    .fco(\cu_ru/m_s_epc/add0/c35 ),
    .fx({\cu_ru/m_s_epc/n0 [34],\cu_ru/m_s_epc/n0 [32]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u35_al_u9846  (
    .a({wb_ins_pc[39],wb_ins_pc[37]}),
    .b({wb_ins_pc[40],wb_ins_pc[38]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c35 ),
    .f({\cu_ru/m_s_epc/n0 [37],\cu_ru/m_s_epc/n0 [35]}),
    .fco(\cu_ru/m_s_epc/add0/c39 ),
    .fx({\cu_ru/m_s_epc/n0 [38],\cu_ru/m_s_epc/n0 [36]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u39_al_u9847  (
    .a({wb_ins_pc[43],wb_ins_pc[41]}),
    .b({wb_ins_pc[44],wb_ins_pc[42]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c39 ),
    .f({\cu_ru/m_s_epc/n0 [41],\cu_ru/m_s_epc/n0 [39]}),
    .fco(\cu_ru/m_s_epc/add0/c43 ),
    .fx({\cu_ru/m_s_epc/n0 [42],\cu_ru/m_s_epc/n0 [40]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u3_al_u9838  (
    .a({wb_ins_pc[7],wb_ins_pc[5]}),
    .b({wb_ins_pc[8],wb_ins_pc[6]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c3 ),
    .f({\cu_ru/m_s_epc/n0 [5],\cu_ru/m_s_epc/n0 [3]}),
    .fco(\cu_ru/m_s_epc/add0/c7 ),
    .fx({\cu_ru/m_s_epc/n0 [6],\cu_ru/m_s_epc/n0 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u43_al_u9848  (
    .a({wb_ins_pc[47],wb_ins_pc[45]}),
    .b({wb_ins_pc[48],wb_ins_pc[46]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c43 ),
    .f({\cu_ru/m_s_epc/n0 [45],\cu_ru/m_s_epc/n0 [43]}),
    .fco(\cu_ru/m_s_epc/add0/c47 ),
    .fx({\cu_ru/m_s_epc/n0 [46],\cu_ru/m_s_epc/n0 [44]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u47_al_u9849  (
    .a({wb_ins_pc[51],wb_ins_pc[49]}),
    .b({wb_ins_pc[52],wb_ins_pc[50]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c47 ),
    .f({\cu_ru/m_s_epc/n0 [49],\cu_ru/m_s_epc/n0 [47]}),
    .fco(\cu_ru/m_s_epc/add0/c51 ),
    .fx({\cu_ru/m_s_epc/n0 [50],\cu_ru/m_s_epc/n0 [48]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u51_al_u9850  (
    .a({wb_ins_pc[55],wb_ins_pc[53]}),
    .b({wb_ins_pc[56],wb_ins_pc[54]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c51 ),
    .f({\cu_ru/m_s_epc/n0 [53],\cu_ru/m_s_epc/n0 [51]}),
    .fco(\cu_ru/m_s_epc/add0/c55 ),
    .fx({\cu_ru/m_s_epc/n0 [54],\cu_ru/m_s_epc/n0 [52]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u55_al_u9851  (
    .a({wb_ins_pc[59],wb_ins_pc[57]}),
    .b({wb_ins_pc[60],wb_ins_pc[58]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c55 ),
    .f({\cu_ru/m_s_epc/n0 [57],\cu_ru/m_s_epc/n0 [55]}),
    .fco(\cu_ru/m_s_epc/add0/c59 ),
    .fx({\cu_ru/m_s_epc/n0 [58],\cu_ru/m_s_epc/n0 [56]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u59_al_u9852  (
    .a({wb_ins_pc[63],wb_ins_pc[61]}),
    .b({open_n85943,wb_ins_pc[62]}),
    .c(2'b00),
    .d(2'b00),
    .e({open_n85946,1'b0}),
    .fci(\cu_ru/m_s_epc/add0/c59 ),
    .f({\cu_ru/m_s_epc/n0 [61],\cu_ru/m_s_epc/n0 [59]}),
    .fx({open_n85962,\cu_ru/m_s_epc/n0 [60]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \cu_ru/m_s_epc/add0/u7_al_u9839  (
    .a({wb_ins_pc[11],wb_ins_pc[9]}),
    .b({wb_ins_pc[12],wb_ins_pc[10]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\cu_ru/m_s_epc/add0/c7 ),
    .f({\cu_ru/m_s_epc/n0 [9],\cu_ru/m_s_epc/n0 [7]}),
    .fco(\cu_ru/m_s_epc/add0/c11 ),
    .fx({\cu_ru/m_s_epc/n0 [10],\cu_ru/m_s_epc/n0 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("cu_ru/m_s_epc/add0/ucin_al_u9837"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_epc/add0/ucin_al_u9837  (
    .a({wb_ins_pc[3],1'b0}),
    .b({wb_ins_pc[4],wb_ins_pc[2]}),
    .c(2'b00),
    .clk(clk_pad),
    .d(2'b01),
    .e(2'b01),
    .mi(ex_ins_pc[3:2]),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n0 [1],open_n85996}),
    .fco(\cu_ru/m_s_epc/add0/c3 ),
    .fx({\cu_ru/m_s_epc/n0 [2],\cu_ru/m_s_epc/n0 [0]}),
    .q(wb_ins_pc[3:2]));
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IDDRPIPEMODE("NONE"),
    .INCEMUX("INV"),
    .INPCLKMUX("CLK"),
    .INRSTMUX("RST"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("RESET"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .SRMODE("SYNC"),
    .TSMUX("1"))
    \cu_ru/m_s_ip/meip_reg_IN  (
    .ce(\cu_ru/m_s_ip/u12_sel_is_2_o ),
    .ipad(m_ext_int),
    .ipclk(clk_pad),
    .rst(rst_pad),
    .diq({open_n86006,open_n86007,open_n86008,\cu_ru/m_sip [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IDDRPIPEMODE("NONE"),
    .INCEMUX("INV"),
    .INPCLKMUX("CLK"),
    .INRSTMUX("RST"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("RESET"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .SRMODE("SYNC"),
    .TSMUX("1"))
    \cu_ru/m_s_ip/msip_reg_IN  (
    .ce(\cu_ru/m_s_ip/u12_sel_is_2_o ),
    .ipad(m_soft_int),
    .ipclk(clk_pad),
    .rst(rst_pad),
    .diq({open_n86020,open_n86021,open_n86022,\cu_ru/m_sip [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IDDRPIPEMODE("NONE"),
    .INCEMUX("INV"),
    .INPCLKMUX("CLK"),
    .INRSTMUX("RST"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("RESET"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .SRMODE("SYNC"),
    .TSMUX("1"))
    \cu_ru/m_s_ip/mtip_reg_IN  (
    .ce(\cu_ru/m_s_ip/u12_sel_is_2_o ),
    .ipad(m_time_int),
    .ipclk(clk_pad),
    .rst(rst_pad),
    .diq({open_n86034,open_n86035,open_n86036,\cu_ru/m_sip [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_ip/seip_reg|cu_ru/m_s_ip/stip_reg  (
    .c({data_csr[9],_al_u3191_o}),
    .ce(\cu_ru/m_s_ip/n0 ),
    .clk(clk_pad),
    .d({s_ext_int_pad,_al_u3190_o}),
    .mi({open_n86046,data_csr[5]}),
    .sr(rst_pad),
    .f({open_n86058,\cu_ru/m_s_ip/n0 }),
    .q({\cu_ru/m_s_ip/seip ,\cu_ru/m_sip [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg0_b0|cu_ru/m_s_scratch/reg0_b47  (
    .a({open_n86062,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({open_n86063,\cu_ru/trap_target_m }),
    .c({_al_u3190_o,\cu_ru/mtval [47]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({_al_u3185_o,data_csr[47]}),
    .mi({data_csr[0],data_csr[47]}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_scratch/n0 ,_al_u6485_o}),
    .q({\cu_ru/mscratch [0],\cu_ru/mscratch [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg0_b44|cu_ru/m_s_scratch/reg0_b59  (
    .a({\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux5_b0_sel_is_2_o }),
    .b({\cu_ru/trap_target_m ,\cu_ru/trap_target_m }),
    .c({\cu_ru/mtval [44],\cu_ru/mtval [59]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({data_csr[44],data_csr[59]}),
    .mi({data_csr[44],data_csr[59]}),
    .sr(rst_pad),
    .f({_al_u6491_o,_al_u6459_o}),
    .q({\cu_ru/mscratch [44],\cu_ru/mscratch [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg0_b7|cu_ru/m_s_scratch/reg0_b5  (
    .b({\cu_ru/stval [7],\cu_ru/stval [5]}),
    .c({data_csr[7],data_csr[5]}),
    .ce(\cu_ru/m_s_scratch/n0 ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[7],data_csr[5]}),
    .sr(rst_pad),
    .f({_al_u5167_o,_al_u5215_o}),
    .q({\cu_ru/mscratch [7],\cu_ru/mscratch [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b0|cu_ru/m_s_scratch/reg1_b6  (
    .b({open_n86115,\cu_ru/stval [6]}),
    .c({_al_u3420_o,data_csr[6]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({_al_u3185_o,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[0],data_csr[6]}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ,_al_u5182_o}),
    .q({\cu_ru/sscratch [0],\cu_ru/sscratch [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b14|cu_ru/m_s_scratch/reg1_b9  (
    .b({\cu_ru/stval [14],\cu_ru/stval [9]}),
    .c({data_csr[14],data_csr[9]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[14],data_csr[9]}),
    .sr(rst_pad),
    .f({_al_u5332_o,_al_u5160_o}),
    .q({\cu_ru/sscratch [14],\cu_ru/sscratch [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b15|cu_ru/m_s_scratch/reg1_b4  (
    .b({\cu_ru/stval [15],\cu_ru/stval [4]}),
    .c({data_csr[15],data_csr[4]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[15],data_csr[4]}),
    .sr(rst_pad),
    .f({_al_u5329_o,_al_u5248_o}),
    .q({\cu_ru/sscratch [15],\cu_ru/sscratch [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b16|cu_ru/m_s_scratch/reg1_b18  (
    .b({\cu_ru/stval [16],\cu_ru/stval [18]}),
    .c({data_csr[16],data_csr[18]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[16],data_csr[18]}),
    .sr(rst_pad),
    .f({_al_u5326_o,_al_u5320_o}),
    .q({\cu_ru/sscratch [16],\cu_ru/sscratch [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b23|cu_ru/m_s_scratch/reg1_b61  (
    .b({\cu_ru/stval [23],\cu_ru/stval [61]}),
    .c({data_csr[23],data_csr[61]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[23],data_csr[61]}),
    .sr(rst_pad),
    .f({_al_u5302_o,_al_u5176_o}),
    .q({\cu_ru/sscratch [23],\cu_ru/sscratch [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b24|cu_ru/m_s_scratch/reg1_b60  (
    .b({\cu_ru/stval [24],\cu_ru/stval [60]}),
    .c({data_csr[24],data_csr[60]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[24],data_csr[60]}),
    .sr(rst_pad),
    .f({_al_u5299_o,_al_u5179_o}),
    .q({\cu_ru/sscratch [24],\cu_ru/sscratch [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b25|cu_ru/m_s_scratch/reg1_b42  (
    .b({\cu_ru/stval [25],\cu_ru/stval [42]}),
    .c({data_csr[25],data_csr[42]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[25],data_csr[42]}),
    .sr(rst_pad),
    .f({_al_u5296_o,_al_u5239_o}),
    .q({\cu_ru/sscratch [25],\cu_ru/sscratch [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b26|cu_ru/m_s_scratch/reg1_b38  (
    .b({\cu_ru/stval [26],\cu_ru/stval [38]}),
    .c({data_csr[26],data_csr[38]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[26],data_csr[38]}),
    .sr(rst_pad),
    .f({_al_u5293_o,_al_u5254_o}),
    .q({\cu_ru/sscratch [26],\cu_ru/sscratch [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b27|cu_ru/m_s_scratch/reg1_b34  (
    .b({\cu_ru/stval [27],\cu_ru/stval [34]}),
    .c({data_csr[27],data_csr[34]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[27],data_csr[34]}),
    .sr(rst_pad),
    .f({_al_u5290_o,_al_u5266_o}),
    .q({\cu_ru/sscratch [27],\cu_ru/sscratch [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b28|cu_ru/m_s_scratch/reg1_b32  (
    .b({\cu_ru/stval [28],\cu_ru/stval [32]}),
    .c({data_csr[28],data_csr[32]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[28],data_csr[32]}),
    .sr(rst_pad),
    .f({_al_u5287_o,_al_u5272_o}),
    .q({\cu_ru/sscratch [28],\cu_ru/sscratch [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_scratch/reg1_b29|cu_ru/m_s_scratch/reg1_b30  (
    .b({\cu_ru/stval [29],\cu_ru/stval [30]}),
    .c({data_csr[29],data_csr[30]}),
    .ce(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ,\cu_ru/m_s_tval/mux3_b0_sel_is_2_o }),
    .mi({data_csr[29],data_csr[30]}),
    .sr(rst_pad),
    .f({_al_u5284_o,_al_u5278_o}),
    .q({\cu_ru/sscratch [29],\cu_ru/sscratch [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*B)*~(C*A))"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001001101011111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_status/mprv_reg|cu_ru/m_s_status/tsr_reg  (
    .a({open_n86299,\cu_ru/read_minstret_sel_lutinv }),
    .b({open_n86300,\cu_ru/n90 [32]}),
    .c({_al_u3195_o,\cu_ru/minstret [22]}),
    .ce(\cu_ru/m_s_status/n0 ),
    .clk(clk_pad),
    .d({_al_u3185_o,tsr}),
    .mi({data_csr[17],data_csr[22]}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_status/n0 ,_al_u7602_o}),
    .q({mprv,tsr}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  EG_PHY_MSLICE #(
    //.LUT0("~(~(D*~B)*~(C*A))"),
    //.LUT1("~(~B*~(~C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011001110100000),
    .INIT_LUT1(16'b1100111111001100),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_status/reg1_b1|cu_ru/m_s_status/reg1_b3  (
    .a({open_n86314,_al_u2841_o}),
    .b({_al_u2845_o,_al_u2842_o}),
    .c({\cu_ru/mstatus [12],\cu_ru/mstatus [12]}),
    .clk(clk_pad),
    .d({_al_u2841_o,priv[3]}),
    .sr(rst_pad),
    .q({priv[1],priv[3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_status/tvm_reg  (
    .ce(\cu_ru/m_s_status/n0 ),
    .clk(clk_pad),
    .mi({open_n86351,data_csr[20]}),
    .sr(rst_pad),
    .q({open_n86357,tvm}));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000001001100),
    .INIT_LUTF1(16'b0100000001001100),
    .INIT_LUTG0(16'b0100000001001100),
    .INIT_LUTG1(16'b0100000001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_tvec/reg0_b10|cu_ru/m_s_tvec/reg0_b3  (
    .a({csr_data[10],csr_data[3]}),
    .b({_al_u7141_o,_al_u7141_o}),
    .c({id_system,id_system}),
    .ce(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .clk(clk_pad),
    .d({id_ins_pc[10],id_ins_pc[3]}),
    .mi({csr_data[10],csr_data[3]}),
    .sr(rst_pad),
    .f({_al_u7710_o,_al_u7840_o}),
    .q({\cu_ru/stvec [10],\cu_ru/stvec [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*B*D)"),
    //.LUT1("~(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111111111111),
    .INIT_LUT1(16'b0011111111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \cu_ru/m_s_tvec/reg1_b13|cu_ru/m_s_tvec/reg1_b32  (
    .b({_al_u7282_o,_al_u7421_o}),
    .c({_al_u7283_o,_al_u7422_o}),
    .ce(\cu_ru/m_s_tvec/n0 ),
    .clk(clk_pad),
    .d({_al_u7281_o,_al_u7420_o}),
    .sr(rst_pad),
    .f({csr_data[13],csr_data[32]}),
    .q({\cu_ru/mtvec [13],\cu_ru/mtvec [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/sub0/u0|cu_ru/sub0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \cu_ru/sub0/u0|cu_ru/sub0/ucin  (
    .a({id_rs1_index[0],1'b0}),
    .b({1'b1,open_n86392}),
    .f({\cu_ru/n46 [0],open_n86412}),
    .fco(\cu_ru/sub0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/sub0/u0|cu_ru/sub0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \cu_ru/sub0/u2|cu_ru/sub0/u1  (
    .a(id_rs1_index[2:1]),
    .b(2'b00),
    .fci(\cu_ru/sub0/c1 ),
    .f(\cu_ru/n46 [2:1]),
    .fco(\cu_ru/sub0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/sub0/u0|cu_ru/sub0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \cu_ru/sub0/u4|cu_ru/sub0/u3  (
    .a(id_rs1_index[4:3]),
    .b(2'b00),
    .fci(\cu_ru/sub0/c3 ),
    .f(\cu_ru/n46 [4:3]));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/sub1/u0|cu_ru/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \cu_ru/sub1/u0|cu_ru/sub1/ucin  (
    .a({id_rs2_index[0],1'b0}),
    .b({1'b1,open_n86462}),
    .f({\cu_ru/n49 [0],open_n86482}),
    .fco(\cu_ru/sub1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/sub1/u0|cu_ru/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \cu_ru/sub1/u2|cu_ru/sub1/u1  (
    .a(id_rs2_index[2:1]),
    .b(2'b00),
    .fci(\cu_ru/sub1/c1 ),
    .f(\cu_ru/n49 [2:1]),
    .fco(\cu_ru/sub1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/sub1/u0|cu_ru/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \cu_ru/sub1/u4|cu_ru/sub1/u3  (
    .a(id_rs2_index[4:3]),
    .b(2'b00),
    .fci(\cu_ru/sub1/c3 ),
    .f(\cu_ru/n49 [4:3]));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/sub2/u0|cu_ru/sub2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \cu_ru/sub2/u0|cu_ru/sub2/ucin  (
    .a({wb_rd_index[0],1'b0}),
    .b({1'b1,open_n86532}),
    .f({\cu_ru/n52 [0],open_n86552}),
    .fco(\cu_ru/sub2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/sub2/u0|cu_ru/sub2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \cu_ru/sub2/u2|cu_ru/sub2/u1  (
    .a(wb_rd_index[2:1]),
    .b(2'b00),
    .fci(\cu_ru/sub2/c1 ),
    .f(\cu_ru/n52 [2:1]),
    .fco(\cu_ru/sub2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("cu_ru/sub2/u0|cu_ru/sub2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \cu_ru/sub2/u4|cu_ru/sub2/u3  (
    .a(wb_rd_index[4:3]),
    .b(2'b00),
    .fci(\cu_ru/sub2/c3 ),
    .f(\cu_ru/n52 [4:3]));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u11_al_u9806  (
    .a({ds1[13],ds1[11]}),
    .b({ds1[14],ds1[12]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [13],\exu/alu_au/n17 [11]}),
    .e({\exu/alu_au/n17 [14],\exu/alu_au/n17 [12]}),
    .fci(\exu/alu_au/add0/c11 ),
    .f({\exu/alu_au/add_64 [13],\exu/alu_au/add_64 [11]}),
    .fco(\exu/alu_au/add0/c15 ),
    .fx({\exu/alu_au/add_64 [14],\exu/alu_au/add_64 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u15_al_u9807  (
    .a({ds1[17],ds1[15]}),
    .b({ds1[18],ds1[16]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [17],\exu/alu_au/n17 [15]}),
    .e({\exu/alu_au/n17 [18],\exu/alu_au/n17 [16]}),
    .fci(\exu/alu_au/add0/c15 ),
    .f({\exu/alu_au/add_64 [17],\exu/alu_au/add_64 [15]}),
    .fco(\exu/alu_au/add0/c19 ),
    .fx({\exu/alu_au/add_64 [18],\exu/alu_au/add_64 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u19_al_u9808  (
    .a({ds1[21],ds1[19]}),
    .b({ds1[22],ds1[20]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [21],\exu/alu_au/n17 [19]}),
    .e({\exu/alu_au/n17 [22],\exu/alu_au/n17 [20]}),
    .fci(\exu/alu_au/add0/c19 ),
    .f({\exu/alu_au/add_64 [21],\exu/alu_au/add_64 [19]}),
    .fco(\exu/alu_au/add0/c23 ),
    .fx({\exu/alu_au/add_64 [22],\exu/alu_au/add_64 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u23_al_u9809  (
    .a({ds1[25],ds1[23]}),
    .b({ds1[26],ds1[24]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [25],\exu/alu_au/n17 [23]}),
    .e({\exu/alu_au/n17 [26],\exu/alu_au/n17 [24]}),
    .fci(\exu/alu_au/add0/c23 ),
    .f({\exu/alu_au/add_64 [25],\exu/alu_au/add_64 [23]}),
    .fco(\exu/alu_au/add0/c27 ),
    .fx({\exu/alu_au/add_64 [26],\exu/alu_au/add_64 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u27_al_u9810  (
    .a({ds1[29],ds1[27]}),
    .b({ds1[30],ds1[28]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [29],\exu/alu_au/n17 [27]}),
    .e({\exu/alu_au/n17 [30],\exu/alu_au/n17 [28]}),
    .fci(\exu/alu_au/add0/c27 ),
    .f({\exu/alu_au/add_64 [29],\exu/alu_au/add_64 [27]}),
    .fco(\exu/alu_au/add0/c31 ),
    .fx({\exu/alu_au/add_64 [30],\exu/alu_au/add_64 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u31_al_u9811  (
    .a({ds1[33],ds1[31]}),
    .b({ds1[34],ds1[32]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [33],\exu/alu_au/n17 [31]}),
    .e({\exu/alu_au/n17 [34],\exu/alu_au/n17 [32]}),
    .fci(\exu/alu_au/add0/c31 ),
    .f({\exu/alu_au/add_64 [33],\exu/alu_au/add_64 [31]}),
    .fco(\exu/alu_au/add0/c35 ),
    .fx({\exu/alu_au/add_64 [34],\exu/alu_au/add_64 [32]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u35_al_u9812  (
    .a({ds1[37],ds1[35]}),
    .b({ds1[38],ds1[36]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [37],\exu/alu_au/n17 [35]}),
    .e({\exu/alu_au/n17 [38],\exu/alu_au/n17 [36]}),
    .fci(\exu/alu_au/add0/c35 ),
    .f({\exu/alu_au/add_64 [37],\exu/alu_au/add_64 [35]}),
    .fco(\exu/alu_au/add0/c39 ),
    .fx({\exu/alu_au/add_64 [38],\exu/alu_au/add_64 [36]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u39_al_u9813  (
    .a({ds1[41],ds1[39]}),
    .b({ds1[42],ds1[40]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [41],\exu/alu_au/n17 [39]}),
    .e({\exu/alu_au/n17 [42],\exu/alu_au/n17 [40]}),
    .fci(\exu/alu_au/add0/c39 ),
    .f({\exu/alu_au/add_64 [41],\exu/alu_au/add_64 [39]}),
    .fco(\exu/alu_au/add0/c43 ),
    .fx({\exu/alu_au/add_64 [42],\exu/alu_au/add_64 [40]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u3_al_u9804  (
    .a({ds1[5],ds1[3]}),
    .b({ds1[6],ds1[4]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [5],\exu/alu_au/n17 [3]}),
    .e({\exu/alu_au/n17 [6],\exu/alu_au/n17 [4]}),
    .fci(\exu/alu_au/add0/c3 ),
    .f({\exu/alu_au/add_64 [5],\exu/alu_au/add_64 [3]}),
    .fco(\exu/alu_au/add0/c7 ),
    .fx({\exu/alu_au/add_64 [6],\exu/alu_au/add_64 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u43_al_u9814  (
    .a({ds1[45],ds1[43]}),
    .b({ds1[46],ds1[44]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [45],\exu/alu_au/n17 [43]}),
    .e({\exu/alu_au/n17 [46],\exu/alu_au/n17 [44]}),
    .fci(\exu/alu_au/add0/c43 ),
    .f({\exu/alu_au/add_64 [45],\exu/alu_au/add_64 [43]}),
    .fco(\exu/alu_au/add0/c47 ),
    .fx({\exu/alu_au/add_64 [46],\exu/alu_au/add_64 [44]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u47_al_u9815  (
    .a({ds1[49],ds1[47]}),
    .b({ds1[50],ds1[48]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [49],\exu/alu_au/n17 [47]}),
    .e({\exu/alu_au/n17 [50],\exu/alu_au/n17 [48]}),
    .fci(\exu/alu_au/add0/c47 ),
    .f({\exu/alu_au/add_64 [49],\exu/alu_au/add_64 [47]}),
    .fco(\exu/alu_au/add0/c51 ),
    .fx({\exu/alu_au/add_64 [50],\exu/alu_au/add_64 [48]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u51_al_u9816  (
    .a({ds1[53],ds1[51]}),
    .b({ds1[54],ds1[52]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [53],\exu/alu_au/n17 [51]}),
    .e({\exu/alu_au/n17 [54],\exu/alu_au/n17 [52]}),
    .fci(\exu/alu_au/add0/c51 ),
    .f({\exu/alu_au/add_64 [53],\exu/alu_au/add_64 [51]}),
    .fco(\exu/alu_au/add0/c55 ),
    .fx({\exu/alu_au/add_64 [54],\exu/alu_au/add_64 [52]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u55_al_u9817  (
    .a({ds1[57],ds1[55]}),
    .b({ds1[58],ds1[56]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [57],\exu/alu_au/n17 [55]}),
    .e({\exu/alu_au/n17 [58],\exu/alu_au/n17 [56]}),
    .fci(\exu/alu_au/add0/c55 ),
    .f({\exu/alu_au/add_64 [57],\exu/alu_au/add_64 [55]}),
    .fco(\exu/alu_au/add0/c59 ),
    .fx({\exu/alu_au/add_64 [58],\exu/alu_au/add_64 [56]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u59_al_u9818  (
    .a({ds1[61],ds1[59]}),
    .b({ds1[62],ds1[60]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [61],\exu/alu_au/n17 [59]}),
    .e({\exu/alu_au/n17 [62],\exu/alu_au/n17 [60]}),
    .fci(\exu/alu_au/add0/c59 ),
    .f({\exu/alu_au/add_64 [61],\exu/alu_au/add_64 [59]}),
    .fco(\exu/alu_au/add0/c63 ),
    .fx({\exu/alu_au/add_64 [62],\exu/alu_au/add_64 [60]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y8Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u63_al_u9819  (
    .a({open_n86854,ds1[63]}),
    .c(2'b00),
    .d({open_n86859,\exu/alu_au/n17 [63]}),
    .fci(\exu/alu_au/add0/c63 ),
    .f({open_n86876,\exu/alu_au/add_64 [63]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/u7_al_u9805  (
    .a({ds1[9],ds1[7]}),
    .b({ds1[10],ds1[8]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [9],\exu/alu_au/n17 [7]}),
    .e({\exu/alu_au/n17 [10],\exu/alu_au/n17 [8]}),
    .fci(\exu/alu_au/add0/c7 ),
    .f({\exu/alu_au/add_64 [9],\exu/alu_au/add_64 [7]}),
    .fco(\exu/alu_au/add0/c11 ),
    .fx({\exu/alu_au/add_64 [10],\exu/alu_au/add_64 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add0/ucin_al_u9803"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add0/ucin_al_u9803  (
    .a({ds1[1],1'b0}),
    .b({ds1[2],ds1[0]}),
    .c(2'b00),
    .d({\exu/alu_au/n17 [1],1'b1}),
    .e({\exu/alu_au/n17 [2],\exu/alu_au/n17 [0]}),
    .f({\exu/alu_au/add_64 [1],open_n86917}),
    .fco(\exu/alu_au/add0/c3 ),
    .fx({\exu/alu_au/add_64 [2],\exu/alu_au/add_64 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u0|exu/alu_au/add1/ucin  (
    .a({\exu/alu_au/add_64 [0],1'b0}),
    .b({1'b1,open_n86920}),
    .f({\exu/alu_au/sub_64 [0],open_n86940}),
    .fco(\exu/alu_au/add1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u10|exu/alu_au/add1/u9  (
    .a(\exu/alu_au/add_64 [10:9]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c9 ),
    .f(\exu/alu_au/sub_64 [10:9]),
    .fco(\exu/alu_au/add1/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u12|exu/alu_au/add1/u11  (
    .a(\exu/alu_au/add_64 [12:11]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c11 ),
    .f(\exu/alu_au/sub_64 [12:11]),
    .fco(\exu/alu_au/add1/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u14|exu/alu_au/add1/u13  (
    .a(\exu/alu_au/add_64 [14:13]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c13 ),
    .f(\exu/alu_au/sub_64 [14:13]),
    .fco(\exu/alu_au/add1/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u16|exu/alu_au/add1/u15  (
    .a(\exu/alu_au/add_64 [16:15]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c15 ),
    .f(\exu/alu_au/sub_64 [16:15]),
    .fco(\exu/alu_au/add1/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u18|exu/alu_au/add1/u17  (
    .a(\exu/alu_au/add_64 [18:17]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c17 ),
    .f(\exu/alu_au/sub_64 [18:17]),
    .fco(\exu/alu_au/add1/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u20|exu/alu_au/add1/u19  (
    .a(\exu/alu_au/add_64 [20:19]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c19 ),
    .f(\exu/alu_au/sub_64 [20:19]),
    .fco(\exu/alu_au/add1/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u22|exu/alu_au/add1/u21  (
    .a(\exu/alu_au/add_64 [22:21]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c21 ),
    .f(\exu/alu_au/sub_64 [22:21]),
    .fco(\exu/alu_au/add1/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u24|exu/alu_au/add1/u23  (
    .a(\exu/alu_au/add_64 [24:23]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c23 ),
    .f(\exu/alu_au/sub_64 [24:23]),
    .fco(\exu/alu_au/add1/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u26|exu/alu_au/add1/u25  (
    .a(\exu/alu_au/add_64 [26:25]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c25 ),
    .f(\exu/alu_au/sub_64 [26:25]),
    .fco(\exu/alu_au/add1/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u28|exu/alu_au/add1/u27  (
    .a(\exu/alu_au/add_64 [28:27]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c27 ),
    .f(\exu/alu_au/sub_64 [28:27]),
    .fco(\exu/alu_au/add1/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u2|exu/alu_au/add1/u1  (
    .a(\exu/alu_au/add_64 [2:1]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c1 ),
    .f(\exu/alu_au/sub_64 [2:1]),
    .fco(\exu/alu_au/add1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u30|exu/alu_au/add1/u29  (
    .a(\exu/alu_au/add_64 [30:29]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c29 ),
    .f(\exu/alu_au/sub_64 [30:29]),
    .fco(\exu/alu_au/add1/c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u31_al_u9853  (
    .a({open_n87209,\exu/alu_au/add_64 [31]}),
    .b({open_n87210,1'b0}),
    .fci(\exu/alu_au/add1/c31 ),
    .f({open_n87229,\exu/alu_au/sub_64 [31]}));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u4|exu/alu_au/add1/u3  (
    .a(\exu/alu_au/add_64 [4:3]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c3 ),
    .f(\exu/alu_au/sub_64 [4:3]),
    .fco(\exu/alu_au/add1/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u6|exu/alu_au/add1/u5  (
    .a(\exu/alu_au/add_64 [6:5]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c5 ),
    .f(\exu/alu_au/sub_64 [6:5]),
    .fco(\exu/alu_au/add1/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/add1/u0|exu/alu_au/add1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \exu/alu_au/add1/u8|exu/alu_au/add1/u7  (
    .a(\exu/alu_au/add_64 [8:7]),
    .b(2'b00),
    .fci(\exu/alu_au/add1/c7 ),
    .f(\exu/alu_au/sub_64 [8:7]),
    .fco(\exu/alu_au/add1/c9 ));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u11_al_u9823  (
    .a({as1[13],as1[11]}),
    .b({as1[14],as1[12]}),
    .c(2'b00),
    .d({as2[13],as2[11]}),
    .e({as2[14],as2[12]}),
    .fci(\exu/alu_au/add2/c11 ),
    .f({addr_ex[13],addr_ex[11]}),
    .fco(\exu/alu_au/add2/c15 ),
    .fx({addr_ex[14],addr_ex[12]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u15_al_u9824  (
    .a({as1[17],as1[15]}),
    .b({as1[18],as1[16]}),
    .c(2'b00),
    .d({as2[17],as2[15]}),
    .e({as2[18],as2[16]}),
    .fci(\exu/alu_au/add2/c15 ),
    .f({addr_ex[17],addr_ex[15]}),
    .fco(\exu/alu_au/add2/c19 ),
    .fx({addr_ex[18],addr_ex[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u19_al_u9825  (
    .a({as1[21],as1[19]}),
    .b({as1[22],as1[20]}),
    .c(2'b00),
    .d(as2[20:19]),
    .e({as2[20],as2[20]}),
    .fci(\exu/alu_au/add2/c19 ),
    .f({addr_ex[21],addr_ex[19]}),
    .fco(\exu/alu_au/add2/c23 ),
    .fx({addr_ex[22],addr_ex[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u23_al_u9826  (
    .a({as1[25],as1[23]}),
    .b({as1[26],as1[24]}),
    .c(2'b00),
    .d({as2[20],as2[20]}),
    .e({as2[20],as2[20]}),
    .fci(\exu/alu_au/add2/c23 ),
    .f({addr_ex[25],addr_ex[23]}),
    .fco(\exu/alu_au/add2/c27 ),
    .fx({addr_ex[26],addr_ex[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u27_al_u9827  (
    .a({as1[29],as1[27]}),
    .b({as1[30],as1[28]}),
    .c(2'b00),
    .d({as2[20],as2[20]}),
    .e({as2[20],as2[20]}),
    .fci(\exu/alu_au/add2/c27 ),
    .f({addr_ex[29],addr_ex[27]}),
    .fco(\exu/alu_au/add2/c31 ),
    .fx({addr_ex[30],addr_ex[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u31_al_u9828  (
    .a({as1[33],as1[31]}),
    .b({as1[34],as1[32]}),
    .c(2'b00),
    .d({as2[20],as2[20]}),
    .e({as2[20],as2[20]}),
    .fci(\exu/alu_au/add2/c31 ),
    .f({addr_ex[33],addr_ex[31]}),
    .fco(\exu/alu_au/add2/c35 ),
    .fx({addr_ex[34],addr_ex[32]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u35_al_u9829  (
    .a({as1[37],as1[35]}),
    .b({as1[38],as1[36]}),
    .c(2'b00),
    .d({as2[20],as2[20]}),
    .e({as2[20],as2[20]}),
    .fci(\exu/alu_au/add2/c35 ),
    .f({addr_ex[37],addr_ex[35]}),
    .fco(\exu/alu_au/add2/c39 ),
    .fx({addr_ex[38],addr_ex[36]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u39_al_u9830  (
    .a({as1[41],as1[39]}),
    .b({as1[42],as1[40]}),
    .c(2'b00),
    .d({as2[20],as2[20]}),
    .e({as2[20],as2[20]}),
    .fci(\exu/alu_au/add2/c39 ),
    .f({addr_ex[41],addr_ex[39]}),
    .fco(\exu/alu_au/add2/c43 ),
    .fx({addr_ex[42],addr_ex[40]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u3_al_u9821  (
    .a({as1[5],as1[3]}),
    .b({as1[6],as1[4]}),
    .c(2'b00),
    .d({as2[5],as2[3]}),
    .e({as2[6],as2[4]}),
    .fci(\exu/alu_au/add2/c3 ),
    .f({addr_ex[5],addr_ex[3]}),
    .fco(\exu/alu_au/add2/c7 ),
    .fx({addr_ex[6],addr_ex[4]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u43_al_u9831  (
    .a({as1[45],as1[43]}),
    .b({as1[46],as1[44]}),
    .c(2'b00),
    .d({as2[20],as2[20]}),
    .e({as2[20],as2[20]}),
    .fci(\exu/alu_au/add2/c43 ),
    .f({addr_ex[45],addr_ex[43]}),
    .fco(\exu/alu_au/add2/c47 ),
    .fx({addr_ex[46],addr_ex[44]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u47_al_u9832  (
    .a({as1[49],as1[47]}),
    .b({as1[50],as1[48]}),
    .c(2'b00),
    .d({as2[20],as2[20]}),
    .e({as2[20],as2[20]}),
    .fci(\exu/alu_au/add2/c47 ),
    .f({addr_ex[49],addr_ex[47]}),
    .fco(\exu/alu_au/add2/c51 ),
    .fx({addr_ex[50],addr_ex[48]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u51_al_u9833  (
    .a({as1[53],as1[51]}),
    .b({as1[54],as1[52]}),
    .c(2'b00),
    .d({as2[20],as2[20]}),
    .e({as2[20],as2[20]}),
    .fci(\exu/alu_au/add2/c51 ),
    .f({addr_ex[53],addr_ex[51]}),
    .fco(\exu/alu_au/add2/c55 ),
    .fx({addr_ex[54],addr_ex[52]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u55_al_u9834  (
    .a({as1[57],as1[55]}),
    .b({as1[58],as1[56]}),
    .c(2'b00),
    .d({as2[56],as2[20]}),
    .e({as2[56],as2[56]}),
    .fci(\exu/alu_au/add2/c55 ),
    .f({addr_ex[57],addr_ex[55]}),
    .fco(\exu/alu_au/add2/c59 ),
    .fx({addr_ex[58],addr_ex[56]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u59_al_u9835  (
    .a({as1[61],as1[59]}),
    .b({as1[62],as1[60]}),
    .c(2'b00),
    .d({as2[56],as2[56]}),
    .e({as2[56],as2[56]}),
    .fci(\exu/alu_au/add2/c59 ),
    .f({addr_ex[61],addr_ex[59]}),
    .fco(\exu/alu_au/add2/c63 ),
    .fx({addr_ex[62],addr_ex[60]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y8Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u63_al_u9836  (
    .a({open_n87553,as1[63]}),
    .c(2'b00),
    .d({open_n87558,as2[56]}),
    .fci(\exu/alu_au/add2/c63 ),
    .f({open_n87575,addr_ex[63]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \exu/alu_au/add2/u7_al_u9822  (
    .a({as1[9],as1[7]}),
    .b({as1[10],as1[8]}),
    .c(2'b00),
    .d({as2[9],as2[7]}),
    .e({as2[10],as2[8]}),
    .fci(\exu/alu_au/add2/c7 ),
    .f({addr_ex[9],addr_ex[7]}),
    .fco(\exu/alu_au/add2/c11 ),
    .fx({addr_ex[10],addr_ex[8]}));
  EG_PHY_LSLICE #(
    //.MACRO("exu/alu_au/add2/ucin_al_u9820"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/alu_au/add2/ucin_al_u9820  (
    .a({as1[1],1'b0}),
    .b({as1[2],as1[0]}),
    .c(2'b00),
    .clk(clk_pad),
    .d({as2[1],1'b1}),
    .e({as2[2],as2[0]}),
    .mi({open_n87601,addr_ex[2]}),
    .sr(rst_pad),
    .f({addr_ex[1],open_n87613}),
    .fco(\exu/alu_au/add2/c3 ),
    .fx({addr_ex[2],addr_ex[0]}),
    .q({open_n87614,new_pc[2]}));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_0|exu/alu_au/lt0_cin  (
    .a({ds1[0],1'b0}),
    .b({ds2[0],open_n87615}),
    .fco(\exu/alu_au/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_10|exu/alu_au/lt0_9  (
    .a(ds1[10:9]),
    .b(ds2[10:9]),
    .fci(\exu/alu_au/lt0_c9 ),
    .fco(\exu/alu_au/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_12|exu/alu_au/lt0_11  (
    .a(ds1[12:11]),
    .b(ds2[12:11]),
    .fci(\exu/alu_au/lt0_c11 ),
    .fco(\exu/alu_au/lt0_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_14|exu/alu_au/lt0_13  (
    .a(ds1[14:13]),
    .b(ds2[14:13]),
    .fci(\exu/alu_au/lt0_c13 ),
    .fco(\exu/alu_au/lt0_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_16|exu/alu_au/lt0_15  (
    .a(ds1[16:15]),
    .b(ds2[16:15]),
    .fci(\exu/alu_au/lt0_c15 ),
    .fco(\exu/alu_au/lt0_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_18|exu/alu_au/lt0_17  (
    .a(ds1[18:17]),
    .b(ds2[18:17]),
    .fci(\exu/alu_au/lt0_c17 ),
    .fco(\exu/alu_au/lt0_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_20|exu/alu_au/lt0_19  (
    .a(ds1[20:19]),
    .b(ds2[20:19]),
    .fci(\exu/alu_au/lt0_c19 ),
    .fco(\exu/alu_au/lt0_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_22|exu/alu_au/lt0_21  (
    .a(ds1[22:21]),
    .b(ds2[22:21]),
    .fci(\exu/alu_au/lt0_c21 ),
    .fco(\exu/alu_au/lt0_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_24|exu/alu_au/lt0_23  (
    .a(ds1[24:23]),
    .b(ds2[24:23]),
    .fci(\exu/alu_au/lt0_c23 ),
    .fco(\exu/alu_au/lt0_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_26|exu/alu_au/lt0_25  (
    .a(ds1[26:25]),
    .b(ds2[26:25]),
    .fci(\exu/alu_au/lt0_c25 ),
    .fco(\exu/alu_au/lt0_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_28|exu/alu_au/lt0_27  (
    .a(ds1[28:27]),
    .b(ds2[28:27]),
    .fci(\exu/alu_au/lt0_c27 ),
    .fco(\exu/alu_au/lt0_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_2|exu/alu_au/lt0_1  (
    .a(ds1[2:1]),
    .b(ds2[2:1]),
    .fci(\exu/alu_au/lt0_c1 ),
    .fco(\exu/alu_au/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_30|exu/alu_au/lt0_29  (
    .a(ds1[30:29]),
    .b(ds2[30:29]),
    .fci(\exu/alu_au/lt0_c29 ),
    .fco(\exu/alu_au/lt0_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_32|exu/alu_au/lt0_31  (
    .a(ds1[32:31]),
    .b(ds2[32:31]),
    .fci(\exu/alu_au/lt0_c31 ),
    .fco(\exu/alu_au/lt0_c33 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y8Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_34|exu/alu_au/lt0_33  (
    .a(ds1[34:33]),
    .b(ds2[34:33]),
    .fci(\exu/alu_au/lt0_c33 ),
    .fco(\exu/alu_au/lt0_c35 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y9Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_36|exu/alu_au/lt0_35  (
    .a(ds1[36:35]),
    .b(ds2[36:35]),
    .fci(\exu/alu_au/lt0_c35 ),
    .fco(\exu/alu_au/lt0_c37 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y9Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_38|exu/alu_au/lt0_37  (
    .a(ds1[38:37]),
    .b(ds2[38:37]),
    .fci(\exu/alu_au/lt0_c37 ),
    .fco(\exu/alu_au/lt0_c39 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y10Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_40|exu/alu_au/lt0_39  (
    .a(ds1[40:39]),
    .b(ds2[40:39]),
    .fci(\exu/alu_au/lt0_c39 ),
    .fco(\exu/alu_au/lt0_c41 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y10Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_42|exu/alu_au/lt0_41  (
    .a(ds1[42:41]),
    .b(ds2[42:41]),
    .fci(\exu/alu_au/lt0_c41 ),
    .fco(\exu/alu_au/lt0_c43 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y11Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_44|exu/alu_au/lt0_43  (
    .a(ds1[44:43]),
    .b(ds2[44:43]),
    .fci(\exu/alu_au/lt0_c43 ),
    .fco(\exu/alu_au/lt0_c45 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y11Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_46|exu/alu_au/lt0_45  (
    .a(ds1[46:45]),
    .b(ds2[46:45]),
    .fci(\exu/alu_au/lt0_c45 ),
    .fco(\exu/alu_au/lt0_c47 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y12Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_48|exu/alu_au/lt0_47  (
    .a(ds1[48:47]),
    .b(ds2[48:47]),
    .fci(\exu/alu_au/lt0_c47 ),
    .fco(\exu/alu_au/lt0_c49 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_4|exu/alu_au/lt0_3  (
    .a(ds1[4:3]),
    .b(ds2[4:3]),
    .fci(\exu/alu_au/lt0_c3 ),
    .fco(\exu/alu_au/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y12Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_50|exu/alu_au/lt0_49  (
    .a(ds1[50:49]),
    .b(ds2[50:49]),
    .fci(\exu/alu_au/lt0_c49 ),
    .fco(\exu/alu_au/lt0_c51 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y13Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_52|exu/alu_au/lt0_51  (
    .a(ds1[52:51]),
    .b(ds2[52:51]),
    .fci(\exu/alu_au/lt0_c51 ),
    .fco(\exu/alu_au/lt0_c53 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y13Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_54|exu/alu_au/lt0_53  (
    .a(ds1[54:53]),
    .b(ds2[54:53]),
    .fci(\exu/alu_au/lt0_c53 ),
    .fco(\exu/alu_au/lt0_c55 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y14Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_56|exu/alu_au/lt0_55  (
    .a(ds1[56:55]),
    .b(ds2[56:55]),
    .fci(\exu/alu_au/lt0_c55 ),
    .fco(\exu/alu_au/lt0_c57 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y14Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_58|exu/alu_au/lt0_57  (
    .a(ds1[58:57]),
    .b(ds2[58:57]),
    .fci(\exu/alu_au/lt0_c57 ),
    .fco(\exu/alu_au/lt0_c59 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y15Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_60|exu/alu_au/lt0_59  (
    .a(ds1[60:59]),
    .b(ds2[60:59]),
    .fci(\exu/alu_au/lt0_c59 ),
    .fco(\exu/alu_au/lt0_c61 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y15Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_62|exu/alu_au/lt0_61  (
    .a(ds1[62:61]),
    .b(ds2[62:61]),
    .fci(\exu/alu_au/lt0_c61 ),
    .fco(\exu/alu_au/lt0_c63 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_6|exu/alu_au/lt0_5  (
    .a(ds1[6:5]),
    .b(ds2[6:5]),
    .fci(\exu/alu_au/lt0_c5 ),
    .fco(\exu/alu_au/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_8|exu/alu_au/lt0_7  (
    .a(ds1[8:7]),
    .b(ds2[8:7]),
    .fci(\exu/alu_au/lt0_c7 ),
    .fco(\exu/alu_au/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt0_0|exu/alu_au/lt0_cin"),
    //.R_POSITION("X0Y16Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt0_cout|exu/alu_au/lt0_63  (
    .a({1'b0,ds1[63]}),
    .b({1'b1,ds2[63]}),
    .fci(\exu/alu_au/lt0_c63 ),
    .f({\exu/alu_au/n5 ,open_n88403}));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_0|exu/alu_au/lt1_cin  (
    .a({ds2[0],1'b0}),
    .b({ds1[0],open_n88409}),
    .fco(\exu/alu_au/lt1_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_10|exu/alu_au/lt1_9  (
    .a(ds2[10:9]),
    .b(ds1[10:9]),
    .fci(\exu/alu_au/lt1_c9 ),
    .fco(\exu/alu_au/lt1_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_12|exu/alu_au/lt1_11  (
    .a(ds2[12:11]),
    .b(ds1[12:11]),
    .fci(\exu/alu_au/lt1_c11 ),
    .fco(\exu/alu_au/lt1_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_14|exu/alu_au/lt1_13  (
    .a(ds2[14:13]),
    .b(ds1[14:13]),
    .fci(\exu/alu_au/lt1_c13 ),
    .fco(\exu/alu_au/lt1_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_16|exu/alu_au/lt1_15  (
    .a(ds2[16:15]),
    .b(ds1[16:15]),
    .fci(\exu/alu_au/lt1_c15 ),
    .fco(\exu/alu_au/lt1_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_18|exu/alu_au/lt1_17  (
    .a(ds2[18:17]),
    .b(ds1[18:17]),
    .fci(\exu/alu_au/lt1_c17 ),
    .fco(\exu/alu_au/lt1_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_20|exu/alu_au/lt1_19  (
    .a(ds2[20:19]),
    .b(ds1[20:19]),
    .fci(\exu/alu_au/lt1_c19 ),
    .fco(\exu/alu_au/lt1_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_22|exu/alu_au/lt1_21  (
    .a(ds2[22:21]),
    .b(ds1[22:21]),
    .fci(\exu/alu_au/lt1_c21 ),
    .fco(\exu/alu_au/lt1_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_24|exu/alu_au/lt1_23  (
    .a(ds2[24:23]),
    .b(ds1[24:23]),
    .fci(\exu/alu_au/lt1_c23 ),
    .fco(\exu/alu_au/lt1_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_26|exu/alu_au/lt1_25  (
    .a(ds2[26:25]),
    .b(ds1[26:25]),
    .fci(\exu/alu_au/lt1_c25 ),
    .fco(\exu/alu_au/lt1_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_28|exu/alu_au/lt1_27  (
    .a(ds2[28:27]),
    .b(ds1[28:27]),
    .fci(\exu/alu_au/lt1_c27 ),
    .fco(\exu/alu_au/lt1_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_2|exu/alu_au/lt1_1  (
    .a(ds2[2:1]),
    .b(ds1[2:1]),
    .fci(\exu/alu_au/lt1_c1 ),
    .fco(\exu/alu_au/lt1_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_30|exu/alu_au/lt1_29  (
    .a(ds2[30:29]),
    .b(ds1[30:29]),
    .fci(\exu/alu_au/lt1_c29 ),
    .fco(\exu/alu_au/lt1_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_32|exu/alu_au/lt1_31  (
    .a(ds2[32:31]),
    .b(ds1[32:31]),
    .fci(\exu/alu_au/lt1_c31 ),
    .fco(\exu/alu_au/lt1_c33 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y8Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_34|exu/alu_au/lt1_33  (
    .a(ds2[34:33]),
    .b(ds1[34:33]),
    .fci(\exu/alu_au/lt1_c33 ),
    .fco(\exu/alu_au/lt1_c35 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y9Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_36|exu/alu_au/lt1_35  (
    .a(ds2[36:35]),
    .b(ds1[36:35]),
    .fci(\exu/alu_au/lt1_c35 ),
    .fco(\exu/alu_au/lt1_c37 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y9Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_38|exu/alu_au/lt1_37  (
    .a(ds2[38:37]),
    .b(ds1[38:37]),
    .fci(\exu/alu_au/lt1_c37 ),
    .fco(\exu/alu_au/lt1_c39 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y10Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_40|exu/alu_au/lt1_39  (
    .a(ds2[40:39]),
    .b(ds1[40:39]),
    .fci(\exu/alu_au/lt1_c39 ),
    .fco(\exu/alu_au/lt1_c41 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y10Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_42|exu/alu_au/lt1_41  (
    .a(ds2[42:41]),
    .b(ds1[42:41]),
    .fci(\exu/alu_au/lt1_c41 ),
    .fco(\exu/alu_au/lt1_c43 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y11Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_44|exu/alu_au/lt1_43  (
    .a(ds2[44:43]),
    .b(ds1[44:43]),
    .fci(\exu/alu_au/lt1_c43 ),
    .fco(\exu/alu_au/lt1_c45 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y11Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_46|exu/alu_au/lt1_45  (
    .a(ds2[46:45]),
    .b(ds1[46:45]),
    .fci(\exu/alu_au/lt1_c45 ),
    .fco(\exu/alu_au/lt1_c47 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y12Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_48|exu/alu_au/lt1_47  (
    .a(ds2[48:47]),
    .b(ds1[48:47]),
    .fci(\exu/alu_au/lt1_c47 ),
    .fco(\exu/alu_au/lt1_c49 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_4|exu/alu_au/lt1_3  (
    .a(ds2[4:3]),
    .b(ds1[4:3]),
    .fci(\exu/alu_au/lt1_c3 ),
    .fco(\exu/alu_au/lt1_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y12Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_50|exu/alu_au/lt1_49  (
    .a(ds2[50:49]),
    .b(ds1[50:49]),
    .fci(\exu/alu_au/lt1_c49 ),
    .fco(\exu/alu_au/lt1_c51 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y13Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_52|exu/alu_au/lt1_51  (
    .a(ds2[52:51]),
    .b(ds1[52:51]),
    .fci(\exu/alu_au/lt1_c51 ),
    .fco(\exu/alu_au/lt1_c53 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y13Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_54|exu/alu_au/lt1_53  (
    .a(ds2[54:53]),
    .b(ds1[54:53]),
    .fci(\exu/alu_au/lt1_c53 ),
    .fco(\exu/alu_au/lt1_c55 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y14Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_56|exu/alu_au/lt1_55  (
    .a(ds2[56:55]),
    .b(ds1[56:55]),
    .fci(\exu/alu_au/lt1_c55 ),
    .fco(\exu/alu_au/lt1_c57 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y14Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_58|exu/alu_au/lt1_57  (
    .a(ds2[58:57]),
    .b(ds1[58:57]),
    .fci(\exu/alu_au/lt1_c57 ),
    .fco(\exu/alu_au/lt1_c59 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y15Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_60|exu/alu_au/lt1_59  (
    .a(ds2[60:59]),
    .b(ds1[60:59]),
    .fci(\exu/alu_au/lt1_c59 ),
    .fco(\exu/alu_au/lt1_c61 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y15Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_62|exu/alu_au/lt1_61  (
    .a(ds2[62:61]),
    .b(ds1[62:61]),
    .fci(\exu/alu_au/lt1_c61 ),
    .fco(\exu/alu_au/lt1_c63 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_6|exu/alu_au/lt1_5  (
    .a(ds2[6:5]),
    .b(ds1[6:5]),
    .fci(\exu/alu_au/lt1_c5 ),
    .fco(\exu/alu_au/lt1_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_8|exu/alu_au/lt1_7  (
    .a(ds2[8:7]),
    .b(ds1[8:7]),
    .fci(\exu/alu_au/lt1_c7 ),
    .fco(\exu/alu_au/lt1_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/alu_au/lt1_0|exu/alu_au/lt1_cin"),
    //.R_POSITION("X0Y16Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \exu/alu_au/lt1_cout|exu/alu_au/lt1_63  (
    .a({1'b0,ds2[63]}),
    .b({1'b1,ds1[63]}),
    .fci(\exu/alu_au/lt1_c63 ),
    .f({\exu/alu_au/n12 ,open_n89197}));
  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/ebreak_reg|exu/ecall_reg  (
    .a({ex_ebreak,open_n89203}),
    .b({ex_ecall,open_n89204}),
    .c({ex_jmp,rst_pad}),
    .clk(clk_pad),
    .d({ex_system,ex_nop}),
    .mi({ex_ebreak,ex_ecall}),
    .sr(\exu/n86 ),
    .f({_al_u9192_o,\exu/n86 }),
    .q({wb_ebreak,wb_ecall}));  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/id_jmp_reg|exu/int_acc_reg  (
    .a({open_n89223,_al_u9192_o}),
    .b({wb_system,ex_int_acc}),
    .c({wb_int_acc,1'b0}),
    .clk(clk_pad),
    .d({wb_jmp,1'b0}),
    .mi({ex_jmp,ex_int_acc}),
    .sr(\exu/n86 ),
    .f({_al_u4837_o,_al_u9193_o}),
    .q({wb_jmp,wb_int_acc}));  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/id_system_reg  (
    .clk(clk_pad),
    .mi({open_n89261,ex_system}),
    .sr(\exu/n86 ),
    .q({open_n89267,wb_system}));  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~D))"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/ins_acc_fault_reg|exu/ins_addr_mis_reg  (
    .b({wb_ins_addr_mis,\cu_ru/medeleg [0]}),
    .c({wb_ins_page_fault,wb_ins_addr_mis}),
    .clk(clk_pad),
    .d({wb_ins_acc_fault,priv[3]}),
    .mi({ex_ins_acc_fault,ex_ins_addr_mis}),
    .sr(\exu/n86 ),
    .f({_al_u4133_o,\cu_ru/medeleg_exc_ctrl/iam_target_m_lutinv }),
    .q({wb_ins_acc_fault,wb_ins_addr_mis}));  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*A*~(C*B))"),
    //.LUTF1("~(~C*D)"),
    //.LUTG0("~(~D*A*~(C*B))"),
    //.LUTG1("~(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111010101),
    .INIT_LUTF1(16'b1111000011111111),
    .INIT_LUTG0(16'b1111111111010101),
    .INIT_LUTG1(16'b1111000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/ld_page_fault_reg|exu/st_page_fault_reg  (
    .a({open_n89284,_al_u6724_o}),
    .b({open_n89285,_al_u2910_o}),
    .c({_al_u6725_o,_al_u6725_o}),
    .clk(clk_pad),
    .d({_al_u6724_o,_al_u7195_o}),
    .sr(\exu/n86 ),
    .q({wb_ld_page_fault,wb_st_page_fault}));  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTF1("~(~C*B*~D)"),
    //.LUTG0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG1("~(~C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110011),
    .INIT_LUTF1(16'b1111111111110011),
    .INIT_LUTG0(16'b1111000000110011),
    .INIT_LUTG1(16'b1111111111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg2_b43|cu_ru/m_cycle_event/reg1_b43  (
    .b({_al_u3634_o,_al_u3304_o}),
    .c({\exu/alu_au/n55 [43],data_csr[43]}),
    .clk(clk_pad),
    .d({\exu/alu_au/n53 [43],_al_u3253_o}),
    .sr(rst_pad),
    .f({\exu/alu_data_mem_csr [43],open_n89327}),
    .q({data_csr[43],\cu_ru/mcycle [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUT1("~(~C*B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000110011),
    .INIT_LUT1(16'b1111111111110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg2_b63|cu_ru/m_cycle_event/reg1_b63  (
    .b({_al_u3460_o,_al_u3260_o}),
    .c({\exu/alu_au/n55 [63],data_csr[63]}),
    .clk(clk_pad),
    .d({\exu/alu_au/n53 [63],_al_u3253_o}),
    .sr(rst_pad),
    .f({\exu/alu_data_mem_csr [63],open_n89346}),
    .q({data_csr[63],\cu_ru/mcycle [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b12|exu/reg5_b12  (
    .b({\biu/cache_ctrl_logic/l1i_va [12],addr_ex[12]}),
    .c({addr_ex[12],ex_exc_code[12]}),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_value ,ex_more_exception_neg_lutinv}),
    .mi({addr_ex[12],open_n89356}),
    .sr(rst_pad),
    .f({_al_u6389_o,open_n89368}),
    .q({new_pc[12],wb_exc_code[12]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(C@D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b16|exu/reg5_b16  (
    .b({open_n89374,addr_ex[16]}),
    .c({addr_ex[16],ex_exc_code[16]}),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_va [16],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[16],open_n89386}),
    .sr(rst_pad),
    .f({\biu/cache_ctrl_logic/eq1/xor_i0[4]_i1[4]_o_lutinv ,open_n89387}),
    .q({new_pc[16],wb_exc_code[16]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b17|exu/reg5_b17  (
    .a({\biu/cache_ctrl_logic/l1d_va [17],open_n89391}),
    .b({\biu/cache_ctrl_logic/l1d_va [26],addr_ex[17]}),
    .c({addr_ex[17],ex_exc_code[17]}),
    .clk(clk_pad),
    .d({addr_ex[26],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[17],open_n89403}),
    .sr(rst_pad),
    .f({_al_u6304_o,open_n89404}),
    .q({new_pc[17],wb_exc_code[17]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(~C*A))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~(D*~B)*~(~C*A))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100010011110101),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1100010011110101),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b18|exu/reg3_b36  (
    .a({\biu/cache_ctrl_logic/l1d_va [18],\biu/cache_ctrl_logic/l1d_va [18]}),
    .b({\biu/cache_ctrl_logic/l1d_va [24],\biu/cache_ctrl_logic/l1d_va [36]}),
    .c({addr_ex[18],addr_ex[18]}),
    .clk(clk_pad),
    .d({addr_ex[24],addr_ex[36]}),
    .mi({addr_ex[18],addr_ex[36]}),
    .sr(rst_pad),
    .f({_al_u6281_o,_al_u6249_o}),
    .q({new_pc[18],new_pc[36]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b19|exu/reg5_b19  (
    .a({\biu/cache_ctrl_logic/l1d_va [19],open_n89426}),
    .b({\biu/cache_ctrl_logic/l1d_va [29],addr_ex[19]}),
    .c({addr_ex[19],ex_exc_code[19]}),
    .clk(clk_pad),
    .d({addr_ex[29],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[19],open_n89438}),
    .sr(rst_pad),
    .f({_al_u6268_o,open_n89439}),
    .q({new_pc[19],wb_exc_code[19]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b20|exu/reg5_b20  (
    .a({\biu/cache_ctrl_logic/l1d_va [12],open_n89443}),
    .b({\biu/cache_ctrl_logic/l1d_va [20],addr_ex[20]}),
    .c({addr_ex[12],ex_exc_code[20]}),
    .clk(clk_pad),
    .d({addr_ex[20],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[20],open_n89448}),
    .sr(rst_pad),
    .f({_al_u6247_o,open_n89460}),
    .q({new_pc[20],wb_exc_code[20]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b25|exu/reg5_b53  (
    .a({\biu/cache_ctrl_logic/l1d_va [25],open_n89464}),
    .b({\biu/cache_ctrl_logic/l1d_va [53],open_n89465}),
    .c({addr_ex[25],addr_ex[53]}),
    .clk(clk_pad),
    .d({addr_ex[53],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[25],open_n89477}),
    .sr(rst_pad),
    .f({_al_u6293_o,open_n89478}),
    .q({new_pc[25],wb_exc_code[53]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~(C@D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b27|exu/reg5_b27  (
    .b({open_n89484,addr_ex[27]}),
    .c({addr_ex[27],ex_exc_code[27]}),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1d_va [27],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[27],open_n89496}),
    .sr(rst_pad),
    .f({_al_u6272_o,open_n89497}),
    .q({new_pc[27],wb_exc_code[27]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*~B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1100010011110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b28|exu/reg5_b28  (
    .a({\biu/cache_ctrl_logic/l1d_va [28],open_n89501}),
    .b({\biu/cache_ctrl_logic/l1d_va [38],addr_ex[28]}),
    .c({addr_ex[28],ex_exc_code[28]}),
    .clk(clk_pad),
    .d({addr_ex[38],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[28],open_n89513}),
    .sr(rst_pad),
    .f({_al_u6307_o,open_n89514}),
    .q({new_pc[28],wb_exc_code[28]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b30|exu/reg5_b30  (
    .a({\biu/cache_ctrl_logic/l1i_va [30],open_n89518}),
    .b({\biu/cache_ctrl_logic/l1i_va [34],addr_ex[30]}),
    .c({addr_ex[30],ex_exc_code[30]}),
    .clk(clk_pad),
    .d({addr_ex[34],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[30],open_n89523}),
    .sr(rst_pad),
    .f({_al_u6405_o,open_n89535}),
    .q({new_pc[30],wb_exc_code[30]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b32|exu/reg5_b32  (
    .a({\biu/cache_ctrl_logic/l1d_va [32],open_n89539}),
    .b({\biu/cache_ctrl_logic/l1d_va [50],open_n89540}),
    .c({addr_ex[32],addr_ex[32]}),
    .clk(clk_pad),
    .d({addr_ex[50],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[32],open_n89552}),
    .sr(rst_pad),
    .f({_al_u6303_o,open_n89553}),
    .q({new_pc[32],wb_exc_code[32]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b34|exu/reg3_b38  (
    .a({\biu/cache_ctrl_logic/l1d_va [34],\biu/cache_ctrl_logic/l1d_va [34]}),
    .b({\biu/cache_ctrl_logic/l1d_va [42],\biu/cache_ctrl_logic/l1d_va [38]}),
    .c({addr_ex[34],addr_ex[34]}),
    .clk(clk_pad),
    .d({addr_ex[42],addr_ex[38]}),
    .mi({addr_ex[34],addr_ex[38]}),
    .sr(rst_pad),
    .f({_al_u6306_o,_al_u6277_o}),
    .q({new_pc[34],new_pc[38]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b40|exu/reg3_b24  (
    .a({open_n89571,\biu/cache_ctrl_logic/l1d_va [24]}),
    .b({\biu/cache_ctrl_logic/l1d_va [40],\biu/cache_ctrl_logic/l1d_va [36]}),
    .c({addr_ex[40],addr_ex[24]}),
    .clk(clk_pad),
    .d({_al_u6299_o,addr_ex[36]}),
    .mi({addr_ex[40],addr_ex[24]}),
    .sr(rst_pad),
    .f({_al_u6300_o,_al_u6299_o}),
    .q({new_pc[40],new_pc[24]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b41|exu/reg5_b41  (
    .a({\biu/cache_ctrl_logic/l1d_va [41],open_n89586}),
    .b({\biu/cache_ctrl_logic/l1d_va [62],open_n89587}),
    .c({addr_ex[41],addr_ex[41]}),
    .clk(clk_pad),
    .d({addr_ex[62],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[41],open_n89592}),
    .sr(rst_pad),
    .f({_al_u6296_o,open_n89604}),
    .q({new_pc[41],wb_exc_code[41]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(~D*B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1010111100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b42|exu/reg5_b42  (
    .a({\biu/cache_ctrl_logic/l1d_va [42],open_n89608}),
    .b({\biu/cache_ctrl_logic/l1d_va [54],open_n89609}),
    .c({addr_ex[42],addr_ex[42]}),
    .clk(clk_pad),
    .d({addr_ex[54],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[42],open_n89621}),
    .sr(rst_pad),
    .f({_al_u6275_o,open_n89622}),
    .q({new_pc[42],wb_exc_code[42]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b43|exu/reg5_b43  (
    .a({\biu/cache_ctrl_logic/l1d_va [43],open_n89626}),
    .b({\biu/cache_ctrl_logic/l1d_va [45],open_n89627}),
    .c({addr_ex[43],addr_ex[43]}),
    .clk(clk_pad),
    .d({addr_ex[45],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[43],open_n89632}),
    .sr(rst_pad),
    .f({_al_u6287_o,open_n89644}),
    .q({new_pc[43],wb_exc_code[43]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b45|exu/reg5_b45  (
    .a({\biu/cache_ctrl_logic/l1d_va [45],open_n89648}),
    .b({\biu/cache_ctrl_logic/l1d_va [59],open_n89649}),
    .c({addr_ex[45],addr_ex[45]}),
    .clk(clk_pad),
    .d({addr_ex[59],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[45],open_n89661}),
    .sr(rst_pad),
    .f({_al_u6289_o,open_n89662}),
    .q({new_pc[45],wb_exc_code[45]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(~D*B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1010111100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b46|exu/reg5_b46  (
    .a({\biu/cache_ctrl_logic/l1d_va [43],open_n89666}),
    .b({\biu/cache_ctrl_logic/l1d_va [46],open_n89667}),
    .c({addr_ex[43],addr_ex[46]}),
    .clk(clk_pad),
    .d({addr_ex[46],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[46],open_n89679}),
    .sr(rst_pad),
    .f({_al_u6274_o,open_n89680}),
    .q({new_pc[46],wb_exc_code[46]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b48|exu/reg5_b48  (
    .a({\biu/cache_ctrl_logic/l1d_va [30],open_n89684}),
    .b({\biu/cache_ctrl_logic/l1d_va [48],open_n89685}),
    .c({addr_ex[30],addr_ex[48]}),
    .clk(clk_pad),
    .d({addr_ex[48],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[48],open_n89690}),
    .sr(rst_pad),
    .f({_al_u6284_o,open_n89702}),
    .q({new_pc[48],wb_exc_code[48]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b49|exu/reg5_b57  (
    .a({\biu/cache_ctrl_logic/l1d_va [49],open_n89706}),
    .b({\biu/cache_ctrl_logic/l1d_va [57],open_n89707}),
    .c({addr_ex[49],addr_ex[57]}),
    .clk(clk_pad),
    .d({addr_ex[57],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[49],open_n89712}),
    .sr(rst_pad),
    .f({_al_u6264_o,open_n89724}),
    .q({new_pc[49],wb_exc_code[57]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b50|exu/reg5_b50  (
    .a({\biu/cache_ctrl_logic/l1d_va [50],open_n89728}),
    .b({\biu/cache_ctrl_logic/l1d_va [59],open_n89729}),
    .c({addr_ex[50],addr_ex[50]}),
    .clk(clk_pad),
    .d({addr_ex[59],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[50],open_n89734}),
    .sr(rst_pad),
    .f({_al_u6288_o,open_n89746}),
    .q({new_pc[50],wb_exc_code[50]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b51|exu/reg5_b51  (
    .b({\biu/cache_ctrl_logic/l1d_va [51],open_n89752}),
    .c({addr_ex[51],addr_ex[51]}),
    .clk(clk_pad),
    .d({_al_u6243_o,ex_more_exception_neg_lutinv}),
    .mi({addr_ex[51],open_n89757}),
    .sr(rst_pad),
    .f({_al_u6244_o,open_n89769}),
    .q({new_pc[51],wb_exc_code[51]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(~D*B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1010111100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b52|exu/reg5_b52  (
    .a({\biu/cache_ctrl_logic/l1d_va [46],open_n89773}),
    .b({\biu/cache_ctrl_logic/l1d_va [52],open_n89774}),
    .c({addr_ex[46],addr_ex[52]}),
    .clk(clk_pad),
    .d({addr_ex[52],ex_more_exception_neg_lutinv}),
    .mi({addr_ex[52],open_n89786}),
    .sr(rst_pad),
    .f({_al_u6250_o,open_n89787}),
    .q({new_pc[52],wb_exc_code[52]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/EX/exu.v(342)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(~(D*~B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1100010011110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg3_b58|exu/reg3_b54  (
    .a({\biu/cache_ctrl_logic/l1d_va [48],\biu/cache_ctrl_logic/l1d_va [54]}),
    .b({\biu/cache_ctrl_logic/l1d_va [58],\biu/cache_ctrl_logic/l1d_va [58]}),
    .c({addr_ex[48],addr_ex[54]}),
    .clk(clk_pad),
    .d({addr_ex[58],addr_ex[58]}),
    .mi({addr_ex[58],addr_ex[54]}),
    .sr(rst_pad),
    .f({_al_u6283_o,_al_u6286_o}),
    .q({new_pc[58],new_pc[54]}));  // ../../RTL/CPU/EX/exu.v(342)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTF1("(D*~(C)*~((B*~A))+D*C*~((B*~A))+~(D)*C*(B*~A)+D*C*(B*~A))"),
    //.LUTG0("(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTG1("(D*~(C)*~((B*~A))+D*C*~((B*~A))+~(D)*C*(B*~A)+D*C*(B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001111),
    .INIT_LUTF1(16'b1111101101000000),
    .INIT_LUTG0(16'b1100000011001111),
    .INIT_LUTG1(16'b1111101101000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b0|cu_ru/m_s_epc/reg1_b0  (
    .a({_al_u5353_o,open_n89805}),
    .b({pc_jmp,\cu_ru/m_s_epc/n2 [0]}),
    .c({new_pc[0],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({wb_ins_pc[0],_al_u6696_o}),
    .mi({ex_ins_pc[0],open_n89810}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [0],open_n89822}),
    .q({wb_ins_pc[0],\cu_ru/mepc [0]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b10|cu_ru/m_s_epc/reg1_b10  (
    .b({_al_u5599_o,\cu_ru/m_s_epc/n2 [10]}),
    .c({wb_ins_pc[10],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6694_o}),
    .mi({ex_ins_pc[10],open_n89839}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [10],open_n89840}),
    .q({wb_ins_pc[10],\cu_ru/mepc [10]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b11|cu_ru/m_s_epc/reg1_b11  (
    .b({_al_u5595_o,\cu_ru/m_s_epc/n2 [11]}),
    .c({wb_ins_pc[11],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6692_o}),
    .mi({ex_ins_pc[11],open_n89850}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [11],open_n89862}),
    .q({wb_ins_pc[11],\cu_ru/mepc [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b12|cu_ru/m_s_epc/reg1_b12  (
    .b({_al_u5591_o,\cu_ru/m_s_epc/n2 [12]}),
    .c({wb_ins_pc[12],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6690_o}),
    .mi({ex_ins_pc[12],open_n89872}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [12],open_n89884}),
    .q({wb_ins_pc[12],\cu_ru/mepc [12]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b13|cu_ru/m_s_epc/reg1_b13  (
    .b({_al_u5587_o,\cu_ru/m_s_epc/n2 [13]}),
    .c({wb_ins_pc[13],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6688_o}),
    .mi({ex_ins_pc[13],open_n89901}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [13],open_n89902}),
    .q({wb_ins_pc[13],\cu_ru/mepc [13]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b14|cu_ru/m_s_epc/reg1_b14  (
    .b({_al_u5583_o,\cu_ru/m_s_epc/n2 [14]}),
    .c({wb_ins_pc[14],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6686_o}),
    .mi({ex_ins_pc[14],open_n89919}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [14],open_n89920}),
    .q({wb_ins_pc[14],\cu_ru/mepc [14]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b15|cu_ru/m_s_epc/reg1_b15  (
    .b({_al_u5579_o,\cu_ru/m_s_epc/n2 [15]}),
    .c({wb_ins_pc[15],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6684_o}),
    .mi({ex_ins_pc[15],open_n89930}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [15],open_n89942}),
    .q({wb_ins_pc[15],\cu_ru/mepc [15]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b16|cu_ru/m_s_epc/reg1_b16  (
    .b({_al_u5575_o,\cu_ru/m_s_epc/n2 [16]}),
    .c({wb_ins_pc[16],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6682_o}),
    .mi({ex_ins_pc[16],open_n89952}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [16],open_n89964}),
    .q({wb_ins_pc[16],\cu_ru/mepc [16]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b17|cu_ru/m_s_epc/reg1_b17  (
    .b({_al_u5571_o,\cu_ru/m_s_epc/n2 [17]}),
    .c({wb_ins_pc[17],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6680_o}),
    .mi({ex_ins_pc[17],open_n89981}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [17],open_n89982}),
    .q({wb_ins_pc[17],\cu_ru/mepc [17]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b18|cu_ru/m_s_epc/reg1_b18  (
    .b({_al_u5567_o,\cu_ru/m_s_epc/n2 [18]}),
    .c({wb_ins_pc[18],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6678_o}),
    .mi({ex_ins_pc[18],open_n89999}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [18],open_n90000}),
    .q({wb_ins_pc[18],\cu_ru/mepc [18]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b19|cu_ru/m_s_epc/reg1_b19  (
    .b({_al_u5563_o,\cu_ru/m_s_epc/n2 [19]}),
    .c({wb_ins_pc[19],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6676_o}),
    .mi({ex_ins_pc[19],open_n90010}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [19],open_n90022}),
    .q({wb_ins_pc[19],\cu_ru/mepc [19]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(D*~(C)*~((B*~A))+D*C*~((B*~A))+~(D)*C*(B*~A)+D*C*(B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111101101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b1|cu_ru/m_s_epc/reg1_b1  (
    .a({_al_u5353_o,open_n90026}),
    .b({pc_jmp,\cu_ru/m_s_epc/n2 [1]}),
    .c({new_pc[1],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({wb_ins_pc[1],_al_u6674_o}),
    .mi({ex_ins_pc[1],open_n90038}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [1],open_n90039}),
    .q({wb_ins_pc[1],\cu_ru/mepc [1]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b20|cu_ru/m_s_epc/reg1_b20  (
    .b({_al_u5555_o,\cu_ru/m_s_epc/n2 [20]}),
    .c({wb_ins_pc[20],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6672_o}),
    .mi({ex_ins_pc[20],open_n90056}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [20],open_n90057}),
    .q({wb_ins_pc[20],\cu_ru/mepc [20]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b21|cu_ru/m_s_epc/reg1_b21  (
    .b({_al_u5551_o,\cu_ru/m_s_epc/n2 [21]}),
    .c({wb_ins_pc[21],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6670_o}),
    .mi({ex_ins_pc[21],open_n90074}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [21],open_n90075}),
    .q({wb_ins_pc[21],\cu_ru/mepc [21]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b22|cu_ru/m_s_epc/reg1_b22  (
    .b({_al_u5547_o,\cu_ru/m_s_epc/n2 [22]}),
    .c({wb_ins_pc[22],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6668_o}),
    .mi({ex_ins_pc[22],open_n90085}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [22],open_n90097}),
    .q({wb_ins_pc[22],\cu_ru/mepc [22]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b23|cu_ru/m_s_epc/reg1_b23  (
    .b({_al_u5543_o,\cu_ru/m_s_epc/n2 [23]}),
    .c({wb_ins_pc[23],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6666_o}),
    .mi({ex_ins_pc[23],open_n90107}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [23],open_n90119}),
    .q({wb_ins_pc[23],\cu_ru/mepc [23]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b24|cu_ru/m_s_epc/reg1_b24  (
    .b({_al_u5539_o,\cu_ru/m_s_epc/n2 [24]}),
    .c({wb_ins_pc[24],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6664_o}),
    .mi({ex_ins_pc[24],open_n90136}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [24],open_n90137}),
    .q({wb_ins_pc[24],\cu_ru/mepc [24]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b25|cu_ru/m_s_epc/reg1_b25  (
    .b({_al_u5535_o,\cu_ru/m_s_epc/n2 [25]}),
    .c({wb_ins_pc[25],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6662_o}),
    .mi({ex_ins_pc[25],open_n90154}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [25],open_n90155}),
    .q({wb_ins_pc[25],\cu_ru/mepc [25]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b26|cu_ru/m_s_epc/reg1_b26  (
    .b({_al_u5531_o,\cu_ru/m_s_epc/n2 [26]}),
    .c({wb_ins_pc[26],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6660_o}),
    .mi({ex_ins_pc[26],open_n90165}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [26],open_n90177}),
    .q({wb_ins_pc[26],\cu_ru/mepc [26]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b27|cu_ru/m_s_epc/reg1_b27  (
    .b({_al_u5527_o,\cu_ru/m_s_epc/n2 [27]}),
    .c({wb_ins_pc[27],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6658_o}),
    .mi({ex_ins_pc[27],open_n90187}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [27],open_n90199}),
    .q({wb_ins_pc[27],\cu_ru/mepc [27]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b28|cu_ru/m_s_epc/reg1_b28  (
    .b({_al_u5523_o,\cu_ru/m_s_epc/n2 [28]}),
    .c({wb_ins_pc[28],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6656_o}),
    .mi({ex_ins_pc[28],open_n90216}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [28],open_n90217}),
    .q({wb_ins_pc[28],\cu_ru/mepc [28]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b29|cu_ru/m_s_epc/reg1_b29  (
    .b({_al_u5519_o,\cu_ru/m_s_epc/n2 [29]}),
    .c({wb_ins_pc[29],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6654_o}),
    .mi({ex_ins_pc[29],open_n90234}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [29],open_n90235}),
    .q({wb_ins_pc[29],\cu_ru/mepc [29]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b30|cu_ru/m_s_epc/reg1_b30  (
    .b({_al_u5511_o,\cu_ru/m_s_epc/n2 [30]}),
    .c({wb_ins_pc[30],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6650_o}),
    .mi({ex_ins_pc[30],open_n90245}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [30],open_n90257}),
    .q({wb_ins_pc[30],\cu_ru/mepc [30]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b31|cu_ru/m_s_epc/reg1_b31  (
    .b({_al_u5507_o,\cu_ru/m_s_epc/n2 [31]}),
    .c({wb_ins_pc[31],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6648_o}),
    .mi({ex_ins_pc[31],open_n90274}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [31],open_n90275}),
    .q({wb_ins_pc[31],\cu_ru/mepc [31]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b32|cu_ru/m_s_epc/reg1_b32  (
    .b({_al_u5503_o,\cu_ru/m_s_epc/n2 [32]}),
    .c({wb_ins_pc[32],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6646_o}),
    .mi({ex_ins_pc[32],open_n90292}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [32],open_n90293}),
    .q({wb_ins_pc[32],\cu_ru/mepc [32]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b33|cu_ru/m_s_epc/reg1_b33  (
    .b({_al_u5499_o,\cu_ru/m_s_epc/n2 [33]}),
    .c({wb_ins_pc[33],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6644_o}),
    .mi({ex_ins_pc[33],open_n90303}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [33],open_n90315}),
    .q({wb_ins_pc[33],\cu_ru/mepc [33]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b34|cu_ru/m_s_epc/reg1_b34  (
    .b({_al_u5495_o,\cu_ru/m_s_epc/n2 [34]}),
    .c({wb_ins_pc[34],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6642_o}),
    .mi({ex_ins_pc[34],open_n90325}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [34],open_n90337}),
    .q({wb_ins_pc[34],\cu_ru/mepc [34]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b35|cu_ru/m_s_epc/reg1_b35  (
    .b({_al_u5491_o,\cu_ru/m_s_epc/n2 [35]}),
    .c({wb_ins_pc[35],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6640_o}),
    .mi({ex_ins_pc[35],open_n90354}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [35],open_n90355}),
    .q({wb_ins_pc[35],\cu_ru/mepc [35]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b36|cu_ru/m_s_epc/reg1_b36  (
    .b({_al_u5487_o,\cu_ru/m_s_epc/n2 [36]}),
    .c({wb_ins_pc[36],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6638_o}),
    .mi({ex_ins_pc[36],open_n90372}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [36],open_n90373}),
    .q({wb_ins_pc[36],\cu_ru/mepc [36]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b37|cu_ru/m_s_epc/reg1_b37  (
    .b({_al_u5483_o,\cu_ru/m_s_epc/n2 [37]}),
    .c({wb_ins_pc[37],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6636_o}),
    .mi({ex_ins_pc[37],open_n90383}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [37],open_n90395}),
    .q({wb_ins_pc[37],\cu_ru/mepc [37]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b38|cu_ru/m_s_epc/reg1_b38  (
    .b({_al_u5479_o,\cu_ru/m_s_epc/n2 [38]}),
    .c({wb_ins_pc[38],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6634_o}),
    .mi({ex_ins_pc[38],open_n90405}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [38],open_n90417}),
    .q({wb_ins_pc[38],\cu_ru/mepc [38]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b39|cu_ru/m_s_epc/reg1_b39  (
    .b({_al_u5475_o,\cu_ru/m_s_epc/n2 [39]}),
    .c({wb_ins_pc[39],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6632_o}),
    .mi({ex_ins_pc[39],open_n90434}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [39],open_n90435}),
    .q({wb_ins_pc[39],\cu_ru/mepc [39]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b40|cu_ru/m_s_epc/reg1_b40  (
    .b({_al_u5467_o,\cu_ru/m_s_epc/n2 [40]}),
    .c({wb_ins_pc[40],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6628_o}),
    .mi({ex_ins_pc[40],open_n90445}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [40],open_n90457}),
    .q({wb_ins_pc[40],\cu_ru/mepc [40]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b41|cu_ru/m_s_epc/reg1_b41  (
    .b({_al_u5463_o,\cu_ru/m_s_epc/n2 [41]}),
    .c({wb_ins_pc[41],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6626_o}),
    .mi({ex_ins_pc[41],open_n90467}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [41],open_n90479}),
    .q({wb_ins_pc[41],\cu_ru/mepc [41]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b42|cu_ru/m_s_epc/reg1_b42  (
    .b({_al_u5459_o,\cu_ru/m_s_epc/n2 [42]}),
    .c({wb_ins_pc[42],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6624_o}),
    .mi({ex_ins_pc[42],open_n90496}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [42],open_n90497}),
    .q({wb_ins_pc[42],\cu_ru/mepc [42]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b43|cu_ru/m_s_epc/reg1_b43  (
    .b({_al_u5455_o,\cu_ru/m_s_epc/n2 [43]}),
    .c({wb_ins_pc[43],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6622_o}),
    .mi({ex_ins_pc[43],open_n90514}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [43],open_n90515}),
    .q({wb_ins_pc[43],\cu_ru/mepc [43]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b44|cu_ru/m_s_epc/reg1_b44  (
    .b({_al_u5451_o,\cu_ru/m_s_epc/n2 [44]}),
    .c({wb_ins_pc[44],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6620_o}),
    .mi({ex_ins_pc[44],open_n90525}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [44],open_n90537}),
    .q({wb_ins_pc[44],\cu_ru/mepc [44]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b45|cu_ru/m_s_epc/reg1_b45  (
    .b({_al_u5447_o,\cu_ru/m_s_epc/n2 [45]}),
    .c({wb_ins_pc[45],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6618_o}),
    .mi({ex_ins_pc[45],open_n90547}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [45],open_n90559}),
    .q({wb_ins_pc[45],\cu_ru/mepc [45]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b46|cu_ru/m_s_epc/reg1_b46  (
    .b({_al_u5443_o,\cu_ru/m_s_epc/n2 [46]}),
    .c({wb_ins_pc[46],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6616_o}),
    .mi({ex_ins_pc[46],open_n90576}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [46],open_n90577}),
    .q({wb_ins_pc[46],\cu_ru/mepc [46]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b47|cu_ru/m_s_epc/reg1_b47  (
    .b({_al_u5439_o,\cu_ru/m_s_epc/n2 [47]}),
    .c({wb_ins_pc[47],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6614_o}),
    .mi({ex_ins_pc[47],open_n90594}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [47],open_n90595}),
    .q({wb_ins_pc[47],\cu_ru/mepc [47]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b48|cu_ru/m_s_epc/reg1_b48  (
    .b({_al_u5435_o,\cu_ru/m_s_epc/n2 [48]}),
    .c({wb_ins_pc[48],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6612_o}),
    .mi({ex_ins_pc[48],open_n90605}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [48],open_n90617}),
    .q({wb_ins_pc[48],\cu_ru/mepc [48]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b49|cu_ru/m_s_epc/reg1_b49  (
    .b({_al_u5431_o,\cu_ru/m_s_epc/n2 [49]}),
    .c({wb_ins_pc[49],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6610_o}),
    .mi({ex_ins_pc[49],open_n90627}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [49],open_n90639}),
    .q({wb_ins_pc[49],\cu_ru/mepc [49]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b4|cu_ru/m_s_epc/reg1_b4  (
    .b({_al_u5471_o,\cu_ru/m_s_epc/n2 [4]}),
    .c({wb_ins_pc[4],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6608_o}),
    .mi({ex_ins_pc[4],open_n90656}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [4],open_n90657}),
    .q({wb_ins_pc[4],\cu_ru/mepc [4]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b50|cu_ru/m_s_epc/reg1_b50  (
    .b({_al_u5423_o,\cu_ru/m_s_epc/n2 [50]}),
    .c({wb_ins_pc[50],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6606_o}),
    .mi({ex_ins_pc[50],open_n90674}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [50],open_n90675}),
    .q({wb_ins_pc[50],\cu_ru/mepc [50]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b51|cu_ru/m_s_epc/reg1_b51  (
    .b({_al_u5419_o,\cu_ru/m_s_epc/n2 [51]}),
    .c({wb_ins_pc[51],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6604_o}),
    .mi({ex_ins_pc[51],open_n90685}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [51],open_n90697}),
    .q({wb_ins_pc[51],\cu_ru/mepc [51]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b52|cu_ru/m_s_epc/reg1_b52  (
    .b({_al_u5415_o,\cu_ru/m_s_epc/n2 [52]}),
    .c({wb_ins_pc[52],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6602_o}),
    .mi({ex_ins_pc[52],open_n90707}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [52],open_n90719}),
    .q({wb_ins_pc[52],\cu_ru/mepc [52]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b53|cu_ru/m_s_epc/reg1_b53  (
    .b({_al_u5411_o,\cu_ru/m_s_epc/n2 [53]}),
    .c({wb_ins_pc[53],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6600_o}),
    .mi({ex_ins_pc[53],open_n90736}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [53],open_n90737}),
    .q({wb_ins_pc[53],\cu_ru/mepc [53]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b54|cu_ru/m_s_epc/reg1_b54  (
    .b({_al_u5407_o,\cu_ru/m_s_epc/n2 [54]}),
    .c({wb_ins_pc[54],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6598_o}),
    .mi({ex_ins_pc[54],open_n90754}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [54],open_n90755}),
    .q({wb_ins_pc[54],\cu_ru/mepc [54]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b55|cu_ru/m_s_epc/reg1_b55  (
    .b({_al_u5403_o,\cu_ru/m_s_epc/n2 [55]}),
    .c({wb_ins_pc[55],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6596_o}),
    .mi({ex_ins_pc[55],open_n90765}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [55],open_n90777}),
    .q({wb_ins_pc[55],\cu_ru/mepc [55]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b56|cu_ru/m_s_epc/reg1_b56  (
    .b({_al_u5399_o,\cu_ru/m_s_epc/n2 [56]}),
    .c({wb_ins_pc[56],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6594_o}),
    .mi({ex_ins_pc[56],open_n90787}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [56],open_n90799}),
    .q({wb_ins_pc[56],\cu_ru/mepc [56]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b57|cu_ru/m_s_epc/reg1_b57  (
    .b({_al_u5395_o,\cu_ru/m_s_epc/n2 [57]}),
    .c({wb_ins_pc[57],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6592_o}),
    .mi({ex_ins_pc[57],open_n90816}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [57],open_n90817}),
    .q({wb_ins_pc[57],\cu_ru/mepc [57]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b58|cu_ru/m_s_epc/reg1_b58  (
    .b({_al_u5391_o,\cu_ru/m_s_epc/n2 [58]}),
    .c({wb_ins_pc[58],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6590_o}),
    .mi({ex_ins_pc[58],open_n90834}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [58],open_n90835}),
    .q({wb_ins_pc[58],\cu_ru/mepc [58]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b59|cu_ru/m_s_epc/reg1_b59  (
    .b({_al_u5387_o,\cu_ru/m_s_epc/n2 [59]}),
    .c({wb_ins_pc[59],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6588_o}),
    .mi({ex_ins_pc[59],open_n90845}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [59],open_n90857}),
    .q({wb_ins_pc[59],\cu_ru/mepc [59]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b5|cu_ru/m_s_epc/reg1_b5  (
    .b({_al_u5427_o,\cu_ru/m_s_epc/n2 [5]}),
    .c({wb_ins_pc[5],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6586_o}),
    .mi({ex_ins_pc[5],open_n90874}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [5],open_n90875}),
    .q({wb_ins_pc[5],\cu_ru/mepc [5]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b60|cu_ru/m_s_epc/reg1_b60  (
    .b({_al_u5379_o,\cu_ru/m_s_epc/n2 [60]}),
    .c({wb_ins_pc[60],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6584_o}),
    .mi({ex_ins_pc[60],open_n90892}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [60],open_n90893}),
    .q({wb_ins_pc[60],\cu_ru/mepc [60]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b61|cu_ru/m_s_epc/reg1_b61  (
    .b({_al_u5375_o,\cu_ru/m_s_epc/n2 [61]}),
    .c({wb_ins_pc[61],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6582_o}),
    .mi({ex_ins_pc[61],open_n90910}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [61],open_n90911}),
    .q({wb_ins_pc[61],\cu_ru/mepc [61]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b62|cu_ru/m_s_epc/reg1_b62  (
    .b({_al_u5371_o,\cu_ru/m_s_epc/n2 [62]}),
    .c({wb_ins_pc[62],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6580_o}),
    .mi({ex_ins_pc[62],open_n90921}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [62],open_n90933}),
    .q({wb_ins_pc[62],\cu_ru/mepc [62]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b63|cu_ru/m_s_epc/reg1_b63  (
    .b({_al_u5367_o,\cu_ru/m_s_epc/n2 [63]}),
    .c({wb_ins_pc[63],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6578_o}),
    .mi({ex_ins_pc[63],open_n90943}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [63],open_n90955}),
    .q({wb_ins_pc[63],\cu_ru/mepc [63]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b6|cu_ru/m_s_epc/reg1_b6  (
    .b({_al_u5383_o,\cu_ru/m_s_epc/n2 [6]}),
    .c({wb_ins_pc[6],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6576_o}),
    .mi({ex_ins_pc[6],open_n90965}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [6],open_n90977}),
    .q({wb_ins_pc[6],\cu_ru/mepc [6]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b7|cu_ru/m_s_epc/reg1_b7  (
    .b({_al_u5363_o,\cu_ru/m_s_epc/n2 [7]}),
    .c({wb_ins_pc[7],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6574_o}),
    .mi({ex_ins_pc[7],open_n90994}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [7],open_n90995}),
    .q({wb_ins_pc[7],\cu_ru/mepc [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(C*~B))"),
    //.LUT1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001111),
    .INIT_LUT1(16'b1111000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b8|cu_ru/m_s_epc/reg1_b8  (
    .b({_al_u5359_o,\cu_ru/m_s_epc/n2 [8]}),
    .c({wb_ins_pc[8],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6572_o}),
    .mi({ex_ins_pc[8],open_n91012}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [8],open_n91013}),
    .q({wb_ins_pc[8],\cu_ru/mepc [8]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(C*~B))"),
    //.LUTF1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    //.LUTG0("(~D*~(C*~B))"),
    //.LUTG1("(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000011001111),
    .INIT_LUTG1(16'b1111000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg4_b9|cu_ru/m_s_epc/reg1_b9  (
    .b({_al_u5354_o,\cu_ru/m_s_epc/n2 [9]}),
    .c({wb_ins_pc[9],\cu_ru/trap_target_m }),
    .clk(clk_pad),
    .d({_al_u5353_o,_al_u6570_o}),
    .mi({ex_ins_pc[9],open_n91023}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/n2 [9],open_n91035}),
    .q({wb_ins_pc[9],\cu_ru/mepc [9]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(358)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg5_b33|exu/reg5_b39  (
    .c({addr_ex[33],addr_ex[39]}),
    .clk(clk_pad),
    .d({ex_more_exception_neg_lutinv,ex_more_exception_neg_lutinv}),
    .sr(rst_pad),
    .q({wb_exc_code[33],wb_exc_code[39]}));  // ../../RTL/CPU/EX/exu.v(358)
  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~A)"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(D*~C*~B*~A)"),
    //.LUTG1("(~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000100000000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg6_b0|exu/reg6_b5  (
    .a({csr_index[0],csr_index[0]}),
    .b({csr_index[3],csr_index[1]}),
    .c({csr_index[4],csr_index[2]}),
    .clk(clk_pad),
    .d({csr_index[5],csr_index[5]}),
    .mi({ex_csr_index[0],ex_csr_index[5]}),
    .sr(rst_pad),
    .f({_al_u3200_o,_al_u3197_o}),
    .q({csr_index[0],csr_index[5]}));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*A)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(~D*~C*B*A)"),
    //.LUTG1("(~D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000000000001000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg6_b1|exu/reg6_b2  (
    .a({_al_u5992_o,_al_u5158_o}),
    .b({_al_u3200_o,_al_u3200_o}),
    .c({csr_index[1],csr_index[1]}),
    .clk(clk_pad),
    .d({csr_index[2],csr_index[2]}),
    .mi({ex_csr_index[1],ex_csr_index[2]}),
    .sr(rst_pad),
    .f({\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ,\cu_ru/m_s_epc/mux4_b0_sel_is_2_o }),
    .q({csr_index[1],csr_index[2]}));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(~C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg6_b3|exu/reg6_b4  (
    .a({open_n91097,csr_index[0]}),
    .b({csr_index[3],csr_index[3]}),
    .c({csr_index[4],csr_index[4]}),
    .clk(clk_pad),
    .d({_al_u3197_o,csr_index[5]}),
    .mi({ex_csr_index[3],ex_csr_index[4]}),
    .sr(rst_pad),
    .f({_al_u3198_o,_al_u3183_o}),
    .q({csr_index[3],csr_index[4]}));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg6_b7|exu/reg6_b6  (
    .a({open_n91116,_al_u3186_o}),
    .b(csr_index[7:6]),
    .c(csr_index[8:7]),
    .clk(clk_pad),
    .d({csr_index[6],csr_index[8]}),
    .mi(ex_csr_index[7:6]),
    .sr(rst_pad),
    .f({_al_u3194_o,_al_u3420_o}),
    .q(csr_index[7:6]));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg6_b9|exu/reg6_b10  (
    .a({open_n91135,_al_u3194_o}),
    .b(csr_index[11:10]),
    .c({csr_index[9],csr_index[11]}),
    .clk(clk_pad),
    .d(csr_index[10:9]),
    .mi({ex_csr_index[9],ex_csr_index[10]}),
    .sr(rst_pad),
    .f({_al_u3186_o,_al_u3252_o}),
    .q({csr_index[9],csr_index[10]}));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(383)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C@B)*~(D@A))"),
    //.LUT1("(B*A*~(D@C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000001001000001),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/reg7_b2|exu/reg7_b0  (
    .a({_al_u9183_o,id_rs1_index[3]}),
    .b({_al_u9184_o,id_rs1_index[0]}),
    .c({id_rs1_index[2],ex_rd_index[0]}),
    .clk(clk_pad),
    .d({ex_rd_index[2],ex_rd_index[3]}),
    .mi({ex_rd_index[2],ex_rd_index[0]}),
    .sr(rst_pad),
    .f({\pip_ctrl/n36_lutinv ,_al_u9184_o}),
    .q({wb_rd_index[2],wb_rd_index[0]}));  // ../../RTL/CPU/EX/exu.v(383)
  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*D)"),
    //.LUTF1("~(~(D*C)*~(B*A))"),
    //.LUTG0("(C*~B*D)"),
    //.LUTG1("~(~(D*C)*~(B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000000000000),
    .INIT_LUTF1(16'b1111100010001000),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b1111100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/st_acc_fault_reg|exu/ld_acc_fault_reg  (
    .a({load_acc_fault,open_n91164}),
    .b({_al_u2910_o,\biu/cache_ctrl_logic/statu [0]}),
    .c({_al_u2838_o,\biu/cache_ctrl_logic/statu [1]}),
    .clk(clk_pad),
    .d({_al_u2847_o,_al_u2835_o}),
    .sr(\exu/n86 ),
    .f({open_n91182,load_acc_fault}),
    .q({wb_st_acc_fault,wb_ld_acc_fault}));  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(448)
  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("~(~B*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b1111110011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \exu/st_addr_mis_reg|exu/ld_addr_mis_reg  (
    .b({\exu/store_addr_mis ,amo}),
    .c({_al_u2910_o,load}),
    .clk(clk_pad),
    .d({\exu/load_addr_mis ,_al_u3181_o}),
    .sr(\exu/n86 ),
    .f({open_n91201,\exu/load_addr_mis }),
    .q({wb_st_addr_mis,wb_ld_addr_mis}));  // ../../RTL/CPU/EX/exu.v(448)
  EG_PHY_MSLICE #(
    //.MACRO("exu/sub0/u0|exu/sub0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \exu/sub0/u0|exu/sub0/ucin  (
    .a({\exu/shift_count [0],1'b0}),
    .b({1'b1,open_n91205}),
    .f({\exu/n50 [0],open_n91225}),
    .fco(\exu/sub0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/sub0/u0|exu/sub0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \exu/sub0/u2|exu/sub0/u1  (
    .a(\exu/shift_count [2:1]),
    .b(2'b00),
    .fci(\exu/sub0/c1 ),
    .f(\exu/n50 [2:1]),
    .fco(\exu/sub0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/sub0/u0|exu/sub0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \exu/sub0/u4|exu/sub0/u3  (
    .a(\exu/shift_count [4:3]),
    .b(2'b00),
    .fci(\exu/sub0/c3 ),
    .f(\exu/n50 [4:3]),
    .fco(\exu/sub0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/sub0/u0|exu/sub0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \exu/sub0/u6|exu/sub0/u5  (
    .a(\exu/shift_count [6:5]),
    .b(2'b00),
    .fci(\exu/sub0/c5 ),
    .f(\exu/n50 [6:5]),
    .fco(\exu/sub0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("exu/sub0/u0|exu/sub0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \exu/sub0/u7_al_u9854  (
    .a({open_n91296,\exu/shift_count [7]}),
    .b({open_n91297,1'b0}),
    .fci(\exu/sub0/c7 ),
    .f({open_n91316,\exu/n50 [7]}));
  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("~(~C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/cache_reset_reg|ins_dec/cache_flush_reg  (
    .c({\ins_dec/ins_sfencevma ,\ins_dec/n35_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/ins_fence ,id_system}),
    .sr(\ins_dec/n107 ),
    .f({open_n91342,\ins_dec/ins_fence }),
    .q({cache_reset,cache_flush}));  // ../../RTL/CPU/ID/ins_dec.v(739)
  // ../../RTL/CPU/ID/ins_dec.v(830)
  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/ebreak_reg|ins_dec/ecall_reg  (
    .c({_al_u3395_o,_al_u3397_o}),
    .ce(\ins_dec/u461_sel_is_0_o ),
    .clk(clk_pad),
    .d({_al_u3391_o,_al_u3391_o}),
    .sr(\ins_dec/n107 ),
    .q({ex_ebreak,ex_ecall}));  // ../../RTL/CPU/ID/ins_dec.v(830)
  // ../../RTL/CPU/ID/ins_dec.v(830)
  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~D)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001100),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/ins_addr_mis_reg|ins_dec/int_acc_reg  (
    .b({id_ins_addr_mis,_al_u2695_o}),
    .c({id_ins_page_fault,id_int_acc}),
    .ce(\ins_dec/u461_sel_is_0_o ),
    .clk(clk_pad),
    .d({id_ins_acc_fault,id_system}),
    .mi({id_ins_addr_mis,id_int_acc}),
    .sr(\ins_dec/n107 ),
    .f({_al_u2695_o,_al_u9190_o}),
    .q({ex_ins_addr_mis,ex_int_acc}));  // ../../RTL/CPU/ID/ins_dec.v(830)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/ins_page_fault_reg  (
    .ce(\ins_dec/u461_sel_is_0_o ),
    .clk(clk_pad),
    .mi({open_n91397,id_ins_page_fault}),
    .sr(\ins_dec/n107 ),
    .q({open_n91414,ex_ins_page_fault}));  // ../../RTL/CPU/ID/ins_dec.v(830)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/mem_csr_data_xor_reg|ins_dec/mem_csr_data_max_reg  (
    .b({id_ins[29],id_ins[31]}),
    .c({_al_u3388_o,id_ins[29]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3939_o,_al_u3939_o}),
    .sr(\ins_dec/n107 ),
    .q({mem_csr_data_xor,mem_csr_data_max}));  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(D*C*B))"),
    //.LUTF1("~(~D*~C*~B*~A)"),
    //.LUTG0("~(~A*~(D*C*B))"),
    //.LUTG1("~(~D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110101010101010),
    .INIT_LUTF1(16'b1111111111111110),
    .INIT_LUTG0(16'b1110101010101010),
    .INIT_LUTG1(16'b1111111111111110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/rd_data_add_reg|ins_dec/mem_csr_data_add_reg  (
    .a({_al_u4185_o,\ins_dec/ins_addw }),
    .b({\ins_dec/ins_addw ,_al_u3939_o}),
    .c({\ins_dec/n59 ,_al_u3399_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3955_o,_al_u3384_o}),
    .sr(\ins_dec/n107 ),
    .q({rd_data_add,mem_csr_data_add}));  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*~A)"),
    //.LUTF1("(D*C*B*~A)"),
    //.LUTG0("(~D*~C*B*~A)"),
    //.LUTG1("(D*C*B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0100000000000000),
    .INIT_LUTG0(16'b0000000000000100),
    .INIT_LUTG1(16'b0100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/rd_data_and_reg|ins_dec/rd_data_xor_reg  (
    .a({_al_u3929_o,_al_u3929_o}),
    .b({_al_u3216_o,_al_u3216_o}),
    .c({_al_u3217_o,_al_u3217_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3384_o,_al_u3384_o}),
    .sr(\ins_dec/n107 ),
    .q({rd_data_and,rd_data_xor}));  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*~A)"),
    //.LUTF1("(C*~B*~D)"),
    //.LUTG0("(~D*C*B*~A)"),
    //.LUTG1("(C*~B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000001000000),
    .INIT_LUTF1(16'b0000000000110000),
    .INIT_LUTG0(16'b0000000001000000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/rd_data_slt_reg|ins_dec/rd_data_or_reg  (
    .a({open_n91480,_al_u3929_o}),
    .b({_al_u3216_o,_al_u3216_o}),
    .c({_al_u3217_o,_al_u3217_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3929_o,_al_u3384_o}),
    .sr(\ins_dec/n107 ),
    .q({rd_data_slt,rd_data_or}));  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(689)
  // ../../RTL/CPU/ID/ins_dec.v(689)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~D)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(C*~B*~D)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg0_b0|ins_dec/reg0_b1  (
    .b({_al_u3217_o,_al_u3217_o}),
    .c({_al_u3384_o,_al_u3384_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u3919_o,_al_u3919_o}),
    .sr(\ins_dec/n107 ),
    .q({ex_size[0],ex_size[1]}));  // ../../RTL/CPU/ID/ins_dec.v(689)
  // ../../RTL/CPU/ID/ins_dec.v(689)
  // ../../RTL/CPU/ID/ins_dec.v(689)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~C*~B*~A)"),
    //.LUT1("(~D*~(~C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111111110),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg0_b3|ins_dec/reg0_b2  (
    .a({open_n91525,_al_u4162_o}),
    .b({_al_u3919_o,\ins_dec/op_32_reg_lutinv }),
    .c({_al_u3217_o,\ins_dec/op_32_imm_lutinv }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/qbyte ,\ins_dec/n48_lutinv }),
    .sr(\ins_dec/n107 ),
    .f({open_n91538,\ins_dec/qbyte }),
    .q(ex_size[3:2]));  // ../../RTL/CPU/ID/ins_dec.v(689)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b1  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n91560,id_ins_pc[1]}),
    .sr(\ins_dec/n107 ),
    .q({open_n91566,ex_ins_pc[1]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b10|ins_dec/reg11_b58  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[10],id_ins_pc[58]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[10],ex_ins_pc[58]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b11|ins_dec/reg11_b8  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[11],id_ins_pc[8]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[11],ex_ins_pc[8]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b12|ins_dec/reg11_b54  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[12],id_ins_pc[54]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[12],ex_ins_pc[54]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b13|ins_dec/reg11_b53  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[13],id_ins_pc[53]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[13],ex_ins_pc[53]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b14|ins_dec/reg11_b52  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[14],id_ins_pc[52]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[14],ex_ins_pc[52]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b15|ins_dec/reg11_b49  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[15],id_ins_pc[49]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[15],ex_ins_pc[49]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b16  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n91732,id_ins_pc[16]}),
    .sr(\ins_dec/n107 ),
    .q({open_n91749,ex_ins_pc[16]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b17|ins_dec/reg11_b59  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[17],id_ins_pc[59]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[17],ex_ins_pc[59]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b18  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n91784,id_ins_pc[18]}),
    .sr(\ins_dec/n107 ),
    .q({open_n91801,ex_ins_pc[18]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b19|ins_dec/reg11_b21  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[19],id_ins_pc[21]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[19],ex_ins_pc[21]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b20  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n91843,id_ins_pc[20]}),
    .sr(\ins_dec/n107 ),
    .q({open_n91849,ex_ins_pc[20]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b22  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n91861,id_ins_pc[22]}),
    .sr(\ins_dec/n107 ),
    .q({open_n91878,ex_ins_pc[22]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b23  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n91890,id_ins_pc[23]}),
    .sr(\ins_dec/n107 ),
    .q({open_n91907,ex_ins_pc[23]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b24  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n91926,id_ins_pc[24]}),
    .sr(\ins_dec/n107 ),
    .q({open_n91932,ex_ins_pc[24]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b25|ins_dec/reg11_b51  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[25],id_ins_pc[51]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[25],ex_ins_pc[51]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b26|ins_dec/reg11_b28  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[26],id_ins_pc[28]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[26],ex_ins_pc[28]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b27  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92001,id_ins_pc[27]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92007,ex_ins_pc[27]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b29|ins_dec/reg11_b35  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[29],id_ins_pc[35]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[29],ex_ins_pc[35]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b3  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92046,id_ins_pc[3]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92063,ex_ins_pc[3]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b30|ins_dec/reg11_b46  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[30],id_ins_pc[46]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[30],ex_ins_pc[46]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b32  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92109,id_ins_pc[32]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92115,ex_ins_pc[32]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b33  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92134,id_ins_pc[33]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92140,ex_ins_pc[33]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b4  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92152,id_ins_pc[4]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92169,ex_ins_pc[4]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b42|ins_dec/reg11_b50  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({id_ins_pc[42],id_ins_pc[50]}),
    .sr(\ins_dec/n107 ),
    .q({ex_ins_pc[42],ex_ins_pc[50]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b44  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92215,id_ins_pc[44]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92221,ex_ins_pc[44]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b45  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92240,id_ins_pc[45]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92246,ex_ins_pc[45]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b47  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92258,id_ins_pc[47]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92275,ex_ins_pc[47]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b48  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92294,id_ins_pc[48]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92300,ex_ins_pc[48]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b5  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92312,id_ins_pc[5]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92329,ex_ins_pc[5]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b55  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92348,id_ins_pc[55]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92354,ex_ins_pc[55]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b56  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92373,id_ins_pc[56]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92379,ex_ins_pc[56]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b57  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92391,id_ins_pc[57]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92408,ex_ins_pc[57]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b6  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92427,id_ins_pc[6]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92433,ex_ins_pc[6]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b7  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92445,id_ins_pc[7]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92462,ex_ins_pc[7]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  EG_PHY_MSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg11_b9  (
    .ce(id_hold),
    .clk(clk_pad),
    .mi({open_n92481,id_ins_pc[9]}),
    .sr(\ins_dec/n107 ),
    .q({open_n92487,ex_ins_pc[9]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTF1("(~D*~A*~(~C*~B))"),
    //.LUTG0("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    //.LUTG1("(~D*~A*~(~C*~B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000001001100),
    .INIT_LUTF1(16'b0000000001010100),
    .INIT_LUTG0(16'b0100000001001100),
    .INIT_LUTG1(16'b0000000001010100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg5_b0|ins_dec/reg11_b0  (
    .a({_al_u7889_o,csr_data[0]}),
    .b({rs1_data[0],_al_u7141_o}),
    .c({_al_u7141_o,id_system}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/op_lui_lutinv ,id_ins_pc[0]}),
    .mi({open_n92491,id_ins_pc[0]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92503,_al_u7889_o}),
    .q({ds1[0],ex_ins_pc[0]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(~C*~D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg6_b2|ins_dec/reg9_b2  (
    .b({open_n92509,_al_u5843_o}),
    .c({_al_u5843_o,id_ins[17]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u6181_o,\ins_dec/n57_neg_lutinv }),
    .sr(\ins_dec/n107 ),
    .q({ds2[2],op_count[2]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("~(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1111000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg6_b3|ins_dec/reg9_b3  (
    .b({open_n92533,_al_u5841_o}),
    .c({_al_u5841_o,id_ins[18]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u6147_o,\ins_dec/n57_neg_lutinv }),
    .sr(\ins_dec/n107 ),
    .q({ds2[3],op_count[3]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUT1("~(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011110000),
    .INIT_LUT1(16'b1111000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg6_b4|ins_dec/reg9_b4  (
    .b({open_n92553,_al_u5839_o}),
    .c({_al_u5839_o,id_ins[19]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u6114_o,\ins_dec/n57_neg_lutinv }),
    .sr(\ins_dec/n107 ),
    .q({ds2[4],op_count[4]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTF1("~(~C*D)"),
    //.LUTG0("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG1("~(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011110000),
    .INIT_LUTF1(16'b1111000011111111),
    .INIT_LUTG0(16'b1100110011110000),
    .INIT_LUTG1(16'b1111000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg6_b5|ins_dec/reg9_b5  (
    .b({open_n92573,_al_u5837_o}),
    .c({_al_u5837_o,id_ins[20]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u5885_o,\ins_dec/n57_neg_lutinv }),
    .sr(\ins_dec/n107 ),
    .q({ds2[5],op_count[5]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("~(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1111000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg6_b6|ins_dec/reg9_b6  (
    .a({open_n92595,_al_u5144_o}),
    .b({open_n92596,\cu_ru/al_ram_gpr_al_u0_do_i0_006 }),
    .c({\ins_dec/op_count_decode [6],\cu_ru/al_ram_gpr_al_u0_do_i1_006 }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u5871_o,\cu_ru/n49 [4]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92609,\ins_dec/op_count_decode [6]}),
    .q({ds2[6],op_count[6]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    //.LUT1("~(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010000010001000),
    .INIT_LUT1(16'b1111000011111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg6_b7|ins_dec/reg9_b7  (
    .a({open_n92613,_al_u5144_o}),
    .b({open_n92614,\cu_ru/al_ram_gpr_al_u0_do_i0_007 }),
    .c({\ins_dec/op_count_decode [7],\cu_ru/al_ram_gpr_al_u0_do_i1_007 }),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u5856_o,\cu_ru/n49 [4]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92627,\ins_dec/op_count_decode [7]}),
    .q({ds2[7],op_count[7]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b31|ins_dec/reg11_b31  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[31],id_ins_pc[31]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[31],_al_u7141_o}),
    .mi({open_n92643,id_ins_pc[31]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92644,_al_u7570_o}),
    .q({as1[31],ex_ins_pc[31]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b34|ins_dec/reg11_b34  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[34],id_ins_pc[34]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[34],_al_u7141_o}),
    .mi({open_n92653,id_ins_pc[34]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92665,_al_u7682_o}),
    .q({as1[34],ex_ins_pc[34]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b36|ins_dec/reg11_b36  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[36],id_ins_pc[36]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[36],_al_u7141_o}),
    .mi({open_n92674,id_ins_pc[36]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92686,_al_u7566_o}),
    .q({as1[36],ex_ins_pc[36]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b37|ins_dec/reg11_b37  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[37],id_ins_pc[37]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[37],_al_u7141_o}),
    .mi({open_n92702,id_ins_pc[37]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92703,_al_u7562_o}),
    .q({as1[37],ex_ins_pc[37]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b38|ins_dec/reg11_b38  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[38],id_ins_pc[38]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[38],_al_u7141_o}),
    .mi({open_n92719,id_ins_pc[38]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92720,_al_u7558_o}),
    .q({as1[38],ex_ins_pc[38]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b39|ins_dec/reg11_b39  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[39],id_ins_pc[39]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[39],_al_u7141_o}),
    .mi({open_n92729,id_ins_pc[39]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92741,_al_u7554_o}),
    .q({as1[39],ex_ins_pc[39]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b40|ins_dec/reg11_b40  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[40],id_ins_pc[40]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[40],_al_u7141_o}),
    .mi({open_n92750,id_ins_pc[40]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92762,_al_u7538_o}),
    .q({as1[40],ex_ins_pc[40]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b41|ins_dec/reg11_b41  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[41],id_ins_pc[41]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[41],_al_u7141_o}),
    .mi({open_n92778,id_ins_pc[41]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92779,_al_u7534_o}),
    .q({as1[41],ex_ins_pc[41]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b43|ins_dec/reg11_b43  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[43],id_ins_pc[43]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[43],_al_u7141_o}),
    .mi({open_n92795,id_ins_pc[43]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92796,_al_u7527_o}),
    .q({as1[43],ex_ins_pc[43]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b60|ins_dec/reg11_b60  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[60],id_ins_pc[60]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[60],_al_u7141_o}),
    .mi({open_n92805,id_ins_pc[60]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92817,_al_u7523_o}),
    .q({as1[60],ex_ins_pc[60]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*~B))"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(D*~(~C*~B))"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000000000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000000000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b61|ins_dec/reg11_b61  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[61],id_ins_pc[61]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[61],_al_u7141_o}),
    .mi({open_n92826,id_ins_pc[61]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92838,_al_u7519_o}),
    .q({as1[61],ex_ins_pc[61]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b62|ins_dec/reg11_b62  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[62],id_ins_pc[62]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[62],_al_u7141_o}),
    .mi({open_n92854,id_ins_pc[62]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92855,_al_u7515_o}),
    .q({as1[62],ex_ins_pc[62]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*~B))"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg7_b63|ins_dec/reg11_b63  (
    .b({_al_u4875_o,id_system}),
    .c({id_ins_pc[63],id_ins_pc[63]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({rs1_data[63],_al_u7141_o}),
    .mi({open_n92871,id_ins_pc[63]}),
    .sr(\ins_dec/n107 ),
    .f({open_n92872,_al_u7511_o}),
    .q({as1[63],ex_ins_pc[63]}));  // ../../RTL/CPU/ID/ins_dec.v(848)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*B))"),
    //.LUTF1("~(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG0("~(~D*~(C*B))"),
    //.LUTG1("~(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111000000),
    .INIT_LUTF1(16'b1111101111101010),
    .INIT_LUTG0(16'b1111111111000000),
    .INIT_LUTG1(16'b1111101111101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg8_b11|ins_dec/reg8_b19  (
    .a({_al_u4180_o,open_n92876}),
    .b({_al_u4064_o,_al_u3214_o}),
    .c({id_ins[30],id_ins[30]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4055_o,_al_u4055_o}),
    .sr(\ins_dec/n107 ),
    .q({as2[11],as2[19]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("~(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b1111111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg8_b12|ins_dec/reg8_b18  (
    .b({_al_u3214_o,_al_u3214_o}),
    .c({id_ins[23],id_ins[29]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4055_o,_al_u4055_o}),
    .sr(\ins_dec/n107 ),
    .q({as2[12],as2[18]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("~(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b1111111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg8_b13|ins_dec/reg8_b17  (
    .b({_al_u3214_o,_al_u3214_o}),
    .c({id_ins[24],id_ins[28]}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4055_o,_al_u4055_o}),
    .sr(\ins_dec/n107 ),
    .q({as2[13],as2[17]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*B))"),
    //.LUT1("~(~D*~(C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111000000),
    .INIT_LUT1(16'b1111111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg8_b15|ins_dec/reg8_b14  (
    .b({_al_u3214_o,_al_u3214_o}),
    .c(id_ins[26:25]),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4055_o,_al_u4055_o}),
    .sr(\ins_dec/n107 ),
    .q(as2[15:14]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg8_b1|ins_dec/reg8_b2  (
    .c({_al_u4081_o,_al_u4077_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({_al_u4080_o,_al_u4076_o}),
    .sr(\ins_dec/n107 ),
    .q({as2[1],as2[2]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*~B))"),
    //.LUTF1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    //.LUTG0("(~D*~(~C*~B))"),
    //.LUTG1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011111100),
    .INIT_LUTF1(16'b1100110011110000),
    .INIT_LUTG0(16'b0000000011111100),
    .INIT_LUTG1(16'b1100110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg9_b0|ins_dec/reg6_b0  (
    .b({_al_u5847_o,_al_u5847_o}),
    .c({id_ins[15],_al_u4086_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/n57_neg_lutinv ,_al_u6213_o}),
    .sr(\ins_dec/n107 ),
    .q({op_count[0],ds2[0]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(777)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b1100110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/reg9_b1|ins_dec/reg6_b1  (
    .b({_al_u5845_o,_al_u5845_o}),
    .c({id_ins[16],_al_u4086_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/n57_neg_lutinv ,_al_u6209_o}),
    .sr(\ins_dec/n107 ),
    .q({op_count[1],ds2[1]}));  // ../../RTL/CPU/ID/ins_dec.v(777)
  // ../../RTL/CPU/ID/ins_dec.v(636)
  // ../../RTL/CPU/ID/ins_dec.v(739)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~A*~(D*C))"),
    //.LUT1("~(B*A*~(D*C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111101110111011),
    .INIT_LUT1(16'b1111011101110111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_dec/shift_r_reg|ins_dec/rd_data_ds1_reg  (
    .a({_al_u4802_o,\ins_dec/n232 }),
    .b({_al_u4806_o,_al_u7731_o}),
    .c({\ins_dec/funct7_0_lutinv ,_al_u3384_o}),
    .ce(id_hold),
    .clk(clk_pad),
    .d({\ins_dec/n38 ,_al_u3939_o}),
    .sr(\ins_dec/n107 ),
    .f({\ins_dec/n232 ,open_n93030}),
    .q({shift_r,rd_data_ds1}));  // ../../RTL/CPU/ID/ins_dec.v(636)
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/add0/u0|ins_fetch/add0/ucin  (
    .a({addr_if[2],1'b0}),
    .b({1'b1,open_n93034}),
    .ce(if_hold),
    .clk(clk_pad),
    .mi({open_n93049,addr_if[2]}),
    .sr(rst_pad),
    .f({\ins_fetch/n1 [0],open_n93050}),
    .fco(\ins_fetch/add0/c1 ),
    .q({open_n93053,id_ins_pc[2]}));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u10|ins_fetch/add0/u9  (
    .a(addr_if[12:11]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c9 ),
    .f(\ins_fetch/n1 [10:9]),
    .fco(\ins_fetch/add0/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u12|ins_fetch/add0/u11  (
    .a(addr_if[14:13]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c11 ),
    .f(\ins_fetch/n1 [12:11]),
    .fco(\ins_fetch/add0/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u14|ins_fetch/add0/u13  (
    .a(addr_if[16:15]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c13 ),
    .f(\ins_fetch/n1 [14:13]),
    .fco(\ins_fetch/add0/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u16|ins_fetch/add0/u15  (
    .a(addr_if[18:17]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c15 ),
    .f(\ins_fetch/n1 [16:15]),
    .fco(\ins_fetch/add0/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u18|ins_fetch/add0/u17  (
    .a(addr_if[20:19]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c17 ),
    .f(\ins_fetch/n1 [18:17]),
    .fco(\ins_fetch/add0/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u20|ins_fetch/add0/u19  (
    .a(addr_if[22:21]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c19 ),
    .f(\ins_fetch/n1 [20:19]),
    .fco(\ins_fetch/add0/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u22|ins_fetch/add0/u21  (
    .a(addr_if[24:23]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c21 ),
    .f(\ins_fetch/n1 [22:21]),
    .fco(\ins_fetch/add0/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u24|ins_fetch/add0/u23  (
    .a(addr_if[26:25]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c23 ),
    .f(\ins_fetch/n1 [24:23]),
    .fco(\ins_fetch/add0/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u26|ins_fetch/add0/u25  (
    .a(addr_if[28:27]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c25 ),
    .f(\ins_fetch/n1 [26:25]),
    .fco(\ins_fetch/add0/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u28|ins_fetch/add0/u27  (
    .a(addr_if[30:29]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c27 ),
    .f(\ins_fetch/n1 [28:27]),
    .fco(\ins_fetch/add0/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u2|ins_fetch/add0/u1  (
    .a(addr_if[4:3]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c1 ),
    .f(\ins_fetch/n1 [2:1]),
    .fco(\ins_fetch/add0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u30|ins_fetch/add0/u29  (
    .a(addr_if[32:31]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c29 ),
    .f(\ins_fetch/n1 [30:29]),
    .fco(\ins_fetch/add0/c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u32|ins_fetch/add0/u31  (
    .a(addr_if[34:33]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c31 ),
    .f(\ins_fetch/n1 [32:31]),
    .fco(\ins_fetch/add0/c33 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y8Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u34|ins_fetch/add0/u33  (
    .a(addr_if[36:35]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c33 ),
    .f(\ins_fetch/n1 [34:33]),
    .fco(\ins_fetch/add0/c35 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y9Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u36|ins_fetch/add0/u35  (
    .a(addr_if[38:37]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c35 ),
    .f(\ins_fetch/n1 [36:35]),
    .fco(\ins_fetch/add0/c37 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y9Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u38|ins_fetch/add0/u37  (
    .a(addr_if[40:39]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c37 ),
    .f(\ins_fetch/n1 [38:37]),
    .fco(\ins_fetch/add0/c39 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y10Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u40|ins_fetch/add0/u39  (
    .a(addr_if[42:41]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c39 ),
    .f(\ins_fetch/n1 [40:39]),
    .fco(\ins_fetch/add0/c41 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y10Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u42|ins_fetch/add0/u41  (
    .a(addr_if[44:43]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c41 ),
    .f(\ins_fetch/n1 [42:41]),
    .fco(\ins_fetch/add0/c43 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y11Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u44|ins_fetch/add0/u43  (
    .a(addr_if[46:45]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c43 ),
    .f(\ins_fetch/n1 [44:43]),
    .fco(\ins_fetch/add0/c45 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y11Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u46|ins_fetch/add0/u45  (
    .a(addr_if[48:47]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c45 ),
    .f(\ins_fetch/n1 [46:45]),
    .fco(\ins_fetch/add0/c47 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y12Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u48|ins_fetch/add0/u47  (
    .a(addr_if[50:49]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c47 ),
    .f(\ins_fetch/n1 [48:47]),
    .fco(\ins_fetch/add0/c49 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u4|ins_fetch/add0/u3  (
    .a(addr_if[6:5]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c3 ),
    .f(\ins_fetch/n1 [4:3]),
    .fco(\ins_fetch/add0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y12Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u50|ins_fetch/add0/u49  (
    .a(addr_if[52:51]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c49 ),
    .f(\ins_fetch/n1 [50:49]),
    .fco(\ins_fetch/add0/c51 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y13Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u52|ins_fetch/add0/u51  (
    .a(addr_if[54:53]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c51 ),
    .f(\ins_fetch/n1 [52:51]),
    .fco(\ins_fetch/add0/c53 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y13Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u54|ins_fetch/add0/u53  (
    .a(addr_if[56:55]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c53 ),
    .f(\ins_fetch/n1 [54:53]),
    .fco(\ins_fetch/add0/c55 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y14Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u56|ins_fetch/add0/u55  (
    .a(addr_if[58:57]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c55 ),
    .f(\ins_fetch/n1 [56:55]),
    .fco(\ins_fetch/add0/c57 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y14Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u58|ins_fetch/add0/u57  (
    .a(addr_if[60:59]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c57 ),
    .f(\ins_fetch/n1 [58:57]),
    .fco(\ins_fetch/add0/c59 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y15Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u60|ins_fetch/add0/u59  (
    .a(addr_if[62:61]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c59 ),
    .f(\ins_fetch/n1 [60:59]),
    .fco(\ins_fetch/add0/c61 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y15Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u61_al_u9855  (
    .a({open_n93670,addr_if[63]}),
    .b({open_n93671,1'b0}),
    .fci(\ins_fetch/add0/c61 ),
    .f({open_n93690,\ins_fetch/n1 [61]}));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u6|ins_fetch/add0/u5  (
    .a(addr_if[8:7]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c5 ),
    .f(\ins_fetch/n1 [6:5]),
    .fco(\ins_fetch/add0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("ins_fetch/add0/u0|ins_fetch/add0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \ins_fetch/add0/u8|ins_fetch/add0/u7  (
    .a(addr_if[10:9]),
    .b(2'b00),
    .fci(\ins_fetch/add0/c7 ),
    .f(\ins_fetch/n1 [8:7]),
    .fco(\ins_fetch/add0/c9 ));
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(137)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/ins_acc_fault_reg|ins_fetch/reg0_b32  (
    .a({open_n93740,\biu/cache_ctrl_logic/l1i_va [32]}),
    .b({open_n93741,\biu/cache_ctrl_logic/l1i_va [34]}),
    .c({_al_u2838_o,addr_if[32]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u2837_o,addr_if[34]}),
    .mi({open_n93745,addr_if[32]}),
    .sr(rst_pad),
    .f({open_n93757,_al_u9255_o}),
    .q({id_ins_acc_fault,id_ins_pc[32]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(137)
  EG_PHY_MSLICE #(
    //.LUT0("(~D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011111111),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/ins_addr_mis_reg|ins_fetch/reg0_b1  (
    .c({addr_if[1],open_n93765}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[0],if_hold}),
    .mi({open_n93776,addr_if[1]}),
    .sr(rst_pad),
    .f({open_n93777,_al_n0_en}),
    .q({id_ins_addr_mis,id_ins_pc[1]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(137)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("~(~D*~(C*B*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1111111110000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/ins_page_fault_reg|ins_fetch/reg0_b53  (
    .a({_al_u9204_o,\biu/cache_ctrl_logic/l1i_va [53]}),
    .b({_al_u9264_o,\biu/cache_ctrl_logic/l1i_va [57]}),
    .c({_al_u9265_o,addr_if[53]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u9266_o,addr_if[57]}),
    .mi({open_n93791,addr_if[53]}),
    .sr(rst_pad),
    .f({open_n93792,_al_u9237_o}),
    .q({id_ins_page_fault,id_ins_pc[53]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(137)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~B))"),
    //.LUT1("~(C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111100000000),
    .INIT_LUT1(16'b0000111111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/int_acc_reg|ins_fetch/reg0_b63  (
    .b({open_n93798,\biu/cache_ctrl_logic/l1i_va [63]}),
    .c({_al_u3250_o,addr_if[63]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({\cu_ru/mideleg_int_ctrl/n28_lutinv ,\biu/cache_ctrl_logic/l1i_value }),
    .mi({open_n93809,addr_if[63]}),
    .sr(rst_pad),
    .f({int_req,_al_u9239_o}),
    .q({id_int_acc,id_ins_pc[63]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b11|ins_fetch/reg0_b8  (
    .a({\ins_fetch/n27 ,\ins_fetch/n27 }),
    .b({pip_flush,pip_flush}),
    .c({\ins_fetch/n1 [9],\ins_fetch/n1 [6]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[11],addr_if[8]}),
    .mi({addr_if[11],addr_if[8]}),
    .sr(rst_pad),
    .f({_al_u9289_o,_al_u9306_o}),
    .q({id_ins_pc[11],id_ins_pc[8]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b14|ins_fetch/reg0_b40  (
    .a({\biu/cache_ctrl_logic/l1i_va [14],\biu/cache_ctrl_logic/l1i_va [14]}),
    .b({\biu/cache_ctrl_logic/l1i_va [22],\biu/cache_ctrl_logic/l1i_va [40]}),
    .c({addr_if[14],addr_if[14]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[22],addr_if[40]}),
    .mi({addr_if[14],addr_if[40]}),
    .sr(rst_pad),
    .f({_al_u9246_o,_al_u9224_o}),
    .q({id_ins_pc[14],id_ins_pc[40]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100110001),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b15|ins_fetch/reg0_b61  (
    .a({open_n93843,\biu/cache_ctrl_logic/l1i_va [61]}),
    .b({\biu/cache_ctrl_logic/l1i_va [15],\biu/cache_ctrl_logic/l1i_va [63]}),
    .c({addr_if[15],addr_if[61]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u9230_o,addr_if[63]}),
    .mi({addr_if[15],addr_if[61]}),
    .sr(rst_pad),
    .f({_al_u9231_o,_al_u9230_o}),
    .q({id_ins_pc[15],id_ins_pc[61]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b16|ins_fetch/reg0_b36  (
    .a({\biu/cache_ctrl_logic/l1i_va [16],\biu/cache_ctrl_logic/l1i_va [36]}),
    .b({\biu/cache_ctrl_logic/l1i_va [36],\biu/cache_ctrl_logic/l1i_va [60]}),
    .c({addr_if[16],addr_if[36]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[36],addr_if[60]}),
    .mi({addr_if[16],addr_if[36]}),
    .sr(rst_pad),
    .f({_al_u9248_o,_al_u9227_o}),
    .q({id_ins_pc[16],id_ins_pc[36]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~A*~(D@C))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~B*~A*~(D@C))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000000000001),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0001000000000001),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b18|ins_fetch/reg0_b12  (
    .a({open_n93874,_al_u9243_o}),
    .b({open_n93875,_al_u9244_o}),
    .c({addr_if[18],\biu/cache_ctrl_logic/l1i_va [12]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({\biu/cache_ctrl_logic/l1i_va [18],addr_if[12]}),
    .mi({addr_if[18],addr_if[12]}),
    .sr(rst_pad),
    .f({_al_u9243_o,_al_u9245_o}),
    .q({id_ins_pc[18],id_ins_pc[12]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b19|ins_fetch/reg0_b21  (
    .a({\biu/cache_ctrl_logic/l1i_va [19],\biu/cache_ctrl_logic/l1i_va [19]}),
    .b({\biu/cache_ctrl_logic/l1i_va [60],\biu/cache_ctrl_logic/l1i_va [21]}),
    .c({addr_if[19],addr_if[19]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[60],addr_if[21]}),
    .mi({addr_if[19],addr_if[21]}),
    .sr(rst_pad),
    .f({_al_u9226_o,_al_u9220_o}),
    .q({id_ins_pc[19],id_ins_pc[21]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b23|ins_fetch/reg0_b39  (
    .a({\biu/cache_ctrl_logic/l1i_va [23],\biu/cache_ctrl_logic/l1i_va [23]}),
    .b({\biu/cache_ctrl_logic/l1i_va [37],\biu/cache_ctrl_logic/l1i_va [39]}),
    .c({addr_if[23],addr_if[23]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[37],addr_if[39]}),
    .mi({addr_if[23],addr_if[39]}),
    .sr(rst_pad),
    .f({_al_u9217_o,_al_u9216_o}),
    .q({id_ins_pc[23],id_ins_pc[39]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b25|ins_fetch/reg0_b51  (
    .a({open_n93923,\biu/cache_ctrl_logic/l1i_va [51]}),
    .b({\biu/cache_ctrl_logic/l1i_va [25],\biu/cache_ctrl_logic/l1i_va [55]}),
    .c({addr_if[25],addr_if[51]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({_al_u9234_o,addr_if[55]}),
    .mi({addr_if[25],addr_if[51]}),
    .sr(rst_pad),
    .f({_al_u9235_o,_al_u9234_o}),
    .q({id_ins_pc[25],id_ins_pc[51]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(~(~D*B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b1010111100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b26|ins_fetch/reg0_b28  (
    .a({\biu/cache_ctrl_logic/l1i_va [26],\biu/cache_ctrl_logic/l1i_va [26]}),
    .b({\biu/cache_ctrl_logic/l1i_va [28],\biu/cache_ctrl_logic/l1i_va [28]}),
    .c({addr_if[26],addr_if[26]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[28],addr_if[28]}),
    .mi({addr_if[26],addr_if[28]}),
    .sr(rst_pad),
    .f({_al_u9262_o,_al_u9249_o}),
    .q({id_ins_pc[26],id_ins_pc[28]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b30|ins_fetch/reg0_b46  (
    .a({\biu/cache_ctrl_logic/l1i_va [30],\biu/cache_ctrl_logic/l1i_va [46]}),
    .b({\biu/cache_ctrl_logic/l1i_va [46],\biu/cache_ctrl_logic/l1i_va [50]}),
    .c({addr_if[30],addr_if[46]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[46],addr_if[50]}),
    .mi({addr_if[30],addr_if[46]}),
    .sr(rst_pad),
    .f({_al_u9261_o,_al_u9252_o}),
    .q({id_ins_pc[30],id_ins_pc[46]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b33|ins_fetch/reg0_b41  (
    .a({_al_u9239_o,\biu/cache_ctrl_logic/l1i_va [41]}),
    .b({_al_u9240_o,\biu/cache_ctrl_logic/l1i_va [47]}),
    .c({\biu/cache_ctrl_logic/l1i_va [33],addr_if[41]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[33],addr_if[47]}),
    .mi({addr_if[33],addr_if[41]}),
    .sr(rst_pad),
    .f({_al_u9241_o,_al_u9240_o}),
    .q({id_ins_pc[33],id_ins_pc[41]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b34|ins_fetch/reg0_b38  (
    .a({\biu/cache_ctrl_logic/l1i_va [34],\biu/cache_ctrl_logic/l1i_va [38]}),
    .b({\biu/cache_ctrl_logic/l1i_va [38],\biu/cache_ctrl_logic/l1i_va [40]}),
    .c({addr_if[34],addr_if[38]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[38],addr_if[40]}),
    .mi({addr_if[34],addr_if[38]}),
    .sr(rst_pad),
    .f({_al_u9247_o,_al_u9251_o}),
    .q({id_ins_pc[34],id_ins_pc[38]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b35|ins_fetch/reg0_b29  (
    .a({_al_u9212_o,\biu/cache_ctrl_logic/l1i_va [29]}),
    .b({_al_u9213_o,\biu/cache_ctrl_logic/l1i_va [31]}),
    .c({\biu/cache_ctrl_logic/l1i_va [35],addr_if[29]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[35],addr_if[31]}),
    .mi({addr_if[35],addr_if[29]}),
    .sr(rst_pad),
    .f({_al_u9214_o,_al_u9212_o}),
    .q({id_ins_pc[35],id_ins_pc[29]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b42|ins_fetch/reg0_b50  (
    .a({\biu/cache_ctrl_logic/l1i_va [42],open_n94014}),
    .b({\biu/cache_ctrl_logic/l1i_va [50],\biu/bus_unit/mmu/n19_lutinv }),
    .c({addr_if[42],addr_if[50]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[50],_al_u4501_o}),
    .mi({addr_if[42],addr_if[50]}),
    .sr(rst_pad),
    .f({_al_u9259_o,_al_u4502_o}),
    .q({id_ins_pc[42],id_ins_pc[50]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*B))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b43|ins_fetch/reg0_b45  (
    .a({\biu/cache_ctrl_logic/l1i_va [43],open_n94028}),
    .b({\biu/cache_ctrl_logic/l1i_va [45],\biu/bus_unit/mmu/n19_lutinv }),
    .c({addr_if[43],addr_if[45]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[45],_al_u4537_o}),
    .mi({addr_if[43],addr_if[45]}),
    .sr(rst_pad),
    .f({_al_u9215_o,_al_u4538_o}),
    .q({id_ins_pc[43],id_ins_pc[45]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C*B))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(D*~(C*B))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100000000),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b0011111100000000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b48|ins_fetch/reg0_b62  (
    .a({\biu/cache_ctrl_logic/l1i_va [48],open_n94042}),
    .b({\biu/cache_ctrl_logic/l1i_va [62],\biu/bus_unit/mmu/n19_lutinv }),
    .c({addr_if[48],addr_if[62]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[62],_al_u4423_o}),
    .mi({addr_if[48],addr_if[62]}),
    .sr(rst_pad),
    .f({_al_u9213_o,_al_u4424_o}),
    .q({id_ins_pc[48],id_ins_pc[62]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b49|ins_fetch/reg0_b13  (
    .a({\biu/cache_ctrl_logic/l1i_va [39],\biu/cache_ctrl_logic/l1i_va [13]}),
    .b({\biu/cache_ctrl_logic/l1i_va [49],\biu/cache_ctrl_logic/l1i_va [49]}),
    .c({addr_if[39],addr_if[13]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[49],addr_if[49]}),
    .mi({addr_if[49],addr_if[13]}),
    .sr(rst_pad),
    .f({_al_u9210_o,_al_u9206_o}),
    .q({id_ins_pc[49],id_ins_pc[13]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(95)
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(~(D*~B)*~(~C*A))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b1100010011110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg0_b59|ins_fetch/reg0_b17  (
    .a({\biu/cache_ctrl_logic/l1i_va [59],\biu/cache_ctrl_logic/l1i_va [17]}),
    .b({\biu/cache_ctrl_logic/l1i_va [61],\biu/cache_ctrl_logic/l1i_va [59]}),
    .c({addr_if[59],addr_if[17]}),
    .ce(if_hold),
    .clk(clk_pad),
    .d({addr_if[61],addr_if[59]}),
    .mi({addr_if[59],addr_if[17]}),
    .sr(rst_pad),
    .f({_al_u9232_o,_al_u9256_o}),
    .q({id_ins_pc[59],id_ins_pc[17]}));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg1_b0|ins_fetch/reg1_b9  (
    .b({ins_read[32],ins_read[41]}),
    .c({id_ins_pc[2],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({ins_read[0],ins_read[9]}),
    .sr(rst_pad),
    .f({open_n94108,\ins_fetch/ins_shift [9]}),
    .q({\ins_fetch/ins_hold [0],\ins_fetch/ins_hold [9]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg1_b10|ins_fetch/reg1_b8  (
    .b({ins_read[42],ins_read[40]}),
    .c({id_ins_pc[2],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({ins_read[10],ins_read[8]}),
    .sr(rst_pad),
    .f({\ins_fetch/ins_shift [10],\ins_fetch/ins_shift [8]}),
    .q({\ins_fetch/ins_hold [10],\ins_fetch/ins_hold [8]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg1_b11|ins_fetch/reg1_b7  (
    .b({ins_read[43],ins_read[39]}),
    .c({id_ins_pc[2],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({ins_read[11],ins_read[7]}),
    .sr(rst_pad),
    .f({\ins_fetch/ins_shift [11],\ins_fetch/ins_shift [7]}),
    .q({\ins_fetch/ins_hold [11],\ins_fetch/ins_hold [7]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg1_b12|ins_fetch/reg1_b29  (
    .b({ins_read[44],ins_read[61]}),
    .c({id_ins_pc[2],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({ins_read[12],ins_read[29]}),
    .sr(rst_pad),
    .f({\ins_fetch/ins_shift [12],\ins_fetch/ins_shift [29]}),
    .q({\ins_fetch/ins_hold [12],\ins_fetch/ins_hold [29]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg1_b13|ins_fetch/reg1_b28  (
    .b({ins_read[45],ins_read[60]}),
    .c({id_ins_pc[2],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({ins_read[13],ins_read[28]}),
    .sr(rst_pad),
    .f({\ins_fetch/ins_shift [13],\ins_fetch/ins_shift [28]}),
    .q({\ins_fetch/ins_hold [13],\ins_fetch/ins_hold [28]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg1_b14|ins_fetch/reg1_b25  (
    .b({ins_read[46],ins_read[57]}),
    .c({id_ins_pc[2],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({ins_read[14],ins_read[25]}),
    .sr(rst_pad),
    .f({\ins_fetch/ins_shift [14],\ins_fetch/ins_shift [25]}),
    .q({\ins_fetch/ins_hold [14],\ins_fetch/ins_hold [25]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  // ../../RTL/CPU/IF/ins_fetch.v(104)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \ins_fetch/reg1_b15|ins_fetch/reg1_b20  (
    .b({ins_read[47],ins_read[52]}),
    .c({id_ins_pc[2],id_ins_pc[2]}),
    .ce(\ins_fetch/n9 ),
    .clk(clk_pad),
    .d({ins_read[15],ins_read[20]}),
    .sr(rst_pad),
    .f({\ins_fetch/ins_shift [15],\ins_fetch/ins_shift [20]}),
    .q({\ins_fetch/ins_hold [15],\ins_fetch/ins_hold [20]}));  // ../../RTL/CPU/IF/ins_fetch.v(104)

endmodule 

