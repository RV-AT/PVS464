// Verilog netlist created by TD v4.5.12562
// Wed Apr  8 15:22:23 2020

`timescale 1ns / 1ps
module prv464_top  // ../../RTL/CPU/prv464_top.v(15)
  (
  cacheability_block,
  clk,
  hrdata,
  hready,
  hreset_n,
  hresp,
  m_ext_int,
  m_soft_int,
  m_time_int,
  mtime,
  rst,
  s_ext_int,
  haddr,
  hburst,
  hmastlock,
  hprot,
  hsize,
  htrans,
  hwdata,
  hwrite
  );

  input [31:0] cacheability_block;  // ../../RTL/CPU/prv464_top.v(17)
  input clk;  // ../../RTL/CPU/prv464_top.v(19)
  input [63:0] hrdata;  // ../../RTL/CPU/prv464_top.v(34)
  input hready;  // ../../RTL/CPU/prv464_top.v(31)
  input hreset_n;  // ../../RTL/CPU/prv464_top.v(33)
  input hresp;  // ../../RTL/CPU/prv464_top.v(32)
  input m_ext_int;  // ../../RTL/CPU/prv464_top.v(39)
  input m_soft_int;  // ../../RTL/CPU/prv464_top.v(38)
  input m_time_int;  // ../../RTL/CPU/prv464_top.v(37)
  input [63:0] mtime;  // ../../RTL/CPU/prv464_top.v(42)
  input rst;  // ../../RTL/CPU/prv464_top.v(20)
  input s_ext_int;  // ../../RTL/CPU/prv464_top.v(40)
  output [63:0] haddr;  // ../../RTL/CPU/prv464_top.v(22)
  output [2:0] hburst;  // ../../RTL/CPU/prv464_top.v(25)
  output hmastlock;  // ../../RTL/CPU/prv464_top.v(28)
  output [3:0] hprot;  // ../../RTL/CPU/prv464_top.v(26)
  output [2:0] hsize;  // ../../RTL/CPU/prv464_top.v(24)
  output [1:0] htrans;  // ../../RTL/CPU/prv464_top.v(27)
  output [63:0] hwdata;  // ../../RTL/CPU/prv464_top.v(29)
  output hwrite;  // ../../RTL/CPU/prv464_top.v(23)

  wire [63:0] addr_ex;  // ../../RTL/CPU/prv464_top.v(74)
  wire [63:0] addr_if;  // ../../RTL/CPU/prv464_top.v(65)
  wire [63:0] as1;  // ../../RTL/CPU/prv464_top.v(155)
  wire [63:0] as2;  // ../../RTL/CPU/prv464_top.v(156)
  wire [8:0] \biu/bus_unit/addr_counter ;  // ../../RTL/CPU/BIU/bus_unit.v(117)
  wire [8:0] \biu/bus_unit/last_addr ;  // ../../RTL/CPU/BIU/bus_unit.v(118)
  wire [1:0] \biu/bus_unit/mmu/i ;  // ../../RTL/CPU/BIU/mmu.v(94)
  wire [2:0] \biu/bus_unit/mmu/n39 ;
  wire [3:0] \biu/bus_unit/mmu/n40 ;
  wire [3:0] \biu/bus_unit/mmu/n54 ;
  wire [3:0] \biu/bus_unit/mmu/n56 ;
  wire [1:0] \biu/bus_unit/mmu/n59 ;
  wire [63:0] \biu/bus_unit/mmu/n66 ;
  wire [63:0] \biu/bus_unit/mmu/n71 ;
  wire [63:0] \biu/bus_unit/mmu/n79 ;
  wire [3:0] \biu/bus_unit/mmu/statu ;  // ../../RTL/CPU/BIU/mmu.v(95)
  wire [63:0] \biu/bus_unit/mmu_hwdata ;  // ../../RTL/CPU/BIU/bus_unit.v(106)
  wire [4:0] \biu/bus_unit/n26 ;
  wire [4:0] \biu/bus_unit/n30 ;
  wire [4:0] \biu/bus_unit/n35 ;
  wire [8:0] \biu/bus_unit/n39 ;
  wire [60:0] \biu/bus_unit/n49 ;
  wire [4:0] \biu/bus_unit/statu ;  // ../../RTL/CPU/BIU/bus_unit.v(115)
  wire [7:0] \biu/cache_ctrl_logic/ex_bsel ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(167)
  wire [127:0] \biu/cache_ctrl_logic/l1d_pa ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(143)
  wire [63:0] \biu/cache_ctrl_logic/l1d_pte ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(147)
  wire [63:0] \biu/cache_ctrl_logic/l1d_va ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(142)
  wire [127:0] \biu/cache_ctrl_logic/l1i_pa ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(141)
  wire [63:0] \biu/cache_ctrl_logic/l1i_pte ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(146)
  wire [63:0] \biu/cache_ctrl_logic/l1i_va ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(140)
  wire [4:0] \biu/cache_ctrl_logic/n100 ;
  wire [4:0] \biu/cache_ctrl_logic/n128 ;
  wire [4:0] \biu/cache_ctrl_logic/n132 ;
  wire [63:0] \biu/cache_ctrl_logic/n147 ;
  wire [63:0] \biu/cache_ctrl_logic/n158 ;
  wire [63:0] \biu/cache_ctrl_logic/n165 ;
  wire [127:0] \biu/cache_ctrl_logic/n166 ;
  wire [7:0] \biu/cache_ctrl_logic/n182 ;
  wire [6:0] \biu/cache_ctrl_logic/n185 ;
  wire [6:0] \biu/cache_ctrl_logic/n189 ;
  wire [63:0] \biu/cache_ctrl_logic/n207 ;
  wire [63:0] \biu/cache_ctrl_logic/n209 ;
  wire [63:0] \biu/cache_ctrl_logic/n212 ;
  wire [4:0] \biu/cache_ctrl_logic/n83 ;
  wire [11:0] \biu/cache_ctrl_logic/off ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(165)
  wire [127:0] \biu/cache_ctrl_logic/pa_temp ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(136)
  wire [63:0] \biu/cache_ctrl_logic/pte_temp ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(145)
  wire [4:0] \biu/cache_ctrl_logic/statu ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(133)
  wire [1:0] \biu/ex_data_sel ;  // ../../RTL/CPU/BIU/biu.v(81)
  wire [8:0] \biu/l1d_addr ;  // ../../RTL/CPU/BIU/biu.v(96)
  wire [63:0] \biu/l1d_out ;  // ../../RTL/CPU/BIU/biu.v(92)
  wire [8:0] \biu/l1i_addr ;  // ../../RTL/CPU/BIU/biu.v(95)
  wire [63:0] \biu/l1i_in ;  // ../../RTL/CPU/BIU/biu.v(91)
  wire [63:0] \biu/maddress ;  // ../../RTL/CPU/BIU/biu.v(119)
  wire [127:0] \biu/paddress ;  // ../../RTL/CPU/BIU/biu.v(120)
  wire [31:0] cacheability_block_pad;  // ../../RTL/CPU/prv464_top.v(17)
  wire [63:0] csr_data;  // ../../RTL/CPU/prv464_top.v(54)
  wire [11:0] csr_index;  // ../../RTL/CPU/prv464_top.v(180)
  wire [63:0] \cu_ru/m_cycle_event/n2 ;
  wire [63:0] \cu_ru/m_cycle_event/n4 ;
  wire [63:0] \cu_ru/m_cycle_event/n9 ;
  wire [63:0] \cu_ru/m_s_cause/n5 ;
  wire [63:0] \cu_ru/m_s_cause/n7 ;
  wire [61:0] \cu_ru/m_s_epc/n0 ;
  wire [63:0] \cu_ru/m_s_epc/n10 ;
  wire [63:0] \cu_ru/m_s_epc/n2 ;
  wire [63:0] \cu_ru/m_s_epc/n8 ;
  wire [1:0] \cu_ru/m_s_status/n47 ;
  wire [1:0] \cu_ru/m_s_status/n5 ;
  wire [3:0] \cu_ru/m_s_status/n64 ;
  wire [63:0] \cu_ru/m_s_tval/n11 ;
  wire [63:0] \cu_ru/m_s_tval/n3 ;
  wire [63:0] \cu_ru/m_s_tval/n9 ;
  wire [63:0] \cu_ru/m_sie ;  // ../../RTL/CPU/CU&RU/cu_ru.v(157)
  wire [63:0] \cu_ru/m_sip ;  // ../../RTL/CPU/CU&RU/cu_ru.v(158)
  wire [63:0] \cu_ru/mcause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(161)
  wire [63:0] \cu_ru/mcycle ;  // ../../RTL/CPU/CU&RU/cu_ru.v(170)
  wire [63:0] \cu_ru/medeleg ;  // ../../RTL/CPU/CU&RU/cu_ru.v(156)
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n98 ;
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n99 ;
  wire [63:0] \cu_ru/mepc ;  // ../../RTL/CPU/CU&RU/cu_ru.v(163)
  wire [63:0] \cu_ru/mideleg ;  // ../../RTL/CPU/CU&RU/cu_ru.v(155)
  wire [63:0] \cu_ru/minstret ;  // ../../RTL/CPU/CU&RU/cu_ru.v(171)
  wire [63:0] \cu_ru/mscratch ;  // ../../RTL/CPU/CU&RU/cu_ru.v(172)
  wire [63:0] \cu_ru/mstatus ;  // ../../RTL/CPU/CU&RU/cu_ru.v(153)
  wire [63:0] \cu_ru/mtval ;  // ../../RTL/CPU/CU&RU/cu_ru.v(165)
  wire [63:0] \cu_ru/mtvec ;  // ../../RTL/CPU/CU&RU/cu_ru.v(167)
  wire [61:0] \cu_ru/n43 ;
  wire [4:0] \cu_ru/n46 ;
  wire [4:0] \cu_ru/n49 ;
  wire [4:0] \cu_ru/n52 ;
  wire [63:0] \cu_ru/n64 ;
  wire [63:0] \cu_ru/n82 ;
  wire [63:0] \cu_ru/n84 ;
  wire [63:0] \cu_ru/n90 ;
  wire [63:0] \cu_ru/scause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(162)
  wire [63:0] \cu_ru/sepc ;  // ../../RTL/CPU/CU&RU/cu_ru.v(164)
  wire [63:0] \cu_ru/sscratch ;  // ../../RTL/CPU/CU&RU/cu_ru.v(173)
  wire [63:0] \cu_ru/stval ;  // ../../RTL/CPU/CU&RU/cu_ru.v(166)
  wire [63:0] \cu_ru/stvec ;  // ../../RTL/CPU/CU&RU/cu_ru.v(168)
  wire [63:0] \cu_ru/trap_cause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(131)
  wire [63:0] \cu_ru/tvec ;  // ../../RTL/CPU/CU&RU/cu_ru.v(133)
  wire [63:0] data_csr;  // ../../RTL/CPU/prv464_top.v(182)
  wire [63:0] data_rd;  // ../../RTL/CPU/prv464_top.v(183)
  wire [63:0] ds1;  // ../../RTL/CPU/prv464_top.v(153)
  wire [63:0] ds2;  // ../../RTL/CPU/prv464_top.v(154)
  wire [11:0] ex_csr_index;  // ../../RTL/CPU/prv464_top.v(147)
  wire [63:0] ex_exc_code;  // ../../RTL/CPU/prv464_top.v(99)
  wire [63:0] ex_ins_pc;  // ../../RTL/CPU/prv464_top.v(100)
  wire [4:0] ex_rd_index;  // ../../RTL/CPU/prv464_top.v(150)
  wire [3:0] ex_size;  // ../../RTL/CPU/prv464_top.v(133)
  wire [63:0] \exu/alu_au/add_64 ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(55)
  wire [63:0] \exu/alu_au/alu_and ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(58)
  wire [63:0] \exu/alu_au/n17 ;
  wire [63:0] \exu/alu_au/n31 ;
  wire [63:0] \exu/alu_au/n33 ;
  wire [63:0] \exu/alu_au/n35 ;
  wire [63:0] \exu/alu_au/n37 ;
  wire [63:0] \exu/alu_au/n39 ;
  wire [63:0] \exu/alu_au/n47 ;
  wire [63:0] \exu/alu_au/n53 ;
  wire [63:0] \exu/alu_au/n55 ;
  wire [63:0] \exu/alu_au/sub_64 ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(56)
  wire [63:0] \exu/alu_data_mem_csr ;  // ../../RTL/CPU/EX/exu.v(193)
  wire [63:0] \exu/lsu/n1 ;
  wire [63:0] \exu/lsu/n22 ;
  wire [47:0] \exu/lsu/n25 ;
  wire [63:0] \exu/lsu/n4 ;
  wire [63:0] \exu/lsu/n52 ;
  wire [63:0] \exu/lsu/n59 ;
  wire [3:0] \exu/main_state ;  // ../../RTL/CPU/EX/exu.v(184)
  wire [3:0] \exu/n45 ;
  wire [7:0] \exu/n50 ;
  wire [7:0] \exu/n52 ;
  wire [31:0] \exu/n54 ;
  wire [63:0] \exu/n57 ;
  wire [63:0] \exu/n64 ;
  wire [63:0] \exu/n71 ;
  wire [7:0] \exu/shift_count ;  // ../../RTL/CPU/EX/exu.v(185)
  wire [63:0] flush_pc;  // ../../RTL/CPU/prv464_top.v(61)
  wire [63:0] haddr_pad;  // ../../RTL/CPU/prv464_top.v(22)
  wire [2:0] hburst_pad;  // ../../RTL/CPU/prv464_top.v(25)
  wire [3:0] hprot_pad;  // ../../RTL/CPU/prv464_top.v(26)
  wire [63:0] hrdata_pad;  // ../../RTL/CPU/prv464_top.v(34)
  wire [2:0] hsize_pad;  // ../../RTL/CPU/prv464_top.v(24)
  wire [1:0] htrans_pad;  // ../../RTL/CPU/prv464_top.v(27)
  wire [63:0] hwdata_pad;  // ../../RTL/CPU/prv464_top.v(29)
  wire [31:0] id_ins;  // ../../RTL/CPU/prv464_top.v(90)
  wire [63:0] id_ins_pc;  // ../../RTL/CPU/prv464_top.v(91)
  wire [4:0] id_rs1_index;  // ../../RTL/CPU/prv464_top.v(57)
  wire [4:0] id_rs2_index;  // ../../RTL/CPU/prv464_top.v(59)
  wire [63:0] \ins_dec/n272 ;
  wire [63:0] \ins_dec/n284 ;
  wire [63:0] \ins_dec/n286 ;
  wire [63:0] \ins_dec/n291 ;
  wire [31:0] \ins_dec/n342 ;
  wire [7:0] \ins_dec/op_count_decode ;  // ../../RTL/CPU/ID/ins_dec.v(239)
  wire [31:0] \ins_fetch/ins_hold ;  // ../../RTL/CPU/IF/ins_fetch.v(55)
  wire [31:0] \ins_fetch/ins_shift ;  // ../../RTL/CPU/IF/ins_fetch.v(59)
  wire [61:0] \ins_fetch/n1 ;
  wire [63:0] \ins_fetch/n4 ;
  wire [63:0] ins_read;  // ../../RTL/CPU/prv464_top.v(67)
  wire [63:0] mtime_pad;  // ../../RTL/CPU/prv464_top.v(42)
  wire [63:0] new_pc;  // ../../RTL/CPU/prv464_top.v(184)
  wire [7:0] op_count;  // ../../RTL/CPU/prv464_top.v(157)
  wire [3:0] priv;  // ../../RTL/CPU/prv464_top.v(47)
  wire [63:0] rs1_data;  // ../../RTL/CPU/prv464_top.v(56)
  wire [63:0] satp;  // ../../RTL/CPU/prv464_top.v(46)
  wire [63:0] uncache_data;  // ../../RTL/CPU/prv464_top.v(77)
  wire [63:0] wb_exc_code;  // ../../RTL/CPU/prv464_top.v(185)
  wire [63:0] wb_ins_pc;  // ../../RTL/CPU/prv464_top.v(186)
  wire [4:0] wb_rd_index;  // ../../RTL/CPU/prv464_top.v(181)
  wire _al_n0_en;
  wire _al_u2659_o;
  wire _al_u2660_o;
  wire _al_u2662_o;
  wire _al_u2663_o;
  wire _al_u2667_o;
  wire _al_u2668_o;
  wire _al_u2670_o;
  wire _al_u2671_o;
  wire _al_u2674_o;
  wire _al_u2675_o;
  wire _al_u2677_o;
  wire _al_u2678_o;
  wire _al_u2680_o;
  wire _al_u2681_o;
  wire _al_u2683_o;
  wire _al_u2684_o;
  wire _al_u2691_o;
  wire _al_u2695_o;
  wire _al_u2697_o;
  wire _al_u2698_o;
  wire _al_u2703_o;
  wire _al_u2704_o;
  wire _al_u2705_o;
  wire _al_u2706_o;
  wire _al_u2707_o;
  wire _al_u2833_o;
  wire _al_u2835_o;
  wire _al_u2837_o;
  wire _al_u2838_o;
  wire _al_u2841_o;
  wire _al_u2842_o;
  wire _al_u2844_o;
  wire _al_u2845_o;
  wire _al_u2847_o;
  wire _al_u2848_o;
  wire _al_u2850_o;
  wire _al_u2852_o;
  wire _al_u2855_o;
  wire _al_u2856_o;
  wire _al_u2858_o;
  wire _al_u2860_o;
  wire _al_u2862_o;
  wire _al_u2864_o;
  wire _al_u2866_o;
  wire _al_u2868_o;
  wire _al_u2870_o;
  wire _al_u2873_o;
  wire _al_u2874_o;
  wire _al_u2885_o;
  wire _al_u2886_o;
  wire _al_u2889_o;
  wire _al_u2890_o;
  wire _al_u2891_o;
  wire _al_u2893_o;
  wire _al_u2895_o;
  wire _al_u2897_o;
  wire _al_u2899_o;
  wire _al_u2901_o;
  wire _al_u2903_o;
  wire _al_u2905_o;
  wire _al_u2907_o;
  wire _al_u2909_o;
  wire _al_u2910_o;
  wire _al_u2914_o;
  wire _al_u2915_o;
  wire _al_u2929_o;
  wire _al_u2930_o;
  wire _al_u2931_o;
  wire _al_u2932_o;
  wire _al_u2933_o;
  wire _al_u2934_o;
  wire _al_u2935_o;
  wire _al_u2936_o;
  wire _al_u2937_o;
  wire _al_u2938_o;
  wire _al_u2939_o;
  wire _al_u2940_o;
  wire _al_u2941_o;
  wire _al_u2942_o;
  wire _al_u2943_o;
  wire _al_u2944_o;
  wire _al_u2946_o;
  wire _al_u2948_o;
  wire _al_u2952_o;
  wire _al_u2954_o;
  wire _al_u2955_o;
  wire _al_u2956_o;
  wire _al_u2957_o;
  wire _al_u2958_o;
  wire _al_u2963_o;
  wire _al_u2964_o;
  wire _al_u2966_o;
  wire _al_u2974_o;
  wire _al_u2975_o;
  wire _al_u3033_o;
  wire _al_u3034_o;
  wire _al_u3043_o;
  wire _al_u3044_o;
  wire _al_u3046_o;
  wire _al_u3047_o;
  wire _al_u3049_o;
  wire _al_u3050_o;
  wire _al_u3052_o;
  wire _al_u3053_o;
  wire _al_u3055_o;
  wire _al_u3056_o;
  wire _al_u3058_o;
  wire _al_u3059_o;
  wire _al_u3061_o;
  wire _al_u3062_o;
  wire _al_u3064_o;
  wire _al_u3065_o;
  wire _al_u3067_o;
  wire _al_u3068_o;
  wire _al_u3070_o;
  wire _al_u3071_o;
  wire _al_u3073_o;
  wire _al_u3074_o;
  wire _al_u3076_o;
  wire _al_u3077_o;
  wire _al_u3079_o;
  wire _al_u3080_o;
  wire _al_u3082_o;
  wire _al_u3083_o;
  wire _al_u3085_o;
  wire _al_u3086_o;
  wire _al_u3088_o;
  wire _al_u3089_o;
  wire _al_u3091_o;
  wire _al_u3092_o;
  wire _al_u3094_o;
  wire _al_u3095_o;
  wire _al_u3097_o;
  wire _al_u3098_o;
  wire _al_u3100_o;
  wire _al_u3101_o;
  wire _al_u3103_o;
  wire _al_u3104_o;
  wire _al_u3106_o;
  wire _al_u3107_o;
  wire _al_u3109_o;
  wire _al_u3110_o;
  wire _al_u3112_o;
  wire _al_u3113_o;
  wire _al_u3115_o;
  wire _al_u3116_o;
  wire _al_u3118_o;
  wire _al_u3119_o;
  wire _al_u3121_o;
  wire _al_u3122_o;
  wire _al_u3124_o;
  wire _al_u3125_o;
  wire _al_u3127_o;
  wire _al_u3128_o;
  wire _al_u3130_o;
  wire _al_u3131_o;
  wire _al_u3133_o;
  wire _al_u3134_o;
  wire _al_u3136_o;
  wire _al_u3137_o;
  wire _al_u3139_o;
  wire _al_u3140_o;
  wire _al_u3142_o;
  wire _al_u3143_o;
  wire _al_u3145_o;
  wire _al_u3146_o;
  wire _al_u3148_o;
  wire _al_u3149_o;
  wire _al_u3152_o;
  wire _al_u3153_o;
  wire _al_u3155_o;
  wire _al_u3156_o;
  wire _al_u3158_o;
  wire _al_u3159_o;
  wire _al_u3161_o;
  wire _al_u3162_o;
  wire _al_u3164_o;
  wire _al_u3165_o;
  wire _al_u3167_o;
  wire _al_u3168_o;
  wire _al_u3170_o;
  wire _al_u3171_o;
  wire _al_u3173_o;
  wire _al_u3174_o;
  wire _al_u3179_o;
  wire _al_u3181_o;
  wire _al_u3183_o;
  wire _al_u3184_o;
  wire _al_u3185_o;
  wire _al_u3186_o;
  wire _al_u3187_o;
  wire _al_u3189_o;
  wire _al_u3190_o;
  wire _al_u3191_o;
  wire _al_u3194_o;
  wire _al_u3195_o;
  wire _al_u3197_o;
  wire _al_u3198_o;
  wire _al_u3200_o;
  wire _al_u3201_o;
  wire _al_u3204_o;
  wire _al_u3206_o;
  wire _al_u3209_o;
  wire _al_u3212_o;
  wire _al_u3213_o;
  wire _al_u3214_o;
  wire _al_u3216_o;
  wire _al_u3217_o;
  wire _al_u3222_o;
  wire _al_u3224_o;
  wire _al_u3237_o;
  wire _al_u3238_o;
  wire _al_u3240_o;
  wire _al_u3242_o;
  wire _al_u3244_o;
  wire _al_u3245_o;
  wire _al_u3248_o;
  wire _al_u3250_o;
  wire _al_u3252_o;
  wire _al_u3253_o;
  wire _al_u3254_o;
  wire _al_u3256_o;
  wire _al_u3258_o;
  wire _al_u3260_o;
  wire _al_u3262_o;
  wire _al_u3264_o;
  wire _al_u3266_o;
  wire _al_u3268_o;
  wire _al_u3270_o;
  wire _al_u3272_o;
  wire _al_u3274_o;
  wire _al_u3276_o;
  wire _al_u3278_o;
  wire _al_u3280_o;
  wire _al_u3282_o;
  wire _al_u3284_o;
  wire _al_u3286_o;
  wire _al_u3288_o;
  wire _al_u3290_o;
  wire _al_u3292_o;
  wire _al_u3294_o;
  wire _al_u3296_o;
  wire _al_u3298_o;
  wire _al_u3300_o;
  wire _al_u3302_o;
  wire _al_u3304_o;
  wire _al_u3306_o;
  wire _al_u3308_o;
  wire _al_u3310_o;
  wire _al_u3312_o;
  wire _al_u3314_o;
  wire _al_u3316_o;
  wire _al_u3318_o;
  wire _al_u3320_o;
  wire _al_u3322_o;
  wire _al_u3324_o;
  wire _al_u3326_o;
  wire _al_u3328_o;
  wire _al_u3330_o;
  wire _al_u3332_o;
  wire _al_u3334_o;
  wire _al_u3336_o;
  wire _al_u3338_o;
  wire _al_u3340_o;
  wire _al_u3342_o;
  wire _al_u3344_o;
  wire _al_u3346_o;
  wire _al_u3348_o;
  wire _al_u3350_o;
  wire _al_u3352_o;
  wire _al_u3354_o;
  wire _al_u3356_o;
  wire _al_u3358_o;
  wire _al_u3360_o;
  wire _al_u3362_o;
  wire _al_u3364_o;
  wire _al_u3366_o;
  wire _al_u3368_o;
  wire _al_u3370_o;
  wire _al_u3372_o;
  wire _al_u3374_o;
  wire _al_u3376_o;
  wire _al_u3378_o;
  wire _al_u3380_o;
  wire _al_u3382_o;
  wire _al_u3384_o;
  wire _al_u3387_o;
  wire _al_u3388_o;
  wire _al_u3391_o;
  wire _al_u3392_o;
  wire _al_u3393_o;
  wire _al_u3394_o;
  wire _al_u3395_o;
  wire _al_u3397_o;
  wire _al_u3399_o;
  wire _al_u3400_o;
  wire _al_u3403_o;
  wire _al_u3404_o;
  wire _al_u3407_o;
  wire _al_u3410_o;
  wire _al_u3411_o;
  wire _al_u3415_o;
  wire _al_u3420_o;
  wire _al_u3427_o;
  wire _al_u3430_o;
  wire _al_u3432_o;
  wire _al_u3433_o;
  wire _al_u3434_o;
  wire _al_u3441_o;
  wire _al_u3442_o;
  wire _al_u3443_o;
  wire _al_u3449_o;
  wire _al_u3450_o;
  wire _al_u3451_o;
  wire _al_u3456_o;
  wire _al_u3457_o;
  wire _al_u3459_o;
  wire _al_u3460_o;
  wire _al_u3464_o;
  wire _al_u3465_o;
  wire _al_u3467_o;
  wire _al_u3468_o;
  wire _al_u3472_o;
  wire _al_u3473_o;
  wire _al_u3475_o;
  wire _al_u3476_o;
  wire _al_u3480_o;
  wire _al_u3481_o;
  wire _al_u3483_o;
  wire _al_u3484_o;
  wire _al_u3488_o;
  wire _al_u3489_o;
  wire _al_u3490_o;
  wire _al_u3495_o;
  wire _al_u3496_o;
  wire _al_u3498_o;
  wire _al_u3499_o;
  wire _al_u3503_o;
  wire _al_u3504_o;
  wire _al_u3506_o;
  wire _al_u3507_o;
  wire _al_u3511_o;
  wire _al_u3512_o;
  wire _al_u3514_o;
  wire _al_u3515_o;
  wire _al_u3519_o;
  wire _al_u3520_o;
  wire _al_u3522_o;
  wire _al_u3523_o;
  wire _al_u3527_o;
  wire _al_u3528_o;
  wire _al_u3530_o;
  wire _al_u3531_o;
  wire _al_u3535_o;
  wire _al_u3536_o;
  wire _al_u3538_o;
  wire _al_u3539_o;
  wire _al_u3543_o;
  wire _al_u3544_o;
  wire _al_u3546_o;
  wire _al_u3547_o;
  wire _al_u3551_o;
  wire _al_u3552_o;
  wire _al_u3554_o;
  wire _al_u3555_o;
  wire _al_u3559_o;
  wire _al_u3560_o;
  wire _al_u3562_o;
  wire _al_u3563_o;
  wire _al_u3567_o;
  wire _al_u3568_o;
  wire _al_u3570_o;
  wire _al_u3571_o;
  wire _al_u3575_o;
  wire _al_u3576_o;
  wire _al_u3577_o;
  wire _al_u3582_o;
  wire _al_u3583_o;
  wire _al_u3585_o;
  wire _al_u3586_o;
  wire _al_u3590_o;
  wire _al_u3591_o;
  wire _al_u3593_o;
  wire _al_u3594_o;
  wire _al_u3598_o;
  wire _al_u3599_o;
  wire _al_u3601_o;
  wire _al_u3602_o;
  wire _al_u3606_o;
  wire _al_u3607_o;
  wire _al_u3609_o;
  wire _al_u3610_o;
  wire _al_u3614_o;
  wire _al_u3615_o;
  wire _al_u3617_o;
  wire _al_u3618_o;
  wire _al_u3622_o;
  wire _al_u3623_o;
  wire _al_u3625_o;
  wire _al_u3626_o;
  wire _al_u3630_o;
  wire _al_u3631_o;
  wire _al_u3633_o;
  wire _al_u3634_o;
  wire _al_u3638_o;
  wire _al_u3639_o;
  wire _al_u3641_o;
  wire _al_u3642_o;
  wire _al_u3646_o;
  wire _al_u3647_o;
  wire _al_u3649_o;
  wire _al_u3650_o;
  wire _al_u3654_o;
  wire _al_u3655_o;
  wire _al_u3657_o;
  wire _al_u3658_o;
  wire _al_u3662_o;
  wire _al_u3663_o;
  wire _al_u3664_o;
  wire _al_u3669_o;
  wire _al_u3670_o;
  wire _al_u3672_o;
  wire _al_u3673_o;
  wire _al_u3677_o;
  wire _al_u3678_o;
  wire _al_u3680_o;
  wire _al_u3681_o;
  wire _al_u3685_o;
  wire _al_u3686_o;
  wire _al_u3688_o;
  wire _al_u3689_o;
  wire _al_u3693_o;
  wire _al_u3694_o;
  wire _al_u3696_o;
  wire _al_u3697_o;
  wire _al_u3701_o;
  wire _al_u3702_o;
  wire _al_u3704_o;
  wire _al_u3705_o;
  wire _al_u3709_o;
  wire _al_u3710_o;
  wire _al_u3712_o;
  wire _al_u3713_o;
  wire _al_u3717_o;
  wire _al_u3718_o;
  wire _al_u3720_o;
  wire _al_u3721_o;
  wire _al_u3725_o;
  wire _al_u3726_o;
  wire _al_u3728_o;
  wire _al_u3729_o;
  wire _al_u3733_o;
  wire _al_u3734_o;
  wire _al_u3735_o;
  wire _al_u3740_o;
  wire _al_u3741_o;
  wire _al_u3742_o;
  wire _al_u3747_o;
  wire _al_u3748_o;
  wire _al_u3749_o;
  wire _al_u3754_o;
  wire _al_u3755_o;
  wire _al_u3756_o;
  wire _al_u3761_o;
  wire _al_u3762_o;
  wire _al_u3763_o;
  wire _al_u3768_o;
  wire _al_u3769_o;
  wire _al_u3770_o;
  wire _al_u3775_o;
  wire _al_u3776_o;
  wire _al_u3777_o;
  wire _al_u3782_o;
  wire _al_u3783_o;
  wire _al_u3784_o;
  wire _al_u3789_o;
  wire _al_u3790_o;
  wire _al_u3791_o;
  wire _al_u3796_o;
  wire _al_u3797_o;
  wire _al_u3798_o;
  wire _al_u3803_o;
  wire _al_u3804_o;
  wire _al_u3805_o;
  wire _al_u3810_o;
  wire _al_u3811_o;
  wire _al_u3812_o;
  wire _al_u3817_o;
  wire _al_u3818_o;
  wire _al_u3819_o;
  wire _al_u3824_o;
  wire _al_u3825_o;
  wire _al_u3826_o;
  wire _al_u3831_o;
  wire _al_u3832_o;
  wire _al_u3833_o;
  wire _al_u3838_o;
  wire _al_u3839_o;
  wire _al_u3840_o;
  wire _al_u3845_o;
  wire _al_u3846_o;
  wire _al_u3847_o;
  wire _al_u3852_o;
  wire _al_u3853_o;
  wire _al_u3854_o;
  wire _al_u3859_o;
  wire _al_u3860_o;
  wire _al_u3861_o;
  wire _al_u3866_o;
  wire _al_u3867_o;
  wire _al_u3868_o;
  wire _al_u3874_o;
  wire _al_u3875_o;
  wire _al_u3876_o;
  wire _al_u3882_o;
  wire _al_u3883_o;
  wire _al_u3884_o;
  wire _al_u3890_o;
  wire _al_u3891_o;
  wire _al_u3892_o;
  wire _al_u3898_o;
  wire _al_u3899_o;
  wire _al_u3900_o;
  wire _al_u3906_o;
  wire _al_u3907_o;
  wire _al_u3908_o;
  wire _al_u3913_o;
  wire _al_u3914_o;
  wire _al_u3915_o;
  wire _al_u3919_o;
  wire _al_u3923_o;
  wire _al_u3924_o;
  wire _al_u3925_o;
  wire _al_u3926_o;
  wire _al_u3927_o;
  wire _al_u3928_o;
  wire _al_u3929_o;
  wire _al_u3932_o;
  wire _al_u3938_o;
  wire _al_u3939_o;
  wire _al_u3944_o;
  wire _al_u3945_o;
  wire _al_u3947_o;
  wire _al_u3950_o;
  wire _al_u3955_o;
  wire _al_u3956_o;
  wire _al_u3969_o;
  wire _al_u3972_o;
  wire _al_u4055_o;
  wire _al_u4064_o;
  wire _al_u4066_o;
  wire _al_u4067_o;
  wire _al_u4069_o;
  wire _al_u4071_o;
  wire _al_u4072_o;
  wire _al_u4073_o;
  wire _al_u4075_o;
  wire _al_u4076_o;
  wire _al_u4077_o;
  wire _al_u4079_o;
  wire _al_u4080_o;
  wire _al_u4081_o;
  wire _al_u4083_o;
  wire _al_u4084_o;
  wire _al_u4086_o;
  wire _al_u4092_o;
  wire _al_u4094_o;
  wire _al_u4099_o;
  wire _al_u4100_o;
  wire _al_u4101_o;
  wire _al_u4106_o;
  wire _al_u4107_o;
  wire _al_u4108_o;
  wire _al_u4113_o;
  wire _al_u4117_o;
  wire _al_u4119_o;
  wire _al_u4121_o;
  wire _al_u4122_o;
  wire _al_u4123_o;
  wire _al_u4126_o;
  wire _al_u4127_o;
  wire _al_u4128_o;
  wire _al_u4131_o;
  wire _al_u4132_o;
  wire _al_u4133_o;
  wire _al_u4134_o;
  wire _al_u4135_o;
  wire _al_u4136_o;
  wire _al_u4137_o;
  wire _al_u4138_o;
  wire _al_u4139_o;
  wire _al_u4140_o;
  wire _al_u4141_o;
  wire _al_u4142_o;
  wire _al_u4143_o;
  wire _al_u4161_o;
  wire _al_u4162_o;
  wire _al_u4165_o;
  wire _al_u4166_o;
  wire _al_u4167_o;
  wire _al_u4169_o;
  wire _al_u4170_o;
  wire _al_u4172_o;
  wire _al_u4173_o;
  wire _al_u4175_o;
  wire _al_u4177_o;
  wire _al_u4178_o;
  wire _al_u4180_o;
  wire _al_u4182_o;
  wire _al_u4183_o;
  wire _al_u4185_o;
  wire _al_u4191_o;
  wire _al_u4192_o;
  wire _al_u4193_o;
  wire _al_u4194_o;
  wire _al_u4195_o;
  wire _al_u4197_o;
  wire _al_u4199_o;
  wire _al_u4200_o;
  wire _al_u4201_o;
  wire _al_u4203_o;
  wire _al_u4205_o;
  wire _al_u4207_o;
  wire _al_u4208_o;
  wire _al_u4210_o;
  wire _al_u4211_o;
  wire _al_u4213_o;
  wire _al_u4214_o;
  wire _al_u4216_o;
  wire _al_u4217_o;
  wire _al_u4219_o;
  wire _al_u4220_o;
  wire _al_u4222_o;
  wire _al_u4223_o;
  wire _al_u4225_o;
  wire _al_u4226_o;
  wire _al_u4229_o;
  wire _al_u4230_o;
  wire _al_u4232_o;
  wire _al_u4233_o;
  wire _al_u4234_o;
  wire _al_u4236_o;
  wire _al_u4237_o;
  wire _al_u4238_o;
  wire _al_u4240_o;
  wire _al_u4241_o;
  wire _al_u4242_o;
  wire _al_u4244_o;
  wire _al_u4245_o;
  wire _al_u4246_o;
  wire _al_u4248_o;
  wire _al_u4249_o;
  wire _al_u4250_o;
  wire _al_u4252_o;
  wire _al_u4253_o;
  wire _al_u4254_o;
  wire _al_u4256_o;
  wire _al_u4257_o;
  wire _al_u4258_o;
  wire _al_u4260_o;
  wire _al_u4261_o;
  wire _al_u4262_o;
  wire _al_u4264_o;
  wire _al_u4265_o;
  wire _al_u4266_o;
  wire _al_u4268_o;
  wire _al_u4269_o;
  wire _al_u4270_o;
  wire _al_u4272_o;
  wire _al_u4273_o;
  wire _al_u4274_o;
  wire _al_u4276_o;
  wire _al_u4277_o;
  wire _al_u4278_o;
  wire _al_u4280_o;
  wire _al_u4281_o;
  wire _al_u4282_o;
  wire _al_u4284_o;
  wire _al_u4285_o;
  wire _al_u4286_o;
  wire _al_u4288_o;
  wire _al_u4289_o;
  wire _al_u4290_o;
  wire _al_u4292_o;
  wire _al_u4293_o;
  wire _al_u4294_o;
  wire _al_u4296_o;
  wire _al_u4297_o;
  wire _al_u4298_o;
  wire _al_u4300_o;
  wire _al_u4301_o;
  wire _al_u4302_o;
  wire _al_u4304_o;
  wire _al_u4305_o;
  wire _al_u4306_o;
  wire _al_u4308_o;
  wire _al_u4309_o;
  wire _al_u4310_o;
  wire _al_u4312_o;
  wire _al_u4313_o;
  wire _al_u4314_o;
  wire _al_u4316_o;
  wire _al_u4317_o;
  wire _al_u4318_o;
  wire _al_u4320_o;
  wire _al_u4321_o;
  wire _al_u4322_o;
  wire _al_u4324_o;
  wire _al_u4325_o;
  wire _al_u4326_o;
  wire _al_u4328_o;
  wire _al_u4329_o;
  wire _al_u4330_o;
  wire _al_u4332_o;
  wire _al_u4333_o;
  wire _al_u4334_o;
  wire _al_u4336_o;
  wire _al_u4337_o;
  wire _al_u4338_o;
  wire _al_u4340_o;
  wire _al_u4341_o;
  wire _al_u4342_o;
  wire _al_u4344_o;
  wire _al_u4345_o;
  wire _al_u4346_o;
  wire _al_u4348_o;
  wire _al_u4349_o;
  wire _al_u4350_o;
  wire _al_u4352_o;
  wire _al_u4353_o;
  wire _al_u4354_o;
  wire _al_u4356_o;
  wire _al_u4357_o;
  wire _al_u4358_o;
  wire _al_u4360_o;
  wire _al_u4361_o;
  wire _al_u4362_o;
  wire _al_u4364_o;
  wire _al_u4365_o;
  wire _al_u4366_o;
  wire _al_u4368_o;
  wire _al_u4369_o;
  wire _al_u4370_o;
  wire _al_u4372_o;
  wire _al_u4373_o;
  wire _al_u4374_o;
  wire _al_u4376_o;
  wire _al_u4377_o;
  wire _al_u4378_o;
  wire _al_u4380_o;
  wire _al_u4381_o;
  wire _al_u4382_o;
  wire _al_u4384_o;
  wire _al_u4385_o;
  wire _al_u4386_o;
  wire _al_u4388_o;
  wire _al_u4389_o;
  wire _al_u4390_o;
  wire _al_u4392_o;
  wire _al_u4393_o;
  wire _al_u4394_o;
  wire _al_u4397_o;
  wire _al_u4398_o;
  wire _al_u4399_o;
  wire _al_u4400_o;
  wire _al_u4401_o;
  wire _al_u4402_o;
  wire _al_u4403_o;
  wire _al_u4405_o;
  wire _al_u4406_o;
  wire _al_u4407_o;
  wire _al_u4408_o;
  wire _al_u4409_o;
  wire _al_u4411_o;
  wire _al_u4412_o;
  wire _al_u4413_o;
  wire _al_u4414_o;
  wire _al_u4415_o;
  wire _al_u4417_o;
  wire _al_u4418_o;
  wire _al_u4419_o;
  wire _al_u4420_o;
  wire _al_u4421_o;
  wire _al_u4423_o;
  wire _al_u4424_o;
  wire _al_u4425_o;
  wire _al_u4426_o;
  wire _al_u4427_o;
  wire _al_u4429_o;
  wire _al_u4430_o;
  wire _al_u4431_o;
  wire _al_u4432_o;
  wire _al_u4433_o;
  wire _al_u4435_o;
  wire _al_u4436_o;
  wire _al_u4437_o;
  wire _al_u4438_o;
  wire _al_u4439_o;
  wire _al_u4441_o;
  wire _al_u4442_o;
  wire _al_u4443_o;
  wire _al_u4444_o;
  wire _al_u4445_o;
  wire _al_u4447_o;
  wire _al_u4448_o;
  wire _al_u4449_o;
  wire _al_u4450_o;
  wire _al_u4451_o;
  wire _al_u4453_o;
  wire _al_u4454_o;
  wire _al_u4455_o;
  wire _al_u4456_o;
  wire _al_u4457_o;
  wire _al_u4459_o;
  wire _al_u4460_o;
  wire _al_u4461_o;
  wire _al_u4462_o;
  wire _al_u4463_o;
  wire _al_u4465_o;
  wire _al_u4466_o;
  wire _al_u4467_o;
  wire _al_u4468_o;
  wire _al_u4469_o;
  wire _al_u4471_o;
  wire _al_u4472_o;
  wire _al_u4473_o;
  wire _al_u4474_o;
  wire _al_u4475_o;
  wire _al_u4477_o;
  wire _al_u4478_o;
  wire _al_u4479_o;
  wire _al_u4480_o;
  wire _al_u4481_o;
  wire _al_u4483_o;
  wire _al_u4484_o;
  wire _al_u4485_o;
  wire _al_u4486_o;
  wire _al_u4487_o;
  wire _al_u4489_o;
  wire _al_u4490_o;
  wire _al_u4491_o;
  wire _al_u4492_o;
  wire _al_u4493_o;
  wire _al_u4495_o;
  wire _al_u4496_o;
  wire _al_u4497_o;
  wire _al_u4498_o;
  wire _al_u4499_o;
  wire _al_u4501_o;
  wire _al_u4502_o;
  wire _al_u4503_o;
  wire _al_u4504_o;
  wire _al_u4505_o;
  wire _al_u4507_o;
  wire _al_u4508_o;
  wire _al_u4509_o;
  wire _al_u4510_o;
  wire _al_u4511_o;
  wire _al_u4513_o;
  wire _al_u4514_o;
  wire _al_u4515_o;
  wire _al_u4516_o;
  wire _al_u4517_o;
  wire _al_u4519_o;
  wire _al_u4520_o;
  wire _al_u4521_o;
  wire _al_u4522_o;
  wire _al_u4523_o;
  wire _al_u4525_o;
  wire _al_u4526_o;
  wire _al_u4527_o;
  wire _al_u4528_o;
  wire _al_u4529_o;
  wire _al_u4531_o;
  wire _al_u4532_o;
  wire _al_u4533_o;
  wire _al_u4534_o;
  wire _al_u4535_o;
  wire _al_u4537_o;
  wire _al_u4538_o;
  wire _al_u4539_o;
  wire _al_u4540_o;
  wire _al_u4541_o;
  wire _al_u4543_o;
  wire _al_u4544_o;
  wire _al_u4545_o;
  wire _al_u4546_o;
  wire _al_u4547_o;
  wire _al_u4549_o;
  wire _al_u4550_o;
  wire _al_u4551_o;
  wire _al_u4552_o;
  wire _al_u4553_o;
  wire _al_u4555_o;
  wire _al_u4556_o;
  wire _al_u4557_o;
  wire _al_u4558_o;
  wire _al_u4559_o;
  wire _al_u4561_o;
  wire _al_u4562_o;
  wire _al_u4563_o;
  wire _al_u4564_o;
  wire _al_u4565_o;
  wire _al_u4567_o;
  wire _al_u4568_o;
  wire _al_u4569_o;
  wire _al_u4570_o;
  wire _al_u4571_o;
  wire _al_u4573_o;
  wire _al_u4574_o;
  wire _al_u4575_o;
  wire _al_u4576_o;
  wire _al_u4577_o;
  wire _al_u4579_o;
  wire _al_u4580_o;
  wire _al_u4581_o;
  wire _al_u4582_o;
  wire _al_u4583_o;
  wire _al_u4585_o;
  wire _al_u4586_o;
  wire _al_u4587_o;
  wire _al_u4588_o;
  wire _al_u4589_o;
  wire _al_u4591_o;
  wire _al_u4592_o;
  wire _al_u4593_o;
  wire _al_u4594_o;
  wire _al_u4595_o;
  wire _al_u4597_o;
  wire _al_u4598_o;
  wire _al_u4599_o;
  wire _al_u4600_o;
  wire _al_u4601_o;
  wire _al_u4603_o;
  wire _al_u4604_o;
  wire _al_u4605_o;
  wire _al_u4606_o;
  wire _al_u4607_o;
  wire _al_u4609_o;
  wire _al_u4610_o;
  wire _al_u4611_o;
  wire _al_u4612_o;
  wire _al_u4613_o;
  wire _al_u4615_o;
  wire _al_u4616_o;
  wire _al_u4617_o;
  wire _al_u4618_o;
  wire _al_u4619_o;
  wire _al_u4621_o;
  wire _al_u4622_o;
  wire _al_u4623_o;
  wire _al_u4624_o;
  wire _al_u4625_o;
  wire _al_u4627_o;
  wire _al_u4628_o;
  wire _al_u4629_o;
  wire _al_u4630_o;
  wire _al_u4631_o;
  wire _al_u4633_o;
  wire _al_u4634_o;
  wire _al_u4635_o;
  wire _al_u4636_o;
  wire _al_u4637_o;
  wire _al_u4639_o;
  wire _al_u4640_o;
  wire _al_u4641_o;
  wire _al_u4642_o;
  wire _al_u4643_o;
  wire _al_u4645_o;
  wire _al_u4646_o;
  wire _al_u4647_o;
  wire _al_u4648_o;
  wire _al_u4649_o;
  wire _al_u4651_o;
  wire _al_u4652_o;
  wire _al_u4653_o;
  wire _al_u4654_o;
  wire _al_u4655_o;
  wire _al_u4657_o;
  wire _al_u4658_o;
  wire _al_u4659_o;
  wire _al_u4660_o;
  wire _al_u4661_o;
  wire _al_u4663_o;
  wire _al_u4664_o;
  wire _al_u4665_o;
  wire _al_u4666_o;
  wire _al_u4667_o;
  wire _al_u4669_o;
  wire _al_u4670_o;
  wire _al_u4671_o;
  wire _al_u4672_o;
  wire _al_u4673_o;
  wire _al_u4675_o;
  wire _al_u4676_o;
  wire _al_u4677_o;
  wire _al_u4678_o;
  wire _al_u4679_o;
  wire _al_u4681_o;
  wire _al_u4682_o;
  wire _al_u4683_o;
  wire _al_u4684_o;
  wire _al_u4685_o;
  wire _al_u4687_o;
  wire _al_u4688_o;
  wire _al_u4689_o;
  wire _al_u4690_o;
  wire _al_u4691_o;
  wire _al_u4693_o;
  wire _al_u4694_o;
  wire _al_u4695_o;
  wire _al_u4696_o;
  wire _al_u4697_o;
  wire _al_u4699_o;
  wire _al_u4700_o;
  wire _al_u4701_o;
  wire _al_u4702_o;
  wire _al_u4703_o;
  wire _al_u4705_o;
  wire _al_u4706_o;
  wire _al_u4707_o;
  wire _al_u4708_o;
  wire _al_u4709_o;
  wire _al_u4711_o;
  wire _al_u4712_o;
  wire _al_u4713_o;
  wire _al_u4714_o;
  wire _al_u4715_o;
  wire _al_u4717_o;
  wire _al_u4718_o;
  wire _al_u4719_o;
  wire _al_u4720_o;
  wire _al_u4721_o;
  wire _al_u4723_o;
  wire _al_u4724_o;
  wire _al_u4725_o;
  wire _al_u4726_o;
  wire _al_u4727_o;
  wire _al_u4729_o;
  wire _al_u4730_o;
  wire _al_u4731_o;
  wire _al_u4732_o;
  wire _al_u4733_o;
  wire _al_u4735_o;
  wire _al_u4736_o;
  wire _al_u4737_o;
  wire _al_u4738_o;
  wire _al_u4739_o;
  wire _al_u4741_o;
  wire _al_u4742_o;
  wire _al_u4743_o;
  wire _al_u4744_o;
  wire _al_u4745_o;
  wire _al_u4747_o;
  wire _al_u4748_o;
  wire _al_u4749_o;
  wire _al_u4750_o;
  wire _al_u4751_o;
  wire _al_u4753_o;
  wire _al_u4754_o;
  wire _al_u4755_o;
  wire _al_u4756_o;
  wire _al_u4757_o;
  wire _al_u4759_o;
  wire _al_u4760_o;
  wire _al_u4761_o;
  wire _al_u4762_o;
  wire _al_u4763_o;
  wire _al_u4765_o;
  wire _al_u4766_o;
  wire _al_u4768_o;
  wire _al_u4769_o;
  wire _al_u4770_o;
  wire _al_u4772_o;
  wire _al_u4773_o;
  wire _al_u4774_o;
  wire _al_u4776_o;
  wire _al_u4777_o;
  wire _al_u4778_o;
  wire _al_u4780_o;
  wire _al_u4781_o;
  wire _al_u4782_o;
  wire _al_u4784_o;
  wire _al_u4785_o;
  wire _al_u4786_o;
  wire _al_u4788_o;
  wire _al_u4789_o;
  wire _al_u4790_o;
  wire _al_u4792_o;
  wire _al_u4793_o;
  wire _al_u4794_o;
  wire _al_u4796_o;
  wire _al_u4797_o;
  wire _al_u4798_o;
  wire _al_u4801_o;
  wire _al_u4802_o;
  wire _al_u4804_o;
  wire _al_u4806_o;
  wire _al_u4808_o;
  wire _al_u4809_o;
  wire _al_u4810_o;
  wire _al_u4811_o;
  wire _al_u4812_o;
  wire _al_u4813_o;
  wire _al_u4815_o;
  wire _al_u4816_o;
  wire _al_u4817_o;
  wire _al_u4818_o;
  wire _al_u4819_o;
  wire _al_u4820_o;
  wire _al_u4822_o;
  wire _al_u4823_o;
  wire _al_u4824_o;
  wire _al_u4825_o;
  wire _al_u4826_o;
  wire _al_u4827_o;
  wire _al_u4829_o;
  wire _al_u4830_o;
  wire _al_u4831_o;
  wire _al_u4832_o;
  wire _al_u4833_o;
  wire _al_u4834_o;
  wire _al_u4835_o;
  wire _al_u4837_o;
  wire _al_u4838_o;
  wire _al_u4840_o;
  wire _al_u4841_o;
  wire _al_u4842_o;
  wire _al_u4844_o;
  wire _al_u4845_o;
  wire _al_u4846_o;
  wire _al_u4848_o;
  wire _al_u4849_o;
  wire _al_u4850_o;
  wire _al_u4852_o;
  wire _al_u4853_o;
  wire _al_u4854_o;
  wire _al_u4856_o;
  wire _al_u4857_o;
  wire _al_u4858_o;
  wire _al_u4860_o;
  wire _al_u4861_o;
  wire _al_u4862_o;
  wire _al_u4864_o;
  wire _al_u4865_o;
  wire _al_u4866_o;
  wire _al_u4868_o;
  wire _al_u4869_o;
  wire _al_u4870_o;
  wire _al_u4872_o;
  wire _al_u4875_o;
  wire _al_u5003_o;
  wire _al_u5005_o;
  wire _al_u5007_o;
  wire _al_u5009_o;
  wire _al_u5011_o;
  wire _al_u5013_o;
  wire _al_u5015_o;
  wire _al_u5017_o;
  wire _al_u5019_o;
  wire _al_u5020_o;
  wire _al_u5022_o;
  wire _al_u5023_o;
  wire _al_u5025_o;
  wire _al_u5026_o;
  wire _al_u5028_o;
  wire _al_u5029_o;
  wire _al_u5031_o;
  wire _al_u5032_o;
  wire _al_u5034_o;
  wire _al_u5035_o;
  wire _al_u5037_o;
  wire _al_u5038_o;
  wire _al_u5040_o;
  wire _al_u5041_o;
  wire _al_u5043_o;
  wire _al_u5044_o;
  wire _al_u5046_o;
  wire _al_u5047_o;
  wire _al_u5049_o;
  wire _al_u5050_o;
  wire _al_u5052_o;
  wire _al_u5053_o;
  wire _al_u5055_o;
  wire _al_u5056_o;
  wire _al_u5058_o;
  wire _al_u5059_o;
  wire _al_u5061_o;
  wire _al_u5062_o;
  wire _al_u5064_o;
  wire _al_u5065_o;
  wire _al_u5067_o;
  wire _al_u5068_o;
  wire _al_u5070_o;
  wire _al_u5071_o;
  wire _al_u5073_o;
  wire _al_u5074_o;
  wire _al_u5076_o;
  wire _al_u5077_o;
  wire _al_u5079_o;
  wire _al_u5080_o;
  wire _al_u5082_o;
  wire _al_u5083_o;
  wire _al_u5085_o;
  wire _al_u5086_o;
  wire _al_u5088_o;
  wire _al_u5089_o;
  wire _al_u5091_o;
  wire _al_u5092_o;
  wire _al_u5094_o;
  wire _al_u5095_o;
  wire _al_u5098_o;
  wire _al_u5099_o;
  wire _al_u5100_o;
  wire _al_u5101_o;
  wire _al_u5102_o;
  wire _al_u5104_o;
  wire _al_u5105_o;
  wire _al_u5106_o;
  wire _al_u5107_o;
  wire _al_u5108_o;
  wire _al_u5110_o;
  wire _al_u5111_o;
  wire _al_u5112_o;
  wire _al_u5114_o;
  wire _al_u5115_o;
  wire _al_u5116_o;
  wire _al_u5118_o;
  wire _al_u5119_o;
  wire _al_u5120_o;
  wire _al_u5122_o;
  wire _al_u5123_o;
  wire _al_u5124_o;
  wire _al_u5126_o;
  wire _al_u5127_o;
  wire _al_u5128_o;
  wire _al_u5130_o;
  wire _al_u5131_o;
  wire _al_u5132_o;
  wire _al_u5134_o;
  wire _al_u5135_o;
  wire _al_u5136_o;
  wire _al_u5138_o;
  wire _al_u5139_o;
  wire _al_u5140_o;
  wire _al_u5142_o;
  wire _al_u5143_o;
  wire _al_u5144_o;
  wire _al_u5147_o;
  wire _al_u5149_o;
  wire _al_u5151_o;
  wire _al_u5152_o;
  wire _al_u5154_o;
  wire _al_u5155_o;
  wire _al_u5156_o;
  wire _al_u5157_o;
  wire _al_u5158_o;
  wire _al_u5160_o;
  wire _al_u5161_o;
  wire _al_u5164_o;
  wire _al_u5167_o;
  wire _al_u5170_o;
  wire _al_u5173_o;
  wire _al_u5176_o;
  wire _al_u5179_o;
  wire _al_u5182_o;
  wire _al_u5185_o;
  wire _al_u5188_o;
  wire _al_u5191_o;
  wire _al_u5194_o;
  wire _al_u5197_o;
  wire _al_u5200_o;
  wire _al_u5203_o;
  wire _al_u5206_o;
  wire _al_u5209_o;
  wire _al_u5212_o;
  wire _al_u5215_o;
  wire _al_u5218_o;
  wire _al_u5221_o;
  wire _al_u5224_o;
  wire _al_u5227_o;
  wire _al_u5230_o;
  wire _al_u5233_o;
  wire _al_u5236_o;
  wire _al_u5239_o;
  wire _al_u5242_o;
  wire _al_u5245_o;
  wire _al_u5248_o;
  wire _al_u5251_o;
  wire _al_u5254_o;
  wire _al_u5257_o;
  wire _al_u5260_o;
  wire _al_u5263_o;
  wire _al_u5266_o;
  wire _al_u5269_o;
  wire _al_u5272_o;
  wire _al_u5275_o;
  wire _al_u5278_o;
  wire _al_u5281_o;
  wire _al_u5284_o;
  wire _al_u5287_o;
  wire _al_u5290_o;
  wire _al_u5293_o;
  wire _al_u5296_o;
  wire _al_u5299_o;
  wire _al_u5302_o;
  wire _al_u5305_o;
  wire _al_u5308_o;
  wire _al_u5311_o;
  wire _al_u5314_o;
  wire _al_u5317_o;
  wire _al_u5320_o;
  wire _al_u5323_o;
  wire _al_u5326_o;
  wire _al_u5329_o;
  wire _al_u5332_o;
  wire _al_u5335_o;
  wire _al_u5338_o;
  wire _al_u5341_o;
  wire _al_u5344_o;
  wire _al_u5347_o;
  wire _al_u5350_o;
  wire _al_u5353_o;
  wire _al_u5354_o;
  wire _al_u5357_o;
  wire _al_u5359_o;
  wire _al_u5361_o;
  wire _al_u5363_o;
  wire _al_u5365_o;
  wire _al_u5367_o;
  wire _al_u5369_o;
  wire _al_u5371_o;
  wire _al_u5373_o;
  wire _al_u5375_o;
  wire _al_u5377_o;
  wire _al_u5379_o;
  wire _al_u5381_o;
  wire _al_u5383_o;
  wire _al_u5385_o;
  wire _al_u5387_o;
  wire _al_u5389_o;
  wire _al_u5391_o;
  wire _al_u5393_o;
  wire _al_u5395_o;
  wire _al_u5397_o;
  wire _al_u5399_o;
  wire _al_u5401_o;
  wire _al_u5403_o;
  wire _al_u5405_o;
  wire _al_u5407_o;
  wire _al_u5409_o;
  wire _al_u5411_o;
  wire _al_u5413_o;
  wire _al_u5415_o;
  wire _al_u5417_o;
  wire _al_u5419_o;
  wire _al_u5421_o;
  wire _al_u5423_o;
  wire _al_u5425_o;
  wire _al_u5427_o;
  wire _al_u5429_o;
  wire _al_u5431_o;
  wire _al_u5433_o;
  wire _al_u5435_o;
  wire _al_u5437_o;
  wire _al_u5439_o;
  wire _al_u5441_o;
  wire _al_u5443_o;
  wire _al_u5445_o;
  wire _al_u5447_o;
  wire _al_u5449_o;
  wire _al_u5451_o;
  wire _al_u5453_o;
  wire _al_u5455_o;
  wire _al_u5457_o;
  wire _al_u5459_o;
  wire _al_u5461_o;
  wire _al_u5463_o;
  wire _al_u5465_o;
  wire _al_u5467_o;
  wire _al_u5469_o;
  wire _al_u5471_o;
  wire _al_u5473_o;
  wire _al_u5475_o;
  wire _al_u5477_o;
  wire _al_u5479_o;
  wire _al_u5481_o;
  wire _al_u5483_o;
  wire _al_u5485_o;
  wire _al_u5487_o;
  wire _al_u5489_o;
  wire _al_u5491_o;
  wire _al_u5493_o;
  wire _al_u5495_o;
  wire _al_u5497_o;
  wire _al_u5499_o;
  wire _al_u5501_o;
  wire _al_u5503_o;
  wire _al_u5505_o;
  wire _al_u5507_o;
  wire _al_u5509_o;
  wire _al_u5511_o;
  wire _al_u5513_o;
  wire _al_u5515_o;
  wire _al_u5517_o;
  wire _al_u5519_o;
  wire _al_u5521_o;
  wire _al_u5523_o;
  wire _al_u5525_o;
  wire _al_u5527_o;
  wire _al_u5529_o;
  wire _al_u5531_o;
  wire _al_u5533_o;
  wire _al_u5535_o;
  wire _al_u5537_o;
  wire _al_u5539_o;
  wire _al_u5541_o;
  wire _al_u5543_o;
  wire _al_u5545_o;
  wire _al_u5547_o;
  wire _al_u5549_o;
  wire _al_u5551_o;
  wire _al_u5553_o;
  wire _al_u5555_o;
  wire _al_u5557_o;
  wire _al_u5559_o;
  wire _al_u5561_o;
  wire _al_u5563_o;
  wire _al_u5565_o;
  wire _al_u5567_o;
  wire _al_u5569_o;
  wire _al_u5571_o;
  wire _al_u5573_o;
  wire _al_u5575_o;
  wire _al_u5577_o;
  wire _al_u5579_o;
  wire _al_u5581_o;
  wire _al_u5583_o;
  wire _al_u5585_o;
  wire _al_u5587_o;
  wire _al_u5589_o;
  wire _al_u5591_o;
  wire _al_u5593_o;
  wire _al_u5595_o;
  wire _al_u5597_o;
  wire _al_u5599_o;
  wire _al_u5601_o;
  wire _al_u5604_o;
  wire _al_u5607_o;
  wire _al_u5614_o;
  wire _al_u5662_o;
  wire _al_u5674_o;
  wire _al_u5676_o;
  wire _al_u5677_o;
  wire _al_u5678_o;
  wire _al_u5680_o;
  wire _al_u5681_o;
  wire _al_u5682_o;
  wire _al_u5684_o;
  wire _al_u5685_o;
  wire _al_u5686_o;
  wire _al_u5688_o;
  wire _al_u5689_o;
  wire _al_u5690_o;
  wire _al_u5692_o;
  wire _al_u5693_o;
  wire _al_u5694_o;
  wire _al_u5696_o;
  wire _al_u5697_o;
  wire _al_u5698_o;
  wire _al_u5700_o;
  wire _al_u5701_o;
  wire _al_u5702_o;
  wire _al_u5704_o;
  wire _al_u5705_o;
  wire _al_u5706_o;
  wire _al_u5708_o;
  wire _al_u5709_o;
  wire _al_u5710_o;
  wire _al_u5712_o;
  wire _al_u5713_o;
  wire _al_u5714_o;
  wire _al_u5716_o;
  wire _al_u5717_o;
  wire _al_u5718_o;
  wire _al_u5720_o;
  wire _al_u5721_o;
  wire _al_u5722_o;
  wire _al_u5724_o;
  wire _al_u5725_o;
  wire _al_u5726_o;
  wire _al_u5728_o;
  wire _al_u5729_o;
  wire _al_u5730_o;
  wire _al_u5732_o;
  wire _al_u5733_o;
  wire _al_u5734_o;
  wire _al_u5736_o;
  wire _al_u5737_o;
  wire _al_u5738_o;
  wire _al_u5740_o;
  wire _al_u5741_o;
  wire _al_u5742_o;
  wire _al_u5744_o;
  wire _al_u5745_o;
  wire _al_u5746_o;
  wire _al_u5748_o;
  wire _al_u5749_o;
  wire _al_u5750_o;
  wire _al_u5752_o;
  wire _al_u5753_o;
  wire _al_u5754_o;
  wire _al_u5756_o;
  wire _al_u5757_o;
  wire _al_u5758_o;
  wire _al_u5760_o;
  wire _al_u5761_o;
  wire _al_u5762_o;
  wire _al_u5764_o;
  wire _al_u5765_o;
  wire _al_u5766_o;
  wire _al_u5768_o;
  wire _al_u5769_o;
  wire _al_u5770_o;
  wire _al_u5772_o;
  wire _al_u5773_o;
  wire _al_u5774_o;
  wire _al_u5776_o;
  wire _al_u5777_o;
  wire _al_u5778_o;
  wire _al_u5780_o;
  wire _al_u5781_o;
  wire _al_u5782_o;
  wire _al_u5784_o;
  wire _al_u5785_o;
  wire _al_u5786_o;
  wire _al_u5788_o;
  wire _al_u5789_o;
  wire _al_u5790_o;
  wire _al_u5792_o;
  wire _al_u5793_o;
  wire _al_u5794_o;
  wire _al_u5796_o;
  wire _al_u5797_o;
  wire _al_u5798_o;
  wire _al_u5800_o;
  wire _al_u5801_o;
  wire _al_u5802_o;
  wire _al_u5804_o;
  wire _al_u5805_o;
  wire _al_u5806_o;
  wire _al_u5808_o;
  wire _al_u5809_o;
  wire _al_u5810_o;
  wire _al_u5812_o;
  wire _al_u5813_o;
  wire _al_u5814_o;
  wire _al_u5816_o;
  wire _al_u5817_o;
  wire _al_u5818_o;
  wire _al_u5820_o;
  wire _al_u5821_o;
  wire _al_u5822_o;
  wire _al_u5824_o;
  wire _al_u5825_o;
  wire _al_u5826_o;
  wire _al_u5828_o;
  wire _al_u5829_o;
  wire _al_u5830_o;
  wire _al_u5832_o;
  wire _al_u5833_o;
  wire _al_u5834_o;
  wire _al_u5837_o;
  wire _al_u5839_o;
  wire _al_u5841_o;
  wire _al_u5843_o;
  wire _al_u5845_o;
  wire _al_u5847_o;
  wire _al_u5850_o;
  wire _al_u5851_o;
  wire _al_u5853_o;
  wire _al_u5854_o;
  wire _al_u5856_o;
  wire _al_u5858_o;
  wire _al_u5859_o;
  wire _al_u5860_o;
  wire _al_u5862_o;
  wire _al_u5863_o;
  wire _al_u5865_o;
  wire _al_u5866_o;
  wire _al_u5868_o;
  wire _al_u5869_o;
  wire _al_u5871_o;
  wire _al_u5873_o;
  wire _al_u5874_o;
  wire _al_u5876_o;
  wire _al_u5877_o;
  wire _al_u5879_o;
  wire _al_u5880_o;
  wire _al_u5882_o;
  wire _al_u5883_o;
  wire _al_u5885_o;
  wire _al_u5887_o;
  wire _al_u5888_o;
  wire _al_u5890_o;
  wire _al_u5891_o;
  wire _al_u5893_o;
  wire _al_u5894_o;
  wire _al_u5895_o;
  wire _al_u5896_o;
  wire _al_u5898_o;
  wire _al_u5899_o;
  wire _al_u5900_o;
  wire _al_u5901_o;
  wire _al_u5903_o;
  wire _al_u5904_o;
  wire _al_u5905_o;
  wire _al_u5906_o;
  wire _al_u5908_o;
  wire _al_u5909_o;
  wire _al_u5910_o;
  wire _al_u5911_o;
  wire _al_u5913_o;
  wire _al_u5914_o;
  wire _al_u5915_o;
  wire _al_u5916_o;
  wire _al_u5918_o;
  wire _al_u5919_o;
  wire _al_u5920_o;
  wire _al_u5921_o;
  wire _al_u5923_o;
  wire _al_u5924_o;
  wire _al_u5925_o;
  wire _al_u5926_o;
  wire _al_u5928_o;
  wire _al_u5929_o;
  wire _al_u5930_o;
  wire _al_u5931_o;
  wire _al_u5933_o;
  wire _al_u5934_o;
  wire _al_u5935_o;
  wire _al_u5936_o;
  wire _al_u5938_o;
  wire _al_u5939_o;
  wire _al_u5940_o;
  wire _al_u5941_o;
  wire _al_u5942_o;
  wire _al_u5944_o;
  wire _al_u5945_o;
  wire _al_u5946_o;
  wire _al_u5947_o;
  wire _al_u5948_o;
  wire _al_u5950_o;
  wire _al_u5951_o;
  wire _al_u5952_o;
  wire _al_u5953_o;
  wire _al_u5954_o;
  wire _al_u5956_o;
  wire _al_u5957_o;
  wire _al_u5958_o;
  wire _al_u5959_o;
  wire _al_u5960_o;
  wire _al_u5962_o;
  wire _al_u5963_o;
  wire _al_u5964_o;
  wire _al_u5965_o;
  wire _al_u5966_o;
  wire _al_u5968_o;
  wire _al_u5969_o;
  wire _al_u5970_o;
  wire _al_u5971_o;
  wire _al_u5972_o;
  wire _al_u5974_o;
  wire _al_u5975_o;
  wire _al_u5976_o;
  wire _al_u5977_o;
  wire _al_u5978_o;
  wire _al_u5980_o;
  wire _al_u5981_o;
  wire _al_u5982_o;
  wire _al_u5983_o;
  wire _al_u5984_o;
  wire _al_u5986_o;
  wire _al_u5987_o;
  wire _al_u5988_o;
  wire _al_u5989_o;
  wire _al_u5990_o;
  wire _al_u5992_o;
  wire _al_u6055_o;
  wire _al_u6058_o;
  wire _al_u6059_o;
  wire _al_u6061_o;
  wire _al_u6063_o;
  wire _al_u6064_o;
  wire _al_u6065_o;
  wire _al_u6067_o;
  wire _al_u6068_o;
  wire _al_u6070_o;
  wire _al_u6071_o;
  wire _al_u6073_o;
  wire _al_u6074_o;
  wire _al_u6076_o;
  wire _al_u6077_o;
  wire _al_u6079_o;
  wire _al_u6080_o;
  wire _al_u6082_o;
  wire _al_u6083_o;
  wire _al_u6085_o;
  wire _al_u6086_o;
  wire _al_u6088_o;
  wire _al_u6089_o;
  wire _al_u6091_o;
  wire _al_u6092_o;
  wire _al_u6094_o;
  wire _al_u6095_o;
  wire _al_u6097_o;
  wire _al_u6098_o;
  wire _al_u6100_o;
  wire _al_u6101_o;
  wire _al_u6103_o;
  wire _al_u6104_o;
  wire _al_u6106_o;
  wire _al_u6107_o;
  wire _al_u6109_o;
  wire _al_u6110_o;
  wire _al_u6112_o;
  wire _al_u6113_o;
  wire _al_u6114_o;
  wire _al_u6116_o;
  wire _al_u6117_o;
  wire _al_u6119_o;
  wire _al_u6120_o;
  wire _al_u6122_o;
  wire _al_u6123_o;
  wire _al_u6125_o;
  wire _al_u6126_o;
  wire _al_u6128_o;
  wire _al_u6129_o;
  wire _al_u6131_o;
  wire _al_u6132_o;
  wire _al_u6134_o;
  wire _al_u6135_o;
  wire _al_u6137_o;
  wire _al_u6138_o;
  wire _al_u6140_o;
  wire _al_u6141_o;
  wire _al_u6143_o;
  wire _al_u6144_o;
  wire _al_u6146_o;
  wire _al_u6147_o;
  wire _al_u6149_o;
  wire _al_u6150_o;
  wire _al_u6152_o;
  wire _al_u6153_o;
  wire _al_u6155_o;
  wire _al_u6156_o;
  wire _al_u6158_o;
  wire _al_u6159_o;
  wire _al_u6161_o;
  wire _al_u6162_o;
  wire _al_u6164_o;
  wire _al_u6165_o;
  wire _al_u6167_o;
  wire _al_u6168_o;
  wire _al_u6170_o;
  wire _al_u6171_o;
  wire _al_u6173_o;
  wire _al_u6174_o;
  wire _al_u6176_o;
  wire _al_u6177_o;
  wire _al_u6179_o;
  wire _al_u6180_o;
  wire _al_u6181_o;
  wire _al_u6183_o;
  wire _al_u6184_o;
  wire _al_u6186_o;
  wire _al_u6187_o;
  wire _al_u6189_o;
  wire _al_u6190_o;
  wire _al_u6192_o;
  wire _al_u6193_o;
  wire _al_u6195_o;
  wire _al_u6196_o;
  wire _al_u6198_o;
  wire _al_u6199_o;
  wire _al_u6201_o;
  wire _al_u6202_o;
  wire _al_u6204_o;
  wire _al_u6205_o;
  wire _al_u6207_o;
  wire _al_u6208_o;
  wire _al_u6209_o;
  wire _al_u6211_o;
  wire _al_u6212_o;
  wire _al_u6213_o;
  wire _al_u6215_o;
  wire _al_u6216_o;
  wire _al_u6218_o;
  wire _al_u6219_o;
  wire _al_u6221_o;
  wire _al_u6222_o;
  wire _al_u6224_o;
  wire _al_u6225_o;
  wire _al_u6227_o;
  wire _al_u6228_o;
  wire _al_u6230_o;
  wire _al_u6231_o;
  wire _al_u6233_o;
  wire _al_u6234_o;
  wire _al_u6236_o;
  wire _al_u6237_o;
  wire _al_u6239_o;
  wire _al_u6240_o;
  wire _al_u6243_o;
  wire _al_u6244_o;
  wire _al_u6245_o;
  wire _al_u6246_o;
  wire _al_u6247_o;
  wire _al_u6248_o;
  wire _al_u6249_o;
  wire _al_u6250_o;
  wire _al_u6251_o;
  wire _al_u6254_o;
  wire _al_u6255_o;
  wire _al_u6257_o;
  wire _al_u6258_o;
  wire _al_u6259_o;
  wire _al_u6260_o;
  wire _al_u6261_o;
  wire _al_u6262_o;
  wire _al_u6263_o;
  wire _al_u6264_o;
  wire _al_u6265_o;
  wire _al_u6267_o;
  wire _al_u6268_o;
  wire _al_u6269_o;
  wire _al_u6270_o;
  wire _al_u6271_o;
  wire _al_u6272_o;
  wire _al_u6273_o;
  wire _al_u6274_o;
  wire _al_u6275_o;
  wire _al_u6276_o;
  wire _al_u6277_o;
  wire _al_u6278_o;
  wire _al_u6279_o;
  wire _al_u6280_o;
  wire _al_u6281_o;
  wire _al_u6282_o;
  wire _al_u6283_o;
  wire _al_u6284_o;
  wire _al_u6285_o;
  wire _al_u6286_o;
  wire _al_u6287_o;
  wire _al_u6288_o;
  wire _al_u6289_o;
  wire _al_u6290_o;
  wire _al_u6291_o;
  wire _al_u6292_o;
  wire _al_u6293_o;
  wire _al_u6294_o;
  wire _al_u6295_o;
  wire _al_u6296_o;
  wire _al_u6297_o;
  wire _al_u6298_o;
  wire _al_u6299_o;
  wire _al_u6300_o;
  wire _al_u6301_o;
  wire _al_u6302_o;
  wire _al_u6303_o;
  wire _al_u6304_o;
  wire _al_u6305_o;
  wire _al_u6306_o;
  wire _al_u6307_o;
  wire _al_u6308_o;
  wire _al_u6309_o;
  wire _al_u6311_o;
  wire _al_u6313_o;
  wire _al_u6319_o;
  wire _al_u6320_o;
  wire _al_u6321_o;
  wire _al_u6323_o;
  wire _al_u6326_o;
  wire _al_u6331_o;
  wire _al_u6334_o;
  wire _al_u6336_o;
  wire _al_u6339_o;
  wire _al_u6340_o;
  wire _al_u6341_o;
  wire _al_u6344_o;
  wire _al_u6346_o;
  wire _al_u6348_o;
  wire _al_u6349_o;
  wire _al_u6351_o;
  wire _al_u6352_o;
  wire _al_u6354_o;
  wire _al_u6357_o;
  wire _al_u6359_o;
  wire _al_u6360_o;
  wire _al_u6362_o;
  wire _al_u6363_o;
  wire _al_u6365_o;
  wire _al_u6366_o;
  wire _al_u6367_o;
  wire _al_u6368_o;
  wire _al_u6369_o;
  wire _al_u6370_o;
  wire _al_u6371_o;
  wire _al_u6372_o;
  wire _al_u6373_o;
  wire _al_u6374_o;
  wire _al_u6375_o;
  wire _al_u6376_o;
  wire _al_u6377_o;
  wire _al_u6378_o;
  wire _al_u6379_o;
  wire _al_u6380_o;
  wire _al_u6381_o;
  wire _al_u6382_o;
  wire _al_u6383_o;
  wire _al_u6384_o;
  wire _al_u6385_o;
  wire _al_u6386_o;
  wire _al_u6387_o;
  wire _al_u6388_o;
  wire _al_u6389_o;
  wire _al_u6390_o;
  wire _al_u6391_o;
  wire _al_u6392_o;
  wire _al_u6393_o;
  wire _al_u6394_o;
  wire _al_u6395_o;
  wire _al_u6396_o;
  wire _al_u6397_o;
  wire _al_u6398_o;
  wire _al_u6399_o;
  wire _al_u6400_o;
  wire _al_u6401_o;
  wire _al_u6402_o;
  wire _al_u6403_o;
  wire _al_u6404_o;
  wire _al_u6405_o;
  wire _al_u6406_o;
  wire _al_u6407_o;
  wire _al_u6408_o;
  wire _al_u6409_o;
  wire _al_u6410_o;
  wire _al_u6411_o;
  wire _al_u6412_o;
  wire _al_u6413_o;
  wire _al_u6414_o;
  wire _al_u6415_o;
  wire _al_u6416_o;
  wire _al_u6417_o;
  wire _al_u6418_o;
  wire _al_u6419_o;
  wire _al_u6420_o;
  wire _al_u6423_o;
  wire _al_u6425_o;
  wire _al_u6426_o;
  wire _al_u6436_o;
  wire _al_u6438_o;
  wire _al_u6441_o;
  wire _al_u6443_o;
  wire _al_u6445_o;
  wire _al_u6447_o;
  wire _al_u6449_o;
  wire _al_u6451_o;
  wire _al_u6453_o;
  wire _al_u6455_o;
  wire _al_u6457_o;
  wire _al_u6459_o;
  wire _al_u6461_o;
  wire _al_u6463_o;
  wire _al_u6465_o;
  wire _al_u6467_o;
  wire _al_u6469_o;
  wire _al_u6471_o;
  wire _al_u6473_o;
  wire _al_u6475_o;
  wire _al_u6477_o;
  wire _al_u6479_o;
  wire _al_u6481_o;
  wire _al_u6483_o;
  wire _al_u6485_o;
  wire _al_u6487_o;
  wire _al_u6489_o;
  wire _al_u6491_o;
  wire _al_u6493_o;
  wire _al_u6495_o;
  wire _al_u6497_o;
  wire _al_u6499_o;
  wire _al_u6501_o;
  wire _al_u6503_o;
  wire _al_u6505_o;
  wire _al_u6507_o;
  wire _al_u6509_o;
  wire _al_u6511_o;
  wire _al_u6513_o;
  wire _al_u6515_o;
  wire _al_u6517_o;
  wire _al_u6519_o;
  wire _al_u6521_o;
  wire _al_u6523_o;
  wire _al_u6525_o;
  wire _al_u6527_o;
  wire _al_u6529_o;
  wire _al_u6531_o;
  wire _al_u6533_o;
  wire _al_u6535_o;
  wire _al_u6537_o;
  wire _al_u6539_o;
  wire _al_u6541_o;
  wire _al_u6543_o;
  wire _al_u6545_o;
  wire _al_u6547_o;
  wire _al_u6549_o;
  wire _al_u6551_o;
  wire _al_u6553_o;
  wire _al_u6555_o;
  wire _al_u6557_o;
  wire _al_u6559_o;
  wire _al_u6561_o;
  wire _al_u6563_o;
  wire _al_u6565_o;
  wire _al_u6567_o;
  wire _al_u6570_o;
  wire _al_u6572_o;
  wire _al_u6574_o;
  wire _al_u6576_o;
  wire _al_u6578_o;
  wire _al_u6580_o;
  wire _al_u6582_o;
  wire _al_u6584_o;
  wire _al_u6586_o;
  wire _al_u6588_o;
  wire _al_u6590_o;
  wire _al_u6592_o;
  wire _al_u6594_o;
  wire _al_u6596_o;
  wire _al_u6598_o;
  wire _al_u6600_o;
  wire _al_u6602_o;
  wire _al_u6604_o;
  wire _al_u6606_o;
  wire _al_u6608_o;
  wire _al_u6610_o;
  wire _al_u6612_o;
  wire _al_u6614_o;
  wire _al_u6616_o;
  wire _al_u6618_o;
  wire _al_u6620_o;
  wire _al_u6622_o;
  wire _al_u6624_o;
  wire _al_u6626_o;
  wire _al_u6628_o;
  wire _al_u6630_o;
  wire _al_u6632_o;
  wire _al_u6634_o;
  wire _al_u6636_o;
  wire _al_u6638_o;
  wire _al_u6640_o;
  wire _al_u6642_o;
  wire _al_u6644_o;
  wire _al_u6646_o;
  wire _al_u6648_o;
  wire _al_u6650_o;
  wire _al_u6652_o;
  wire _al_u6654_o;
  wire _al_u6656_o;
  wire _al_u6658_o;
  wire _al_u6660_o;
  wire _al_u6662_o;
  wire _al_u6664_o;
  wire _al_u6666_o;
  wire _al_u6668_o;
  wire _al_u6670_o;
  wire _al_u6672_o;
  wire _al_u6674_o;
  wire _al_u6676_o;
  wire _al_u6678_o;
  wire _al_u6680_o;
  wire _al_u6682_o;
  wire _al_u6684_o;
  wire _al_u6686_o;
  wire _al_u6688_o;
  wire _al_u6690_o;
  wire _al_u6692_o;
  wire _al_u6694_o;
  wire _al_u6696_o;
  wire _al_u6698_o;
  wire _al_u6700_o;
  wire _al_u6702_o;
  wire _al_u6704_o;
  wire _al_u6706_o;
  wire _al_u6708_o;
  wire _al_u6710_o;
  wire _al_u6712_o;
  wire _al_u6714_o;
  wire _al_u6716_o;
  wire _al_u6718_o;
  wire _al_u6720_o;
  wire _al_u6722_o;
  wire _al_u6724_o;
  wire _al_u6725_o;
  wire _al_u6727_o;
  wire _al_u6729_o;
  wire _al_u6731_o;
  wire _al_u6732_o;
  wire _al_u6733_o;
  wire _al_u6734_o;
  wire _al_u6736_o;
  wire _al_u6737_o;
  wire _al_u6738_o;
  wire _al_u6739_o;
  wire _al_u6742_o;
  wire _al_u6743_o;
  wire _al_u6744_o;
  wire _al_u6746_o;
  wire _al_u6747_o;
  wire _al_u6748_o;
  wire _al_u6750_o;
  wire _al_u6751_o;
  wire _al_u6752_o;
  wire _al_u6754_o;
  wire _al_u6755_o;
  wire _al_u6757_o;
  wire _al_u6758_o;
  wire _al_u6760_o;
  wire _al_u6761_o;
  wire _al_u6763_o;
  wire _al_u6764_o;
  wire _al_u6765_o;
  wire _al_u6766_o;
  wire _al_u6768_o;
  wire _al_u6769_o;
  wire _al_u6772_o;
  wire _al_u6775_o;
  wire _al_u6777_o;
  wire _al_u6778_o;
  wire _al_u6780_o;
  wire _al_u6781_o;
  wire _al_u6784_o;
  wire _al_u6785_o;
  wire _al_u6788_o;
  wire _al_u6790_o;
  wire _al_u6791_o;
  wire _al_u6794_o;
  wire _al_u6795_o;
  wire _al_u6796_o;
  wire _al_u6797_o;
  wire _al_u6798_o;
  wire _al_u6799_o;
  wire _al_u6800_o;
  wire _al_u6801_o;
  wire _al_u6803_o;
  wire _al_u6804_o;
  wire _al_u6805_o;
  wire _al_u6806_o;
  wire _al_u6807_o;
  wire _al_u6808_o;
  wire _al_u6809_o;
  wire _al_u6810_o;
  wire _al_u6812_o;
  wire _al_u6813_o;
  wire _al_u6814_o;
  wire _al_u6815_o;
  wire _al_u6816_o;
  wire _al_u6817_o;
  wire _al_u6818_o;
  wire _al_u6819_o;
  wire _al_u6820_o;
  wire _al_u6822_o;
  wire _al_u6823_o;
  wire _al_u6824_o;
  wire _al_u6825_o;
  wire _al_u6826_o;
  wire _al_u6827_o;
  wire _al_u6828_o;
  wire _al_u6829_o;
  wire _al_u6831_o;
  wire _al_u6832_o;
  wire _al_u6833_o;
  wire _al_u6834_o;
  wire _al_u6835_o;
  wire _al_u6836_o;
  wire _al_u6837_o;
  wire _al_u6838_o;
  wire _al_u6839_o;
  wire _al_u6841_o;
  wire _al_u6842_o;
  wire _al_u6843_o;
  wire _al_u6844_o;
  wire _al_u6845_o;
  wire _al_u6846_o;
  wire _al_u6847_o;
  wire _al_u6848_o;
  wire _al_u6850_o;
  wire _al_u6851_o;
  wire _al_u6852_o;
  wire _al_u6853_o;
  wire _al_u6854_o;
  wire _al_u6855_o;
  wire _al_u6856_o;
  wire _al_u6857_o;
  wire _al_u6858_o;
  wire _al_u6860_o;
  wire _al_u6861_o;
  wire _al_u6862_o;
  wire _al_u6863_o;
  wire _al_u6864_o;
  wire _al_u6865_o;
  wire _al_u6866_o;
  wire _al_u6867_o;
  wire _al_u6868_o;
  wire _al_u6870_o;
  wire _al_u6871_o;
  wire _al_u6872_o;
  wire _al_u6873_o;
  wire _al_u6874_o;
  wire _al_u6875_o;
  wire _al_u6876_o;
  wire _al_u6877_o;
  wire _al_u6878_o;
  wire _al_u6880_o;
  wire _al_u6881_o;
  wire _al_u6882_o;
  wire _al_u6883_o;
  wire _al_u6884_o;
  wire _al_u6885_o;
  wire _al_u6886_o;
  wire _al_u6887_o;
  wire _al_u6888_o;
  wire _al_u6890_o;
  wire _al_u6891_o;
  wire _al_u6892_o;
  wire _al_u6893_o;
  wire _al_u6894_o;
  wire _al_u6895_o;
  wire _al_u6896_o;
  wire _al_u6897_o;
  wire _al_u6899_o;
  wire _al_u6900_o;
  wire _al_u6901_o;
  wire _al_u6902_o;
  wire _al_u6903_o;
  wire _al_u6904_o;
  wire _al_u6905_o;
  wire _al_u6906_o;
  wire _al_u6908_o;
  wire _al_u6909_o;
  wire _al_u6910_o;
  wire _al_u6911_o;
  wire _al_u6912_o;
  wire _al_u6913_o;
  wire _al_u6914_o;
  wire _al_u6915_o;
  wire _al_u6917_o;
  wire _al_u6918_o;
  wire _al_u6919_o;
  wire _al_u6920_o;
  wire _al_u6921_o;
  wire _al_u6922_o;
  wire _al_u6923_o;
  wire _al_u6924_o;
  wire _al_u6926_o;
  wire _al_u6927_o;
  wire _al_u6928_o;
  wire _al_u6929_o;
  wire _al_u6930_o;
  wire _al_u6931_o;
  wire _al_u6932_o;
  wire _al_u6933_o;
  wire _al_u6935_o;
  wire _al_u6936_o;
  wire _al_u6938_o;
  wire _al_u6939_o;
  wire _al_u6940_o;
  wire _al_u6942_o;
  wire _al_u6943_o;
  wire _al_u6945_o;
  wire _al_u6947_o;
  wire _al_u6948_o;
  wire _al_u6949_o;
  wire _al_u6950_o;
  wire _al_u6951_o;
  wire _al_u6952_o;
  wire _al_u6953_o;
  wire _al_u6954_o;
  wire _al_u6955_o;
  wire _al_u6957_o;
  wire _al_u6958_o;
  wire _al_u6959_o;
  wire _al_u6960_o;
  wire _al_u6961_o;
  wire _al_u6962_o;
  wire _al_u6963_o;
  wire _al_u6964_o;
  wire _al_u6965_o;
  wire _al_u6967_o;
  wire _al_u6968_o;
  wire _al_u6969_o;
  wire _al_u6970_o;
  wire _al_u6971_o;
  wire _al_u6972_o;
  wire _al_u6973_o;
  wire _al_u6974_o;
  wire _al_u6975_o;
  wire _al_u6977_o;
  wire _al_u6978_o;
  wire _al_u6979_o;
  wire _al_u6980_o;
  wire _al_u6981_o;
  wire _al_u6982_o;
  wire _al_u6983_o;
  wire _al_u6984_o;
  wire _al_u6985_o;
  wire _al_u6987_o;
  wire _al_u6988_o;
  wire _al_u6989_o;
  wire _al_u6990_o;
  wire _al_u6991_o;
  wire _al_u6992_o;
  wire _al_u6993_o;
  wire _al_u6994_o;
  wire _al_u6995_o;
  wire _al_u6997_o;
  wire _al_u6998_o;
  wire _al_u6999_o;
  wire _al_u7000_o;
  wire _al_u7001_o;
  wire _al_u7002_o;
  wire _al_u7003_o;
  wire _al_u7004_o;
  wire _al_u7005_o;
  wire _al_u7006_o;
  wire _al_u7008_o;
  wire _al_u7009_o;
  wire _al_u7010_o;
  wire _al_u7011_o;
  wire _al_u7012_o;
  wire _al_u7013_o;
  wire _al_u7014_o;
  wire _al_u7015_o;
  wire _al_u7016_o;
  wire _al_u7018_o;
  wire _al_u7019_o;
  wire _al_u7020_o;
  wire _al_u7021_o;
  wire _al_u7022_o;
  wire _al_u7023_o;
  wire _al_u7024_o;
  wire _al_u7025_o;
  wire _al_u7026_o;
  wire _al_u7028_o;
  wire _al_u7029_o;
  wire _al_u7030_o;
  wire _al_u7031_o;
  wire _al_u7032_o;
  wire _al_u7033_o;
  wire _al_u7034_o;
  wire _al_u7035_o;
  wire _al_u7036_o;
  wire _al_u7038_o;
  wire _al_u7039_o;
  wire _al_u7040_o;
  wire _al_u7041_o;
  wire _al_u7042_o;
  wire _al_u7043_o;
  wire _al_u7044_o;
  wire _al_u7045_o;
  wire _al_u7046_o;
  wire _al_u7048_o;
  wire _al_u7049_o;
  wire _al_u7050_o;
  wire _al_u7051_o;
  wire _al_u7052_o;
  wire _al_u7053_o;
  wire _al_u7054_o;
  wire _al_u7055_o;
  wire _al_u7056_o;
  wire _al_u7058_o;
  wire _al_u7059_o;
  wire _al_u7060_o;
  wire _al_u7061_o;
  wire _al_u7062_o;
  wire _al_u7063_o;
  wire _al_u7064_o;
  wire _al_u7065_o;
  wire _al_u7066_o;
  wire _al_u7068_o;
  wire _al_u7069_o;
  wire _al_u7070_o;
  wire _al_u7071_o;
  wire _al_u7072_o;
  wire _al_u7073_o;
  wire _al_u7074_o;
  wire _al_u7075_o;
  wire _al_u7076_o;
  wire _al_u7078_o;
  wire _al_u7079_o;
  wire _al_u7080_o;
  wire _al_u7081_o;
  wire _al_u7082_o;
  wire _al_u7083_o;
  wire _al_u7084_o;
  wire _al_u7085_o;
  wire _al_u7086_o;
  wire _al_u7088_o;
  wire _al_u7089_o;
  wire _al_u7090_o;
  wire _al_u7091_o;
  wire _al_u7092_o;
  wire _al_u7093_o;
  wire _al_u7094_o;
  wire _al_u7095_o;
  wire _al_u7096_o;
  wire _al_u7098_o;
  wire _al_u7099_o;
  wire _al_u7100_o;
  wire _al_u7101_o;
  wire _al_u7102_o;
  wire _al_u7103_o;
  wire _al_u7104_o;
  wire _al_u7105_o;
  wire _al_u7106_o;
  wire _al_u7107_o;
  wire _al_u7109_o;
  wire _al_u7110_o;
  wire _al_u7111_o;
  wire _al_u7112_o;
  wire _al_u7113_o;
  wire _al_u7114_o;
  wire _al_u7115_o;
  wire _al_u7116_o;
  wire _al_u7117_o;
  wire _al_u7118_o;
  wire _al_u7120_o;
  wire _al_u7121_o;
  wire _al_u7122_o;
  wire _al_u7123_o;
  wire _al_u7124_o;
  wire _al_u7125_o;
  wire _al_u7126_o;
  wire _al_u7127_o;
  wire _al_u7128_o;
  wire _al_u7129_o;
  wire _al_u7131_o;
  wire _al_u7132_o;
  wire _al_u7133_o;
  wire _al_u7134_o;
  wire _al_u7135_o;
  wire _al_u7136_o;
  wire _al_u7137_o;
  wire _al_u7138_o;
  wire _al_u7139_o;
  wire _al_u7141_o;
  wire _al_u7142_o;
  wire _al_u7145_o;
  wire _al_u7146_o;
  wire _al_u7147_o;
  wire _al_u7149_o;
  wire _al_u7150_o;
  wire _al_u7151_o;
  wire _al_u7152_o;
  wire _al_u7154_o;
  wire _al_u7155_o;
  wire _al_u7156_o;
  wire _al_u7157_o;
  wire _al_u7158_o;
  wire _al_u7159_o;
  wire _al_u7160_o;
  wire _al_u7161_o;
  wire _al_u7162_o;
  wire _al_u7163_o;
  wire _al_u7164_o;
  wire _al_u7165_o;
  wire _al_u7166_o;
  wire _al_u7167_o;
  wire _al_u7168_o;
  wire _al_u7169_o;
  wire _al_u7170_o;
  wire _al_u7171_o;
  wire _al_u7172_o;
  wire _al_u7173_o;
  wire _al_u7174_o;
  wire _al_u7175_o;
  wire _al_u7176_o;
  wire _al_u7177_o;
  wire _al_u7178_o;
  wire _al_u7179_o;
  wire _al_u7180_o;
  wire _al_u7181_o;
  wire _al_u7182_o;
  wire _al_u7183_o;
  wire _al_u7184_o;
  wire _al_u7185_o;
  wire _al_u7186_o;
  wire _al_u7187_o;
  wire _al_u7188_o;
  wire _al_u7190_o;
  wire _al_u7191_o;
  wire _al_u7192_o;
  wire _al_u7193_o;
  wire _al_u7195_o;
  wire _al_u7198_o;
  wire _al_u7199_o;
  wire _al_u7200_o;
  wire _al_u7201_o;
  wire _al_u7202_o;
  wire _al_u7203_o;
  wire _al_u7205_o;
  wire _al_u7206_o;
  wire _al_u7208_o;
  wire _al_u7210_o;
  wire _al_u7211_o;
  wire _al_u7212_o;
  wire _al_u7214_o;
  wire _al_u7215_o;
  wire _al_u7216_o;
  wire _al_u7218_o;
  wire _al_u7219_o;
  wire _al_u7220_o;
  wire _al_u7221_o;
  wire _al_u7222_o;
  wire _al_u7223_o;
  wire _al_u7224_o;
  wire _al_u7226_o;
  wire _al_u7227_o;
  wire _al_u7228_o;
  wire _al_u7229_o;
  wire _al_u7230_o;
  wire _al_u7231_o;
  wire _al_u7232_o;
  wire _al_u7233_o;
  wire _al_u7234_o;
  wire _al_u7235_o;
  wire _al_u7237_o;
  wire _al_u7238_o;
  wire _al_u7239_o;
  wire _al_u7240_o;
  wire _al_u7242_o;
  wire _al_u7243_o;
  wire _al_u7244_o;
  wire _al_u7245_o;
  wire _al_u7246_o;
  wire _al_u7247_o;
  wire _al_u7248_o;
  wire _al_u7249_o;
  wire _al_u7251_o;
  wire _al_u7252_o;
  wire _al_u7253_o;
  wire _al_u7254_o;
  wire _al_u7255_o;
  wire _al_u7256_o;
  wire _al_u7257_o;
  wire _al_u7258_o;
  wire _al_u7259_o;
  wire _al_u7260_o;
  wire _al_u7262_o;
  wire _al_u7263_o;
  wire _al_u7264_o;
  wire _al_u7266_o;
  wire _al_u7267_o;
  wire _al_u7268_o;
  wire _al_u7269_o;
  wire _al_u7270_o;
  wire _al_u7271_o;
  wire _al_u7272_o;
  wire _al_u7274_o;
  wire _al_u7275_o;
  wire _al_u7276_o;
  wire _al_u7277_o;
  wire _al_u7278_o;
  wire _al_u7279_o;
  wire _al_u7280_o;
  wire _al_u7281_o;
  wire _al_u7282_o;
  wire _al_u7283_o;
  wire _al_u7285_o;
  wire _al_u7287_o;
  wire _al_u7288_o;
  wire _al_u7289_o;
  wire _al_u7290_o;
  wire _al_u7291_o;
  wire _al_u7292_o;
  wire _al_u7293_o;
  wire _al_u7294_o;
  wire _al_u7295_o;
  wire _al_u7296_o;
  wire _al_u7330_o;
  wire _al_u7331_o;
  wire _al_u7333_o;
  wire _al_u7335_o;
  wire _al_u7337_o;
  wire _al_u7339_o;
  wire _al_u7340_o;
  wire _al_u7341_o;
  wire _al_u7342_o;
  wire _al_u7343_o;
  wire _al_u7344_o;
  wire _al_u7345_o;
  wire _al_u7346_o;
  wire _al_u7347_o;
  wire _al_u7348_o;
  wire _al_u7349_o;
  wire _al_u7351_o;
  wire _al_u7352_o;
  wire _al_u7353_o;
  wire _al_u7355_o;
  wire _al_u7356_o;
  wire _al_u7358_o;
  wire _al_u7359_o;
  wire _al_u7361_o;
  wire _al_u7362_o;
  wire _al_u7364_o;
  wire _al_u7365_o;
  wire _al_u7367_o;
  wire _al_u7368_o;
  wire _al_u7370_o;
  wire _al_u7371_o;
  wire _al_u7373_o;
  wire _al_u7374_o;
  wire _al_u7376_o;
  wire _al_u7377_o;
  wire _al_u7379_o;
  wire _al_u7380_o;
  wire _al_u7382_o;
  wire _al_u7383_o;
  wire _al_u7385_o;
  wire _al_u7386_o;
  wire _al_u7388_o;
  wire _al_u7389_o;
  wire _al_u7391_o;
  wire _al_u7392_o;
  wire _al_u7394_o;
  wire _al_u7395_o;
  wire _al_u7397_o;
  wire _al_u7398_o;
  wire _al_u7401_o;
  wire _al_u7402_o;
  wire _al_u7403_o;
  wire _al_u7404_o;
  wire _al_u7405_o;
  wire _al_u7406_o;
  wire _al_u7407_o;
  wire _al_u7408_o;
  wire _al_u7409_o;
  wire _al_u7410_o;
  wire _al_u7411_o;
  wire _al_u7413_o;
  wire _al_u7414_o;
  wire _al_u7415_o;
  wire _al_u7416_o;
  wire _al_u7417_o;
  wire _al_u7418_o;
  wire _al_u7419_o;
  wire _al_u7420_o;
  wire _al_u7421_o;
  wire _al_u7422_o;
  wire _al_u7424_o;
  wire _al_u7425_o;
  wire _al_u7426_o;
  wire _al_u7427_o;
  wire _al_u7428_o;
  wire _al_u7429_o;
  wire _al_u7430_o;
  wire _al_u7431_o;
  wire _al_u7432_o;
  wire _al_u7433_o;
  wire _al_u7434_o;
  wire _al_u7436_o;
  wire _al_u7437_o;
  wire _al_u7438_o;
  wire _al_u7439_o;
  wire _al_u7440_o;
  wire _al_u7441_o;
  wire _al_u7442_o;
  wire _al_u7443_o;
  wire _al_u7444_o;
  wire _al_u7445_o;
  wire _al_u7447_o;
  wire _al_u7448_o;
  wire _al_u7449_o;
  wire _al_u7450_o;
  wire _al_u7451_o;
  wire _al_u7452_o;
  wire _al_u7453_o;
  wire _al_u7454_o;
  wire _al_u7455_o;
  wire _al_u7456_o;
  wire _al_u7457_o;
  wire _al_u7459_o;
  wire _al_u7460_o;
  wire _al_u7461_o;
  wire _al_u7462_o;
  wire _al_u7463_o;
  wire _al_u7464_o;
  wire _al_u7465_o;
  wire _al_u7466_o;
  wire _al_u7467_o;
  wire _al_u7468_o;
  wire _al_u7470_o;
  wire _al_u7471_o;
  wire _al_u7472_o;
  wire _al_u7473_o;
  wire _al_u7474_o;
  wire _al_u7475_o;
  wire _al_u7476_o;
  wire _al_u7477_o;
  wire _al_u7478_o;
  wire _al_u7480_o;
  wire _al_u7481_o;
  wire _al_u7482_o;
  wire _al_u7483_o;
  wire _al_u7485_o;
  wire _al_u7486_o;
  wire _al_u7487_o;
  wire _al_u7488_o;
  wire _al_u7489_o;
  wire _al_u7491_o;
  wire _al_u7492_o;
  wire _al_u7493_o;
  wire _al_u7494_o;
  wire _al_u7495_o;
  wire _al_u7497_o;
  wire _al_u7498_o;
  wire _al_u7499_o;
  wire _al_u7500_o;
  wire _al_u7501_o;
  wire _al_u7502_o;
  wire _al_u7503_o;
  wire _al_u7504_o;
  wire _al_u7505_o;
  wire _al_u7506_o;
  wire _al_u7507_o;
  wire _al_u7508_o;
  wire _al_u7510_o;
  wire _al_u7511_o;
  wire _al_u7512_o;
  wire _al_u7514_o;
  wire _al_u7515_o;
  wire _al_u7516_o;
  wire _al_u7518_o;
  wire _al_u7519_o;
  wire _al_u7520_o;
  wire _al_u7522_o;
  wire _al_u7523_o;
  wire _al_u7524_o;
  wire _al_u7526_o;
  wire _al_u7527_o;
  wire _al_u7528_o;
  wire _al_u7530_o;
  wire _al_u7531_o;
  wire _al_u7533_o;
  wire _al_u7534_o;
  wire _al_u7535_o;
  wire _al_u7537_o;
  wire _al_u7538_o;
  wire _al_u7539_o;
  wire _al_u7541_o;
  wire _al_u7542_o;
  wire _al_u7543_o;
  wire _al_u7544_o;
  wire _al_u7545_o;
  wire _al_u7546_o;
  wire _al_u7547_o;
  wire _al_u7548_o;
  wire _al_u7549_o;
  wire _al_u7550_o;
  wire _al_u7551_o;
  wire _al_u7553_o;
  wire _al_u7554_o;
  wire _al_u7555_o;
  wire _al_u7557_o;
  wire _al_u7558_o;
  wire _al_u7559_o;
  wire _al_u7561_o;
  wire _al_u7562_o;
  wire _al_u7563_o;
  wire _al_u7565_o;
  wire _al_u7566_o;
  wire _al_u7567_o;
  wire _al_u7569_o;
  wire _al_u7570_o;
  wire _al_u7571_o;
  wire _al_u7573_o;
  wire _al_u7574_o;
  wire _al_u7575_o;
  wire _al_u7576_o;
  wire _al_u7577_o;
  wire _al_u7578_o;
  wire _al_u7579_o;
  wire _al_u7580_o;
  wire _al_u7581_o;
  wire _al_u7582_o;
  wire _al_u7583_o;
  wire _al_u7585_o;
  wire _al_u7586_o;
  wire _al_u7588_o;
  wire _al_u7589_o;
  wire _al_u7591_o;
  wire _al_u7592_o;
  wire _al_u7594_o;
  wire _al_u7595_o;
  wire _al_u7597_o;
  wire _al_u7598_o;
  wire _al_u7600_o;
  wire _al_u7601_o;
  wire _al_u7602_o;
  wire _al_u7603_o;
  wire _al_u7604_o;
  wire _al_u7605_o;
  wire _al_u7606_o;
  wire _al_u7607_o;
  wire _al_u7608_o;
  wire _al_u7609_o;
  wire _al_u7610_o;
  wire _al_u7612_o;
  wire _al_u7613_o;
  wire _al_u7614_o;
  wire _al_u7615_o;
  wire _al_u7616_o;
  wire _al_u7617_o;
  wire _al_u7618_o;
  wire _al_u7619_o;
  wire _al_u7620_o;
  wire _al_u7621_o;
  wire _al_u7622_o;
  wire _al_u7624_o;
  wire _al_u7625_o;
  wire _al_u7626_o;
  wire _al_u7627_o;
  wire _al_u7628_o;
  wire _al_u7629_o;
  wire _al_u7630_o;
  wire _al_u7631_o;
  wire _al_u7632_o;
  wire _al_u7633_o;
  wire _al_u7634_o;
  wire _al_u7635_o;
  wire _al_u7637_o;
  wire _al_u7638_o;
  wire _al_u7639_o;
  wire _al_u7640_o;
  wire _al_u7641_o;
  wire _al_u7642_o;
  wire _al_u7643_o;
  wire _al_u7644_o;
  wire _al_u7645_o;
  wire _al_u7646_o;
  wire _al_u7647_o;
  wire _al_u7649_o;
  wire _al_u7650_o;
  wire _al_u7652_o;
  wire _al_u7653_o;
  wire _al_u7654_o;
  wire _al_u7655_o;
  wire _al_u7656_o;
  wire _al_u7657_o;
  wire _al_u7658_o;
  wire _al_u7659_o;
  wire _al_u7660_o;
  wire _al_u7661_o;
  wire _al_u7662_o;
  wire _al_u7663_o;
  wire _al_u7665_o;
  wire _al_u7666_o;
  wire _al_u7667_o;
  wire _al_u7668_o;
  wire _al_u7669_o;
  wire _al_u7670_o;
  wire _al_u7671_o;
  wire _al_u7672_o;
  wire _al_u7673_o;
  wire _al_u7674_o;
  wire _al_u7675_o;
  wire _al_u7676_o;
  wire _al_u7678_o;
  wire _al_u7679_o;
  wire _al_u7681_o;
  wire _al_u7682_o;
  wire _al_u7683_o;
  wire _al_u7685_o;
  wire _al_u7686_o;
  wire _al_u7688_o;
  wire _al_u7689_o;
  wire _al_u7691_o;
  wire _al_u7692_o;
  wire _al_u7693_o;
  wire _al_u7694_o;
  wire _al_u7695_o;
  wire _al_u7696_o;
  wire _al_u7697_o;
  wire _al_u7698_o;
  wire _al_u7699_o;
  wire _al_u7700_o;
  wire _al_u7701_o;
  wire _al_u7702_o;
  wire _al_u7704_o;
  wire _al_u7705_o;
  wire _al_u7707_o;
  wire _al_u7708_o;
  wire _al_u7710_o;
  wire _al_u7712_o;
  wire _al_u7713_o;
  wire _al_u7715_o;
  wire _al_u7716_o;
  wire _al_u7717_o;
  wire _al_u7718_o;
  wire _al_u7719_o;
  wire _al_u7720_o;
  wire _al_u7721_o;
  wire _al_u7722_o;
  wire _al_u7723_o;
  wire _al_u7724_o;
  wire _al_u7725_o;
  wire _al_u7726_o;
  wire _al_u7728_o;
  wire _al_u7729_o;
  wire _al_u7730_o;
  wire _al_u7731_o;
  wire _al_u7733_o;
  wire _al_u7734_o;
  wire _al_u7800_o;
  wire _al_u7801_o;
  wire _al_u7803_o;
  wire _al_u7804_o;
  wire _al_u7805_o;
  wire _al_u7806_o;
  wire _al_u7807_o;
  wire _al_u7808_o;
  wire _al_u7809_o;
  wire _al_u7810_o;
  wire _al_u7811_o;
  wire _al_u7812_o;
  wire _al_u7814_o;
  wire _al_u7816_o;
  wire _al_u7817_o;
  wire _al_u7819_o;
  wire _al_u7820_o;
  wire _al_u7822_o;
  wire _al_u7823_o;
  wire _al_u7825_o;
  wire _al_u7826_o;
  wire _al_u7828_o;
  wire _al_u7829_o;
  wire _al_u7831_o;
  wire _al_u7832_o;
  wire _al_u7834_o;
  wire _al_u7836_o;
  wire _al_u7838_o;
  wire _al_u7840_o;
  wire _al_u7842_o;
  wire _al_u7843_o;
  wire _al_u7845_o;
  wire _al_u7846_o;
  wire _al_u7848_o;
  wire _al_u7849_o;
  wire _al_u7851_o;
  wire _al_u7852_o;
  wire _al_u7854_o;
  wire _al_u7855_o;
  wire _al_u7857_o;
  wire _al_u7858_o;
  wire _al_u7859_o;
  wire _al_u7860_o;
  wire _al_u7861_o;
  wire _al_u7862_o;
  wire _al_u7863_o;
  wire _al_u7864_o;
  wire _al_u7865_o;
  wire _al_u7866_o;
  wire _al_u7867_o;
  wire _al_u7868_o;
  wire _al_u7869_o;
  wire _al_u7871_o;
  wire _al_u7873_o;
  wire _al_u7874_o;
  wire _al_u7875_o;
  wire _al_u7876_o;
  wire _al_u7877_o;
  wire _al_u7878_o;
  wire _al_u7879_o;
  wire _al_u7880_o;
  wire _al_u7881_o;
  wire _al_u7882_o;
  wire _al_u7883_o;
  wire _al_u7884_o;
  wire _al_u7885_o;
  wire _al_u7887_o;
  wire _al_u7889_o;
  wire _al_u7891_o;
  wire _al_u7893_o;
  wire _al_u7895_o;
  wire _al_u7897_o;
  wire _al_u7898_o;
  wire _al_u7899_o;
  wire _al_u7900_o;
  wire _al_u7901_o;
  wire _al_u7902_o;
  wire _al_u7905_o;
  wire _al_u7906_o;
  wire _al_u7907_o;
  wire _al_u7908_o;
  wire _al_u7909_o;
  wire _al_u7910_o;
  wire _al_u7911_o;
  wire _al_u7912_o;
  wire _al_u7913_o;
  wire _al_u7915_o;
  wire _al_u7916_o;
  wire _al_u7918_o;
  wire _al_u7919_o;
  wire _al_u7920_o;
  wire _al_u7921_o;
  wire _al_u7922_o;
  wire _al_u7923_o;
  wire _al_u7924_o;
  wire _al_u7925_o;
  wire _al_u7926_o;
  wire _al_u7927_o;
  wire _al_u7928_o;
  wire _al_u7930_o;
  wire _al_u7932_o;
  wire _al_u7933_o;
  wire _al_u7934_o;
  wire _al_u7935_o;
  wire _al_u7936_o;
  wire _al_u7937_o;
  wire _al_u7938_o;
  wire _al_u7939_o;
  wire _al_u7940_o;
  wire _al_u7941_o;
  wire _al_u7942_o;
  wire _al_u7943_o;
  wire _al_u7944_o;
  wire _al_u7945_o;
  wire _al_u7946_o;
  wire _al_u7947_o;
  wire _al_u7948_o;
  wire _al_u7949_o;
  wire _al_u7951_o;
  wire _al_u7953_o;
  wire _al_u7954_o;
  wire _al_u7955_o;
  wire _al_u7956_o;
  wire _al_u7957_o;
  wire _al_u7958_o;
  wire _al_u7959_o;
  wire _al_u7960_o;
  wire _al_u7961_o;
  wire _al_u7963_o;
  wire _al_u7965_o;
  wire _al_u7967_o;
  wire _al_u7968_o;
  wire _al_u7969_o;
  wire _al_u7970_o;
  wire _al_u7971_o;
  wire _al_u7973_o;
  wire _al_u7974_o;
  wire _al_u7975_o;
  wire _al_u7976_o;
  wire _al_u7977_o;
  wire _al_u7978_o;
  wire _al_u7979_o;
  wire _al_u7980_o;
  wire _al_u7981_o;
  wire _al_u7982_o;
  wire _al_u7985_o;
  wire _al_u7986_o;
  wire _al_u7987_o;
  wire _al_u7988_o;
  wire _al_u7990_o;
  wire _al_u7991_o;
  wire _al_u7993_o;
  wire _al_u7994_o;
  wire _al_u7995_o;
  wire _al_u7997_o;
  wire _al_u8000_o;
  wire _al_u8001_o;
  wire _al_u8002_o;
  wire _al_u8005_o;
  wire _al_u8007_o;
  wire _al_u8009_o;
  wire _al_u8011_o;
  wire _al_u8012_o;
  wire _al_u8013_o;
  wire _al_u8014_o;
  wire _al_u8016_o;
  wire _al_u8018_o;
  wire _al_u8019_o;
  wire _al_u8020_o;
  wire _al_u8022_o;
  wire _al_u8025_o;
  wire _al_u8027_o;
  wire _al_u8028_o;
  wire _al_u8029_o;
  wire _al_u8030_o;
  wire _al_u8031_o;
  wire _al_u8032_o;
  wire _al_u8034_o;
  wire _al_u8036_o;
  wire _al_u8037_o;
  wire _al_u8038_o;
  wire _al_u8040_o;
  wire _al_u8041_o;
  wire _al_u8042_o;
  wire _al_u8043_o;
  wire _al_u8045_o;
  wire _al_u8046_o;
  wire _al_u8047_o;
  wire _al_u8048_o;
  wire _al_u8050_o;
  wire _al_u8052_o;
  wire _al_u8053_o;
  wire _al_u8054_o;
  wire _al_u8056_o;
  wire _al_u8057_o;
  wire _al_u8058_o;
  wire _al_u8059_o;
  wire _al_u8061_o;
  wire _al_u8062_o;
  wire _al_u8063_o;
  wire _al_u8064_o;
  wire _al_u8066_o;
  wire _al_u8068_o;
  wire _al_u8069_o;
  wire _al_u8070_o;
  wire _al_u8072_o;
  wire _al_u8074_o;
  wire _al_u8075_o;
  wire _al_u8077_o;
  wire _al_u8078_o;
  wire _al_u8079_o;
  wire _al_u8080_o;
  wire _al_u8082_o;
  wire _al_u8084_o;
  wire _al_u8085_o;
  wire _al_u8086_o;
  wire _al_u8088_o;
  wire _al_u8090_o;
  wire _al_u8091_o;
  wire _al_u8093_o;
  wire _al_u8094_o;
  wire _al_u8095_o;
  wire _al_u8096_o;
  wire _al_u8098_o;
  wire _al_u8100_o;
  wire _al_u8101_o;
  wire _al_u8102_o;
  wire _al_u8104_o;
  wire _al_u8106_o;
  wire _al_u8107_o;
  wire _al_u8109_o;
  wire _al_u8110_o;
  wire _al_u8111_o;
  wire _al_u8112_o;
  wire _al_u8114_o;
  wire _al_u8116_o;
  wire _al_u8117_o;
  wire _al_u8118_o;
  wire _al_u8120_o;
  wire _al_u8122_o;
  wire _al_u8123_o;
  wire _al_u8125_o;
  wire _al_u8126_o;
  wire _al_u8127_o;
  wire _al_u8128_o;
  wire _al_u8129_o;
  wire _al_u8130_o;
  wire _al_u8131_o;
  wire _al_u8132_o;
  wire _al_u8133_o;
  wire _al_u8134_o;
  wire _al_u8136_o;
  wire _al_u8137_o;
  wire _al_u8138_o;
  wire _al_u8140_o;
  wire _al_u8142_o;
  wire _al_u8143_o;
  wire _al_u8145_o;
  wire _al_u8146_o;
  wire _al_u8147_o;
  wire _al_u8148_o;
  wire _al_u8149_o;
  wire _al_u8150_o;
  wire _al_u8151_o;
  wire _al_u8153_o;
  wire _al_u8154_o;
  wire _al_u8155_o;
  wire _al_u8157_o;
  wire _al_u8159_o;
  wire _al_u8160_o;
  wire _al_u8162_o;
  wire _al_u8163_o;
  wire _al_u8164_o;
  wire _al_u8165_o;
  wire _al_u8166_o;
  wire _al_u8167_o;
  wire _al_u8168_o;
  wire _al_u8169_o;
  wire _al_u8171_o;
  wire _al_u8172_o;
  wire _al_u8173_o;
  wire _al_u8175_o;
  wire _al_u8177_o;
  wire _al_u8178_o;
  wire _al_u8180_o;
  wire _al_u8181_o;
  wire _al_u8182_o;
  wire _al_u8183_o;
  wire _al_u8184_o;
  wire _al_u8185_o;
  wire _al_u8186_o;
  wire _al_u8188_o;
  wire _al_u8189_o;
  wire _al_u8190_o;
  wire _al_u8192_o;
  wire _al_u8194_o;
  wire _al_u8195_o;
  wire _al_u8197_o;
  wire _al_u8198_o;
  wire _al_u8199_o;
  wire _al_u8200_o;
  wire _al_u8201_o;
  wire _al_u8202_o;
  wire _al_u8203_o;
  wire _al_u8205_o;
  wire _al_u8206_o;
  wire _al_u8207_o;
  wire _al_u8209_o;
  wire _al_u8211_o;
  wire _al_u8212_o;
  wire _al_u8214_o;
  wire _al_u8215_o;
  wire _al_u8216_o;
  wire _al_u8217_o;
  wire _al_u8218_o;
  wire _al_u8219_o;
  wire _al_u8220_o;
  wire _al_u8222_o;
  wire _al_u8223_o;
  wire _al_u8224_o;
  wire _al_u8226_o;
  wire _al_u8228_o;
  wire _al_u8229_o;
  wire _al_u8231_o;
  wire _al_u8232_o;
  wire _al_u8233_o;
  wire _al_u8234_o;
  wire _al_u8235_o;
  wire _al_u8236_o;
  wire _al_u8237_o;
  wire _al_u8239_o;
  wire _al_u8240_o;
  wire _al_u8241_o;
  wire _al_u8243_o;
  wire _al_u8245_o;
  wire _al_u8246_o;
  wire _al_u8248_o;
  wire _al_u8249_o;
  wire _al_u8250_o;
  wire _al_u8251_o;
  wire _al_u8252_o;
  wire _al_u8253_o;
  wire _al_u8254_o;
  wire _al_u8256_o;
  wire _al_u8257_o;
  wire _al_u8258_o;
  wire _al_u8260_o;
  wire _al_u8262_o;
  wire _al_u8263_o;
  wire _al_u8265_o;
  wire _al_u8266_o;
  wire _al_u8267_o;
  wire _al_u8268_o;
  wire _al_u8269_o;
  wire _al_u8270_o;
  wire _al_u8271_o;
  wire _al_u8272_o;
  wire _al_u8274_o;
  wire _al_u8276_o;
  wire _al_u8277_o;
  wire _al_u8278_o;
  wire _al_u8280_o;
  wire _al_u8282_o;
  wire _al_u8283_o;
  wire _al_u8285_o;
  wire _al_u8286_o;
  wire _al_u8287_o;
  wire _al_u8288_o;
  wire _al_u8289_o;
  wire _al_u8290_o;
  wire _al_u8291_o;
  wire _al_u8293_o;
  wire _al_u8295_o;
  wire _al_u8296_o;
  wire _al_u8297_o;
  wire _al_u8299_o;
  wire _al_u8301_o;
  wire _al_u8302_o;
  wire _al_u8304_o;
  wire _al_u8305_o;
  wire _al_u8306_o;
  wire _al_u8307_o;
  wire _al_u8308_o;
  wire _al_u8309_o;
  wire _al_u8310_o;
  wire _al_u8311_o;
  wire _al_u8313_o;
  wire _al_u8315_o;
  wire _al_u8316_o;
  wire _al_u8317_o;
  wire _al_u8319_o;
  wire _al_u8321_o;
  wire _al_u8322_o;
  wire _al_u8324_o;
  wire _al_u8325_o;
  wire _al_u8326_o;
  wire _al_u8327_o;
  wire _al_u8328_o;
  wire _al_u8329_o;
  wire _al_u8330_o;
  wire _al_u8331_o;
  wire _al_u8333_o;
  wire _al_u8335_o;
  wire _al_u8336_o;
  wire _al_u8337_o;
  wire _al_u8339_o;
  wire _al_u8341_o;
  wire _al_u8342_o;
  wire _al_u8344_o;
  wire _al_u8345_o;
  wire _al_u8346_o;
  wire _al_u8347_o;
  wire _al_u8348_o;
  wire _al_u8349_o;
  wire _al_u8350_o;
  wire _al_u8352_o;
  wire _al_u8354_o;
  wire _al_u8355_o;
  wire _al_u8356_o;
  wire _al_u8358_o;
  wire _al_u8360_o;
  wire _al_u8361_o;
  wire _al_u8363_o;
  wire _al_u8364_o;
  wire _al_u8365_o;
  wire _al_u8366_o;
  wire _al_u8367_o;
  wire _al_u8368_o;
  wire _al_u8369_o;
  wire _al_u8371_o;
  wire _al_u8373_o;
  wire _al_u8374_o;
  wire _al_u8375_o;
  wire _al_u8377_o;
  wire _al_u8379_o;
  wire _al_u8380_o;
  wire _al_u8382_o;
  wire _al_u8383_o;
  wire _al_u8384_o;
  wire _al_u8385_o;
  wire _al_u8386_o;
  wire _al_u8387_o;
  wire _al_u8388_o;
  wire _al_u8390_o;
  wire _al_u8391_o;
  wire _al_u8392_o;
  wire _al_u8393_o;
  wire _al_u8395_o;
  wire _al_u8396_o;
  wire _al_u8397_o;
  wire _al_u8399_o;
  wire _al_u8401_o;
  wire _al_u8402_o;
  wire _al_u8403_o;
  wire _al_u8404_o;
  wire _al_u8405_o;
  wire _al_u8406_o;
  wire _al_u8407_o;
  wire _al_u8409_o;
  wire _al_u8410_o;
  wire _al_u8411_o;
  wire _al_u8412_o;
  wire _al_u8414_o;
  wire _al_u8415_o;
  wire _al_u8416_o;
  wire _al_u8418_o;
  wire _al_u8420_o;
  wire _al_u8421_o;
  wire _al_u8422_o;
  wire _al_u8423_o;
  wire _al_u8424_o;
  wire _al_u8425_o;
  wire _al_u8426_o;
  wire _al_u8427_o;
  wire _al_u8428_o;
  wire _al_u8429_o;
  wire _al_u8430_o;
  wire _al_u8431_o;
  wire _al_u8432_o;
  wire _al_u8433_o;
  wire _al_u8434_o;
  wire _al_u8436_o;
  wire _al_u8437_o;
  wire _al_u8438_o;
  wire _al_u8440_o;
  wire _al_u8442_o;
  wire _al_u8443_o;
  wire _al_u8444_o;
  wire _al_u8445_o;
  wire _al_u8446_o;
  wire _al_u8447_o;
  wire _al_u8448_o;
  wire _al_u8449_o;
  wire _al_u8450_o;
  wire _al_u8451_o;
  wire _al_u8452_o;
  wire _al_u8454_o;
  wire _al_u8455_o;
  wire _al_u8456_o;
  wire _al_u8458_o;
  wire _al_u8459_o;
  wire _al_u8460_o;
  wire _al_u8461_o;
  wire _al_u8463_o;
  wire _al_u8464_o;
  wire _al_u8465_o;
  wire _al_u8466_o;
  wire _al_u8467_o;
  wire _al_u8468_o;
  wire _al_u8469_o;
  wire _al_u8470_o;
  wire _al_u8471_o;
  wire _al_u8472_o;
  wire _al_u8473_o;
  wire _al_u8474_o;
  wire _al_u8476_o;
  wire _al_u8477_o;
  wire _al_u8478_o;
  wire _al_u8480_o;
  wire _al_u8481_o;
  wire _al_u8482_o;
  wire _al_u8483_o;
  wire _al_u8485_o;
  wire _al_u8486_o;
  wire _al_u8487_o;
  wire _al_u8488_o;
  wire _al_u8489_o;
  wire _al_u8490_o;
  wire _al_u8491_o;
  wire _al_u8492_o;
  wire _al_u8493_o;
  wire _al_u8494_o;
  wire _al_u8495_o;
  wire _al_u8496_o;
  wire _al_u8497_o;
  wire _al_u8499_o;
  wire _al_u8500_o;
  wire _al_u8501_o;
  wire _al_u8503_o;
  wire _al_u8505_o;
  wire _al_u8506_o;
  wire _al_u8508_o;
  wire _al_u8509_o;
  wire _al_u8510_o;
  wire _al_u8511_o;
  wire _al_u8512_o;
  wire _al_u8513_o;
  wire _al_u8514_o;
  wire _al_u8515_o;
  wire _al_u8516_o;
  wire _al_u8517_o;
  wire _al_u8518_o;
  wire _al_u8519_o;
  wire _al_u8520_o;
  wire _al_u8521_o;
  wire _al_u8523_o;
  wire _al_u8524_o;
  wire _al_u8525_o;
  wire _al_u8527_o;
  wire _al_u8529_o;
  wire _al_u8530_o;
  wire _al_u8531_o;
  wire _al_u8532_o;
  wire _al_u8533_o;
  wire _al_u8534_o;
  wire _al_u8535_o;
  wire _al_u8536_o;
  wire _al_u8537_o;
  wire _al_u8538_o;
  wire _al_u8539_o;
  wire _al_u8540_o;
  wire _al_u8541_o;
  wire _al_u8542_o;
  wire _al_u8544_o;
  wire _al_u8545_o;
  wire _al_u8546_o;
  wire _al_u8548_o;
  wire _al_u8550_o;
  wire _al_u8551_o;
  wire _al_u8552_o;
  wire _al_u8553_o;
  wire _al_u8554_o;
  wire _al_u8555_o;
  wire _al_u8556_o;
  wire _al_u8557_o;
  wire _al_u8558_o;
  wire _al_u8559_o;
  wire _al_u8561_o;
  wire _al_u8562_o;
  wire _al_u8563_o;
  wire _al_u8565_o;
  wire _al_u8567_o;
  wire _al_u8568_o;
  wire _al_u8570_o;
  wire _al_u8571_o;
  wire _al_u8572_o;
  wire _al_u8573_o;
  wire _al_u8574_o;
  wire _al_u8575_o;
  wire _al_u8576_o;
  wire _al_u8577_o;
  wire _al_u8578_o;
  wire _al_u8579_o;
  wire _al_u8581_o;
  wire _al_u8582_o;
  wire _al_u8583_o;
  wire _al_u8585_o;
  wire _al_u8587_o;
  wire _al_u8588_o;
  wire _al_u8590_o;
  wire _al_u8591_o;
  wire _al_u8592_o;
  wire _al_u8593_o;
  wire _al_u8594_o;
  wire _al_u8595_o;
  wire _al_u8596_o;
  wire _al_u8597_o;
  wire _al_u8598_o;
  wire _al_u8600_o;
  wire _al_u8601_o;
  wire _al_u8602_o;
  wire _al_u8603_o;
  wire _al_u8605_o;
  wire _al_u8606_o;
  wire _al_u8607_o;
  wire _al_u8608_o;
  wire _al_u8609_o;
  wire _al_u8610_o;
  wire _al_u8611_o;
  wire _al_u8612_o;
  wire _al_u8613_o;
  wire _al_u8614_o;
  wire _al_u8615_o;
  wire _al_u8616_o;
  wire _al_u8617_o;
  wire _al_u8618_o;
  wire _al_u8620_o;
  wire _al_u8622_o;
  wire _al_u8624_o;
  wire _al_u8625_o;
  wire _al_u8626_o;
  wire _al_u8627_o;
  wire _al_u8628_o;
  wire _al_u8629_o;
  wire _al_u8630_o;
  wire _al_u8631_o;
  wire _al_u8632_o;
  wire _al_u8633_o;
  wire _al_u8634_o;
  wire _al_u8635_o;
  wire _al_u8636_o;
  wire _al_u8637_o;
  wire _al_u8638_o;
  wire _al_u8640_o;
  wire _al_u8642_o;
  wire _al_u8644_o;
  wire _al_u8645_o;
  wire _al_u8646_o;
  wire _al_u8647_o;
  wire _al_u8648_o;
  wire _al_u8649_o;
  wire _al_u8650_o;
  wire _al_u8651_o;
  wire _al_u8652_o;
  wire _al_u8653_o;
  wire _al_u8654_o;
  wire _al_u8655_o;
  wire _al_u8656_o;
  wire _al_u8657_o;
  wire _al_u8658_o;
  wire _al_u8660_o;
  wire _al_u8662_o;
  wire _al_u8664_o;
  wire _al_u8665_o;
  wire _al_u8666_o;
  wire _al_u8667_o;
  wire _al_u8668_o;
  wire _al_u8669_o;
  wire _al_u8670_o;
  wire _al_u8671_o;
  wire _al_u8672_o;
  wire _al_u8673_o;
  wire _al_u8674_o;
  wire _al_u8675_o;
  wire _al_u8676_o;
  wire _al_u8677_o;
  wire _al_u8679_o;
  wire _al_u8681_o;
  wire _al_u8683_o;
  wire _al_u8684_o;
  wire _al_u8685_o;
  wire _al_u8686_o;
  wire _al_u8687_o;
  wire _al_u8688_o;
  wire _al_u8689_o;
  wire _al_u8690_o;
  wire _al_u8691_o;
  wire _al_u8692_o;
  wire _al_u8693_o;
  wire _al_u8694_o;
  wire _al_u8695_o;
  wire _al_u8696_o;
  wire _al_u8698_o;
  wire _al_u8700_o;
  wire _al_u8702_o;
  wire _al_u8703_o;
  wire _al_u8704_o;
  wire _al_u8705_o;
  wire _al_u8706_o;
  wire _al_u8707_o;
  wire _al_u8708_o;
  wire _al_u8709_o;
  wire _al_u8710_o;
  wire _al_u8711_o;
  wire _al_u8712_o;
  wire _al_u8713_o;
  wire _al_u8714_o;
  wire _al_u8716_o;
  wire _al_u8718_o;
  wire _al_u8720_o;
  wire _al_u8721_o;
  wire _al_u8722_o;
  wire _al_u8723_o;
  wire _al_u8724_o;
  wire _al_u8725_o;
  wire _al_u8726_o;
  wire _al_u8727_o;
  wire _al_u8728_o;
  wire _al_u8729_o;
  wire _al_u8730_o;
  wire _al_u8731_o;
  wire _al_u8732_o;
  wire _al_u8734_o;
  wire _al_u8736_o;
  wire _al_u8738_o;
  wire _al_u8739_o;
  wire _al_u8740_o;
  wire _al_u8741_o;
  wire _al_u8742_o;
  wire _al_u8743_o;
  wire _al_u8744_o;
  wire _al_u8745_o;
  wire _al_u8746_o;
  wire _al_u8747_o;
  wire _al_u8748_o;
  wire _al_u8749_o;
  wire _al_u8750_o;
  wire _al_u8751_o;
  wire _al_u8752_o;
  wire _al_u8753_o;
  wire _al_u8755_o;
  wire _al_u8757_o;
  wire _al_u8759_o;
  wire _al_u8760_o;
  wire _al_u8761_o;
  wire _al_u8762_o;
  wire _al_u8763_o;
  wire _al_u8764_o;
  wire _al_u8765_o;
  wire _al_u8766_o;
  wire _al_u8767_o;
  wire _al_u8768_o;
  wire _al_u8769_o;
  wire _al_u8770_o;
  wire _al_u8771_o;
  wire _al_u8772_o;
  wire _al_u8774_o;
  wire _al_u8776_o;
  wire _al_u8778_o;
  wire _al_u8779_o;
  wire _al_u8780_o;
  wire _al_u8781_o;
  wire _al_u8782_o;
  wire _al_u8783_o;
  wire _al_u8784_o;
  wire _al_u8785_o;
  wire _al_u8786_o;
  wire _al_u8787_o;
  wire _al_u8788_o;
  wire _al_u8789_o;
  wire _al_u8790_o;
  wire _al_u8791_o;
  wire _al_u8793_o;
  wire _al_u8795_o;
  wire _al_u8797_o;
  wire _al_u8798_o;
  wire _al_u8799_o;
  wire _al_u8800_o;
  wire _al_u8801_o;
  wire _al_u8802_o;
  wire _al_u8803_o;
  wire _al_u8804_o;
  wire _al_u8805_o;
  wire _al_u8806_o;
  wire _al_u8807_o;
  wire _al_u8808_o;
  wire _al_u8809_o;
  wire _al_u8810_o;
  wire _al_u8812_o;
  wire _al_u8814_o;
  wire _al_u8816_o;
  wire _al_u8817_o;
  wire _al_u8818_o;
  wire _al_u8819_o;
  wire _al_u8820_o;
  wire _al_u8821_o;
  wire _al_u8822_o;
  wire _al_u8823_o;
  wire _al_u8824_o;
  wire _al_u8825_o;
  wire _al_u8826_o;
  wire _al_u8827_o;
  wire _al_u8828_o;
  wire _al_u8829_o;
  wire _al_u8831_o;
  wire _al_u8833_o;
  wire _al_u8835_o;
  wire _al_u8836_o;
  wire _al_u8837_o;
  wire _al_u8838_o;
  wire _al_u8839_o;
  wire _al_u8840_o;
  wire _al_u8841_o;
  wire _al_u8842_o;
  wire _al_u8843_o;
  wire _al_u8844_o;
  wire _al_u8845_o;
  wire _al_u8846_o;
  wire _al_u8847_o;
  wire _al_u8848_o;
  wire _al_u8850_o;
  wire _al_u8852_o;
  wire _al_u8854_o;
  wire _al_u8855_o;
  wire _al_u8856_o;
  wire _al_u8857_o;
  wire _al_u8858_o;
  wire _al_u8859_o;
  wire _al_u8860_o;
  wire _al_u8861_o;
  wire _al_u8862_o;
  wire _al_u8863_o;
  wire _al_u8864_o;
  wire _al_u8865_o;
  wire _al_u8866_o;
  wire _al_u8868_o;
  wire _al_u8870_o;
  wire _al_u8872_o;
  wire _al_u8873_o;
  wire _al_u8874_o;
  wire _al_u8875_o;
  wire _al_u8876_o;
  wire _al_u8877_o;
  wire _al_u8878_o;
  wire _al_u8879_o;
  wire _al_u8880_o;
  wire _al_u8881_o;
  wire _al_u8882_o;
  wire _al_u8883_o;
  wire _al_u8884_o;
  wire _al_u8886_o;
  wire _al_u8888_o;
  wire _al_u8890_o;
  wire _al_u8891_o;
  wire _al_u8892_o;
  wire _al_u8893_o;
  wire _al_u8894_o;
  wire _al_u8895_o;
  wire _al_u8896_o;
  wire _al_u8897_o;
  wire _al_u8898_o;
  wire _al_u8900_o;
  wire _al_u8902_o;
  wire _al_u8904_o;
  wire _al_u8905_o;
  wire _al_u8906_o;
  wire _al_u8907_o;
  wire _al_u8908_o;
  wire _al_u8909_o;
  wire _al_u8910_o;
  wire _al_u8911_o;
  wire _al_u8912_o;
  wire _al_u8913_o;
  wire _al_u8914_o;
  wire _al_u8915_o;
  wire _al_u8916_o;
  wire _al_u8918_o;
  wire _al_u8920_o;
  wire _al_u8922_o;
  wire _al_u8923_o;
  wire _al_u8924_o;
  wire _al_u8925_o;
  wire _al_u8926_o;
  wire _al_u8927_o;
  wire _al_u8928_o;
  wire _al_u8929_o;
  wire _al_u8930_o;
  wire _al_u8931_o;
  wire _al_u8932_o;
  wire _al_u8933_o;
  wire _al_u8934_o;
  wire _al_u8935_o;
  wire _al_u8937_o;
  wire _al_u8939_o;
  wire _al_u8940_o;
  wire _al_u8941_o;
  wire _al_u8942_o;
  wire _al_u8943_o;
  wire _al_u8944_o;
  wire _al_u8945_o;
  wire _al_u8946_o;
  wire _al_u8947_o;
  wire _al_u8948_o;
  wire _al_u8949_o;
  wire _al_u8950_o;
  wire _al_u8951_o;
  wire _al_u8952_o;
  wire _al_u8953_o;
  wire _al_u8955_o;
  wire _al_u8957_o;
  wire _al_u8959_o;
  wire _al_u8960_o;
  wire _al_u8961_o;
  wire _al_u8962_o;
  wire _al_u8963_o;
  wire _al_u8964_o;
  wire _al_u8965_o;
  wire _al_u8966_o;
  wire _al_u8967_o;
  wire _al_u8968_o;
  wire _al_u8969_o;
  wire _al_u8970_o;
  wire _al_u8971_o;
  wire _al_u8972_o;
  wire _al_u8974_o;
  wire _al_u8976_o;
  wire _al_u8977_o;
  wire _al_u8978_o;
  wire _al_u8979_o;
  wire _al_u8980_o;
  wire _al_u8981_o;
  wire _al_u8982_o;
  wire _al_u8983_o;
  wire _al_u8984_o;
  wire _al_u8985_o;
  wire _al_u8986_o;
  wire _al_u8987_o;
  wire _al_u8988_o;
  wire _al_u8990_o;
  wire _al_u8992_o;
  wire _al_u8994_o;
  wire _al_u8995_o;
  wire _al_u8996_o;
  wire _al_u8997_o;
  wire _al_u8998_o;
  wire _al_u8999_o;
  wire _al_u9000_o;
  wire _al_u9001_o;
  wire _al_u9002_o;
  wire _al_u9003_o;
  wire _al_u9004_o;
  wire _al_u9005_o;
  wire _al_u9006_o;
  wire _al_u9007_o;
  wire _al_u9009_o;
  wire _al_u9011_o;
  wire _al_u9012_o;
  wire _al_u9013_o;
  wire _al_u9014_o;
  wire _al_u9015_o;
  wire _al_u9016_o;
  wire _al_u9017_o;
  wire _al_u9018_o;
  wire _al_u9019_o;
  wire _al_u9020_o;
  wire _al_u9021_o;
  wire _al_u9022_o;
  wire _al_u9023_o;
  wire _al_u9025_o;
  wire _al_u9027_o;
  wire _al_u9029_o;
  wire _al_u9030_o;
  wire _al_u9031_o;
  wire _al_u9032_o;
  wire _al_u9033_o;
  wire _al_u9034_o;
  wire _al_u9035_o;
  wire _al_u9036_o;
  wire _al_u9037_o;
  wire _al_u9038_o;
  wire _al_u9039_o;
  wire _al_u9040_o;
  wire _al_u9041_o;
  wire _al_u9042_o;
  wire _al_u9044_o;
  wire _al_u9046_o;
  wire _al_u9047_o;
  wire _al_u9048_o;
  wire _al_u9049_o;
  wire _al_u9050_o;
  wire _al_u9051_o;
  wire _al_u9052_o;
  wire _al_u9053_o;
  wire _al_u9054_o;
  wire _al_u9055_o;
  wire _al_u9056_o;
  wire _al_u9057_o;
  wire _al_u9058_o;
  wire _al_u9059_o;
  wire _al_u9060_o;
  wire _al_u9062_o;
  wire _al_u9064_o;
  wire _al_u9066_o;
  wire _al_u9067_o;
  wire _al_u9068_o;
  wire _al_u9069_o;
  wire _al_u9070_o;
  wire _al_u9071_o;
  wire _al_u9072_o;
  wire _al_u9073_o;
  wire _al_u9074_o;
  wire _al_u9075_o;
  wire _al_u9076_o;
  wire _al_u9077_o;
  wire _al_u9078_o;
  wire _al_u9079_o;
  wire _al_u9081_o;
  wire _al_u9083_o;
  wire _al_u9084_o;
  wire _al_u9085_o;
  wire _al_u9086_o;
  wire _al_u9087_o;
  wire _al_u9088_o;
  wire _al_u9089_o;
  wire _al_u9090_o;
  wire _al_u9091_o;
  wire _al_u9092_o;
  wire _al_u9093_o;
  wire _al_u9094_o;
  wire _al_u9095_o;
  wire _al_u9096_o;
  wire _al_u9098_o;
  wire _al_u9100_o;
  wire _al_u9102_o;
  wire _al_u9103_o;
  wire _al_u9104_o;
  wire _al_u9105_o;
  wire _al_u9106_o;
  wire _al_u9107_o;
  wire _al_u9108_o;
  wire _al_u9110_o;
  wire _al_u9111_o;
  wire _al_u9112_o;
  wire _al_u9113_o;
  wire _al_u9114_o;
  wire _al_u9117_o;
  wire _al_u9118_o;
  wire _al_u9119_o;
  wire _al_u9121_o;
  wire _al_u9122_o;
  wire _al_u9125_o;
  wire _al_u9126_o;
  wire _al_u9127_o;
  wire _al_u9128_o;
  wire _al_u9129_o;
  wire _al_u9130_o;
  wire _al_u9131_o;
  wire _al_u9133_o;
  wire _al_u9134_o;
  wire _al_u9135_o;
  wire _al_u9137_o;
  wire _al_u9139_o;
  wire _al_u9141_o;
  wire _al_u9142_o;
  wire _al_u9144_o;
  wire _al_u9146_o;
  wire _al_u9147_o;
  wire _al_u9148_o;
  wire _al_u9149_o;
  wire _al_u9151_o;
  wire _al_u9152_o;
  wire _al_u9153_o;
  wire _al_u9154_o;
  wire _al_u9155_o;
  wire _al_u9156_o;
  wire _al_u9158_o;
  wire _al_u9159_o;
  wire _al_u9160_o;
  wire _al_u9161_o;
  wire _al_u9162_o;
  wire _al_u9164_o;
  wire _al_u9165_o;
  wire _al_u9166_o;
  wire _al_u9167_o;
  wire _al_u9168_o;
  wire _al_u9170_o;
  wire _al_u9171_o;
  wire _al_u9173_o;
  wire _al_u9174_o;
  wire _al_u9175_o;
  wire _al_u9176_o;
  wire _al_u9177_o;
  wire _al_u9178_o;
  wire _al_u9179_o;
  wire _al_u9180_o;
  wire _al_u9181_o;
  wire _al_u9182_o;
  wire _al_u9183_o;
  wire _al_u9184_o;
  wire _al_u9186_o;
  wire _al_u9188_o;
  wire _al_u9189_o;
  wire _al_u9190_o;
  wire _al_u9192_o;
  wire _al_u9193_o;
  wire _al_u9195_o;
  wire _al_u9197_o;
  wire _al_u9204_o;
  wire _al_u9205_o;
  wire _al_u9206_o;
  wire _al_u9207_o;
  wire _al_u9208_o;
  wire _al_u9209_o;
  wire _al_u9210_o;
  wire _al_u9211_o;
  wire _al_u9212_o;
  wire _al_u9213_o;
  wire _al_u9214_o;
  wire _al_u9215_o;
  wire _al_u9216_o;
  wire _al_u9217_o;
  wire _al_u9218_o;
  wire _al_u9219_o;
  wire _al_u9220_o;
  wire _al_u9221_o;
  wire _al_u9222_o;
  wire _al_u9223_o;
  wire _al_u9224_o;
  wire _al_u9225_o;
  wire _al_u9226_o;
  wire _al_u9227_o;
  wire _al_u9228_o;
  wire _al_u9229_o;
  wire _al_u9230_o;
  wire _al_u9231_o;
  wire _al_u9232_o;
  wire _al_u9233_o;
  wire _al_u9234_o;
  wire _al_u9235_o;
  wire _al_u9236_o;
  wire _al_u9237_o;
  wire _al_u9238_o;
  wire _al_u9239_o;
  wire _al_u9240_o;
  wire _al_u9241_o;
  wire _al_u9242_o;
  wire _al_u9243_o;
  wire _al_u9244_o;
  wire _al_u9245_o;
  wire _al_u9246_o;
  wire _al_u9247_o;
  wire _al_u9248_o;
  wire _al_u9249_o;
  wire _al_u9250_o;
  wire _al_u9251_o;
  wire _al_u9252_o;
  wire _al_u9253_o;
  wire _al_u9254_o;
  wire _al_u9255_o;
  wire _al_u9256_o;
  wire _al_u9257_o;
  wire _al_u9258_o;
  wire _al_u9259_o;
  wire _al_u9260_o;
  wire _al_u9261_o;
  wire _al_u9262_o;
  wire _al_u9263_o;
  wire _al_u9264_o;
  wire _al_u9265_o;
  wire _al_u9266_o;
  wire _al_u9268_o;
  wire _al_u9270_o;
  wire _al_u9271_o;
  wire _al_u9272_o;
  wire _al_u9273_o;
  wire _al_u9274_o;
  wire _al_u9275_o;
  wire _al_u9276_o;
  wire _al_u9277_o;
  wire _al_u9278_o;
  wire _al_u9279_o;
  wire _al_u9280_o;
  wire _al_u9281_o;
  wire _al_u9283_o;
  wire _al_u9284_o;
  wire _al_u9285_o;
  wire _al_u9286_o;
  wire _al_u9287_o;
  wire _al_u9289_o;
  wire _al_u9290_o;
  wire _al_u9292_o;
  wire _al_u9293_o;
  wire _al_u9294_o;
  wire _al_u9296_o;
  wire _al_u9297_o;
  wire _al_u9298_o;
  wire _al_u9299_o;
  wire _al_u9301_o;
  wire _al_u9302_o;
  wire _al_u9303_o;
  wire _al_u9304_o;
  wire _al_u9306_o;
  wire _al_u9307_o;
  wire _al_u9308_o;
  wire _al_u9309_o;
  wire _al_u9311_o;
  wire _al_u9312_o;
  wire _al_u9313_o;
  wire _al_u9315_o;
  wire _al_u9316_o;
  wire _al_u9317_o;
  wire _al_u9318_o;
  wire _al_u9320_o;
  wire _al_u9321_o;
  wire _al_u9322_o;
  wire _al_u9323_o;
  wire _al_u9325_o;
  wire _al_u9326_o;
  wire _al_u9327_o;
  wire _al_u9328_o;
  wire _al_u9330_o;
  wire _al_u9331_o;
  wire _al_u9332_o;
  wire _al_u9333_o;
  wire _al_u9335_o;
  wire _al_u9336_o;
  wire _al_u9337_o;
  wire _al_u9338_o;
  wire _al_u9340_o;
  wire _al_u9341_o;
  wire _al_u9342_o;
  wire _al_u9343_o;
  wire _al_u9345_o;
  wire _al_u9346_o;
  wire _al_u9347_o;
  wire _al_u9348_o;
  wire _al_u9349_o;
  wire _al_u9350_o;
  wire _al_u9352_o;
  wire _al_u9353_o;
  wire _al_u9354_o;
  wire _al_u9355_o;
  wire _al_u9356_o;
  wire _al_u9357_o;
  wire _al_u9359_o;
  wire _al_u9360_o;
  wire _al_u9361_o;
  wire _al_u9362_o;
  wire _al_u9363_o;
  wire _al_u9364_o;
  wire _al_u9366_o;
  wire _al_u9367_o;
  wire _al_u9368_o;
  wire _al_u9369_o;
  wire _al_u9371_o;
  wire _al_u9372_o;
  wire _al_u9373_o;
  wire _al_u9374_o;
  wire _al_u9375_o;
  wire _al_u9376_o;
  wire _al_u9378_o;
  wire _al_u9379_o;
  wire _al_u9380_o;
  wire _al_u9381_o;
  wire _al_u9382_o;
  wire _al_u9383_o;
  wire _al_u9385_o;
  wire _al_u9386_o;
  wire _al_u9387_o;
  wire _al_u9388_o;
  wire _al_u9389_o;
  wire _al_u9390_o;
  wire _al_u9392_o;
  wire _al_u9393_o;
  wire _al_u9394_o;
  wire _al_u9395_o;
  wire _al_u9396_o;
  wire _al_u9397_o;
  wire _al_u9399_o;
  wire _al_u9400_o;
  wire _al_u9401_o;
  wire _al_u9402_o;
  wire _al_u9404_o;
  wire _al_u9405_o;
  wire _al_u9406_o;
  wire _al_u9407_o;
  wire _al_u9408_o;
  wire _al_u9409_o;
  wire _al_u9411_o;
  wire _al_u9412_o;
  wire _al_u9413_o;
  wire _al_u9414_o;
  wire _al_u9415_o;
  wire _al_u9416_o;
  wire _al_u9418_o;
  wire _al_u9419_o;
  wire _al_u9420_o;
  wire _al_u9421_o;
  wire _al_u9422_o;
  wire _al_u9423_o;
  wire _al_u9425_o;
  wire _al_u9426_o;
  wire _al_u9427_o;
  wire _al_u9428_o;
  wire _al_u9430_o;
  wire _al_u9431_o;
  wire _al_u9432_o;
  wire _al_u9433_o;
  wire _al_u9434_o;
  wire _al_u9435_o;
  wire _al_u9437_o;
  wire _al_u9438_o;
  wire _al_u9439_o;
  wire _al_u9440_o;
  wire _al_u9441_o;
  wire _al_u9442_o;
  wire _al_u9444_o;
  wire _al_u9445_o;
  wire _al_u9446_o;
  wire _al_u9447_o;
  wire _al_u9449_o;
  wire _al_u9450_o;
  wire _al_u9451_o;
  wire _al_u9452_o;
  wire _al_u9453_o;
  wire _al_u9454_o;
  wire _al_u9456_o;
  wire _al_u9457_o;
  wire _al_u9458_o;
  wire _al_u9459_o;
  wire _al_u9461_o;
  wire _al_u9462_o;
  wire _al_u9463_o;
  wire _al_u9464_o;
  wire _al_u9465_o;
  wire _al_u9466_o;
  wire _al_u9468_o;
  wire _al_u9469_o;
  wire _al_u9470_o;
  wire _al_u9471_o;
  wire _al_u9473_o;
  wire _al_u9474_o;
  wire _al_u9475_o;
  wire _al_u9476_o;
  wire _al_u9477_o;
  wire _al_u9478_o;
  wire _al_u9480_o;
  wire _al_u9481_o;
  wire _al_u9482_o;
  wire _al_u9483_o;
  wire _al_u9484_o;
  wire _al_u9485_o;
  wire _al_u9487_o;
  wire _al_u9488_o;
  wire _al_u9489_o;
  wire _al_u9490_o;
  wire _al_u9491_o;
  wire _al_u9492_o;
  wire _al_u9494_o;
  wire _al_u9495_o;
  wire _al_u9496_o;
  wire _al_u9497_o;
  wire _al_u9499_o;
  wire _al_u9500_o;
  wire _al_u9501_o;
  wire _al_u9502_o;
  wire _al_u9503_o;
  wire _al_u9504_o;
  wire _al_u9506_o;
  wire _al_u9507_o;
  wire _al_u9508_o;
  wire _al_u9509_o;
  wire _al_u9510_o;
  wire _al_u9511_o;
  wire _al_u9513_o;
  wire _al_u9514_o;
  wire _al_u9515_o;
  wire _al_u9516_o;
  wire _al_u9518_o;
  wire _al_u9519_o;
  wire _al_u9520_o;
  wire _al_u9521_o;
  wire _al_u9522_o;
  wire _al_u9523_o;
  wire _al_u9525_o;
  wire _al_u9526_o;
  wire _al_u9527_o;
  wire _al_u9528_o;
  wire _al_u9530_o;
  wire _al_u9531_o;
  wire _al_u9532_o;
  wire _al_u9533_o;
  wire _al_u9534_o;
  wire _al_u9535_o;
  wire _al_u9537_o;
  wire _al_u9538_o;
  wire _al_u9539_o;
  wire _al_u9540_o;
  wire _al_u9541_o;
  wire _al_u9542_o;
  wire _al_u9544_o;
  wire _al_u9545_o;
  wire _al_u9546_o;
  wire _al_u9547_o;
  wire _al_u9548_o;
  wire _al_u9549_o;
  wire _al_u9551_o;
  wire _al_u9552_o;
  wire _al_u9553_o;
  wire _al_u9554_o;
  wire _al_u9555_o;
  wire _al_u9556_o;
  wire _al_u9558_o;
  wire _al_u9559_o;
  wire _al_u9560_o;
  wire _al_u9561_o;
  wire _al_u9562_o;
  wire _al_u9563_o;
  wire _al_u9565_o;
  wire _al_u9566_o;
  wire _al_u9567_o;
  wire _al_u9568_o;
  wire _al_u9569_o;
  wire _al_u9570_o;
  wire _al_u9572_o;
  wire _al_u9573_o;
  wire _al_u9574_o;
  wire _al_u9575_o;
  wire _al_u9576_o;
  wire _al_u9577_o;
  wire _al_u9579_o;
  wire _al_u9580_o;
  wire _al_u9581_o;
  wire _al_u9582_o;
  wire _al_u9583_o;
  wire _al_u9584_o;
  wire _al_u9586_o;
  wire _al_u9587_o;
  wire _al_u9588_o;
  wire _al_u9589_o;
  wire _al_u9591_o;
  wire _al_u9592_o;
  wire _al_u9593_o;
  wire _al_u9594_o;
  wire _al_u9595_o;
  wire _al_u9596_o;
  wire _al_u9598_o;
  wire _al_u9599_o;
  wire _al_u9600_o;
  wire _al_u9601_o;
  wire _al_u9602_o;
  wire _al_u9603_o;
  wire _al_u9605_o;
  wire _al_u9606_o;
  wire _al_u9607_o;
  wire _al_u9608_o;
  wire _al_u9609_o;
  wire _al_u9610_o;
  wire _al_u9612_o;
  wire _al_u9613_o;
  wire _al_u9614_o;
  wire _al_u9615_o;
  wire _al_u9616_o;
  wire _al_u9617_o;
  wire _al_u9619_o;
  wire _al_u9620_o;
  wire _al_u9621_o;
  wire _al_u9622_o;
  wire _al_u9624_o;
  wire _al_u9625_o;
  wire _al_u9626_o;
  wire _al_u9627_o;
  wire _al_u9628_o;
  wire _al_u9629_o;
  wire _al_u9631_o;
  wire _al_u9632_o;
  wire _al_u9633_o;
  wire _al_u9634_o;
  wire _al_u9635_o;
  wire _al_u9636_o;
  wire _al_u9638_o;
  wire _al_u9639_o;
  wire _al_u9640_o;
  wire _al_u9641_o;
  wire _al_u9642_o;
  wire _al_u9643_o;
  wire _al_u9645_o;
  wire _al_u9646_o;
  wire _al_u9647_o;
  wire _al_u9648_o;
  wire _al_u9650_o;
  wire _al_u9651_o;
  wire _al_u9652_o;
  wire _al_u9653_o;
  wire _al_u9654_o;
  wire _al_u9655_o;
  wire _al_u9657_o;
  wire _al_u9658_o;
  wire _al_u9659_o;
  wire _al_u9660_o;
  wire _al_u9661_o;
  wire _al_u9662_o;
  wire _al_u9664_o;
  wire _al_u9665_o;
  wire _al_u9666_o;
  wire _al_u9667_o;
  wire _al_u9669_o;
  wire _al_u9670_o;
  wire _al_u9671_o;
  wire _al_u9672_o;
  wire _al_u9673_o;
  wire _al_u9674_o;
  wire _al_u9676_o;
  wire _al_u9677_o;
  wire _al_u9678_o;
  wire _al_u9679_o;
  wire _al_u9680_o;
  wire _al_u9681_o;
  wire _al_u9682_o;
  wire _al_u9683_o;
  wire _al_u9685_o;
  wire _al_u9686_o;
  wire _al_u9687_o;
  wire _al_u9688_o;
  wire _al_u9689_o;
  wire _al_u9690_o;
  wire _al_u9691_o;
  wire _al_u9692_o;
  wire _al_u9693_o;
  wire _al_u9695_o;
  wire _al_u9696_o;
  wire _al_u9697_o;
  wire _al_u9698_o;
  wire _al_u9699_o;
  wire _al_u9700_o;
  wire _al_u9701_o;
  wire _al_u9702_o;
  wire _al_u9704_o;
  wire _al_u9705_o;
  wire _al_u9706_o;
  wire _al_u9707_o;
  wire _al_u9708_o;
  wire _al_u9709_o;
  wire _al_u9710_o;
  wire _al_u9711_o;
  wire _al_u9712_o;
  wire _al_u9713_o;
  wire amo;  // ../../RTL/CPU/prv464_top.v(138)
  wire and_clr;  // ../../RTL/CPU/prv464_top.v(129)
  wire \biu/bus_unit/add0/c0 ;
  wire \biu/bus_unit/add0/c1 ;
  wire \biu/bus_unit/add0/c2 ;
  wire \biu/bus_unit/add0/c3 ;
  wire \biu/bus_unit/add0/c4 ;
  wire \biu/bus_unit/add0/c5 ;
  wire \biu/bus_unit/add0/c6 ;
  wire \biu/bus_unit/add0/c7 ;
  wire \biu/bus_unit/add0/c8 ;
  wire \biu/bus_unit/add1/c0 ;
  wire \biu/bus_unit/add1/c1 ;
  wire \biu/bus_unit/add1/c10 ;
  wire \biu/bus_unit/add1/c11 ;
  wire \biu/bus_unit/add1/c12 ;
  wire \biu/bus_unit/add1/c13 ;
  wire \biu/bus_unit/add1/c14 ;
  wire \biu/bus_unit/add1/c15 ;
  wire \biu/bus_unit/add1/c16 ;
  wire \biu/bus_unit/add1/c17 ;
  wire \biu/bus_unit/add1/c18 ;
  wire \biu/bus_unit/add1/c19 ;
  wire \biu/bus_unit/add1/c2 ;
  wire \biu/bus_unit/add1/c20 ;
  wire \biu/bus_unit/add1/c21 ;
  wire \biu/bus_unit/add1/c22 ;
  wire \biu/bus_unit/add1/c23 ;
  wire \biu/bus_unit/add1/c24 ;
  wire \biu/bus_unit/add1/c25 ;
  wire \biu/bus_unit/add1/c26 ;
  wire \biu/bus_unit/add1/c27 ;
  wire \biu/bus_unit/add1/c28 ;
  wire \biu/bus_unit/add1/c29 ;
  wire \biu/bus_unit/add1/c3 ;
  wire \biu/bus_unit/add1/c30 ;
  wire \biu/bus_unit/add1/c31 ;
  wire \biu/bus_unit/add1/c32 ;
  wire \biu/bus_unit/add1/c33 ;
  wire \biu/bus_unit/add1/c34 ;
  wire \biu/bus_unit/add1/c35 ;
  wire \biu/bus_unit/add1/c36 ;
  wire \biu/bus_unit/add1/c37 ;
  wire \biu/bus_unit/add1/c38 ;
  wire \biu/bus_unit/add1/c39 ;
  wire \biu/bus_unit/add1/c4 ;
  wire \biu/bus_unit/add1/c40 ;
  wire \biu/bus_unit/add1/c41 ;
  wire \biu/bus_unit/add1/c42 ;
  wire \biu/bus_unit/add1/c43 ;
  wire \biu/bus_unit/add1/c44 ;
  wire \biu/bus_unit/add1/c45 ;
  wire \biu/bus_unit/add1/c46 ;
  wire \biu/bus_unit/add1/c47 ;
  wire \biu/bus_unit/add1/c48 ;
  wire \biu/bus_unit/add1/c49 ;
  wire \biu/bus_unit/add1/c5 ;
  wire \biu/bus_unit/add1/c50 ;
  wire \biu/bus_unit/add1/c51 ;
  wire \biu/bus_unit/add1/c52 ;
  wire \biu/bus_unit/add1/c53 ;
  wire \biu/bus_unit/add1/c54 ;
  wire \biu/bus_unit/add1/c55 ;
  wire \biu/bus_unit/add1/c56 ;
  wire \biu/bus_unit/add1/c57 ;
  wire \biu/bus_unit/add1/c58 ;
  wire \biu/bus_unit/add1/c59 ;
  wire \biu/bus_unit/add1/c6 ;
  wire \biu/bus_unit/add1/c60 ;
  wire \biu/bus_unit/add1/c7 ;
  wire \biu/bus_unit/add1/c8 ;
  wire \biu/bus_unit/add1/c9 ;
  wire \biu/bus_unit/mmu/mux10_b0_sel_is_2_o ;
  wire \biu/bus_unit/mmu/mux18_b3_sel_is_2_o ;
  wire \biu/bus_unit/mmu/mux20_b0_sel_is_3_o ;
  wire \biu/bus_unit/mmu/mux24_b0_sel_is_1_o ;
  wire \biu/bus_unit/mmu/mux34_b0_sel_is_3_o ;
  wire \biu/bus_unit/mmu/n12_lutinv ;
  wire \biu/bus_unit/mmu/n19_lutinv ;
  wire \biu/bus_unit/mmu/n2 ;
  wire \biu/bus_unit/mmu/n31_lutinv ;
  wire \biu/bus_unit/mmu/n37_lutinv ;
  wire \biu/bus_unit/mmu/n45_lutinv ;
  wire \biu/bus_unit/mmu/n58 ;
  wire \biu/bus_unit/mmu/n7_lutinv ;
  wire \biu/bus_unit/mmu/n8_lutinv ;
  wire \biu/bus_unit/mux10_b3_sel_is_0_o ;
  wire \biu/bus_unit/mux11_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux15_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux17_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux1_b1_sel_is_0_o ;
  wire \biu/bus_unit/n15_lutinv ;
  wire \biu/bus_unit/n37 ;
  wire \biu/bus_unit/n39[0]_d ;
  wire \biu/bus_unit/n39[0]_en ;
  wire \biu/bus_unit/n39[1]_d ;
  wire \biu/bus_unit/n39[2]_d ;
  wire \biu/bus_unit/n39[3]_d ;
  wire \biu/bus_unit/n39[4]_d ;
  wire \biu/bus_unit/n39[5]_d ;
  wire \biu/bus_unit/n39[6]_d ;
  wire \biu/bus_unit/n39[7]_d ;
  wire \biu/bus_unit/n39[8]_d ;
  wire \biu/bus_unit/n45_lutinv ;
  wire \biu/bus_unit/sub0/c0 ;
  wire \biu/bus_unit/sub0/c1 ;
  wire \biu/bus_unit/sub0/c2 ;
  wire \biu/bus_unit/sub0/c3 ;
  wire \biu/bus_unit/sub0/c4 ;
  wire \biu/bus_unit/sub0/c5 ;
  wire \biu/bus_unit/sub0/c6 ;
  wire \biu/bus_unit/sub0/c7 ;
  wire \biu/bus_unit/sub0/c8 ;
  wire \biu/cache/n1 ;
  wire \biu/cache/n11 ;
  wire \biu/cache/n13 ;
  wire \biu/cache/n15 ;
  wire \biu/cache/n17 ;
  wire \biu/cache/n19 ;
  wire \biu/cache/n21 ;
  wire \biu/cache/n23 ;
  wire \biu/cache/n25 ;
  wire \biu/cache/n27 ;
  wire \biu/cache/n29 ;
  wire \biu/cache/n3 ;
  wire \biu/cache/n31 ;
  wire \biu/cache/n5 ;
  wire \biu/cache/n7 ;
  wire \biu/cache/n9 ;
  wire \biu/cache_ctrl_logic/add0/c0 ;
  wire \biu/cache_ctrl_logic/add0/c1 ;
  wire \biu/cache_ctrl_logic/add0/c10 ;
  wire \biu/cache_ctrl_logic/add0/c11 ;
  wire \biu/cache_ctrl_logic/add0/c12 ;
  wire \biu/cache_ctrl_logic/add0/c13 ;
  wire \biu/cache_ctrl_logic/add0/c14 ;
  wire \biu/cache_ctrl_logic/add0/c15 ;
  wire \biu/cache_ctrl_logic/add0/c16 ;
  wire \biu/cache_ctrl_logic/add0/c17 ;
  wire \biu/cache_ctrl_logic/add0/c18 ;
  wire \biu/cache_ctrl_logic/add0/c19 ;
  wire \biu/cache_ctrl_logic/add0/c2 ;
  wire \biu/cache_ctrl_logic/add0/c20 ;
  wire \biu/cache_ctrl_logic/add0/c21 ;
  wire \biu/cache_ctrl_logic/add0/c22 ;
  wire \biu/cache_ctrl_logic/add0/c23 ;
  wire \biu/cache_ctrl_logic/add0/c24 ;
  wire \biu/cache_ctrl_logic/add0/c25 ;
  wire \biu/cache_ctrl_logic/add0/c26 ;
  wire \biu/cache_ctrl_logic/add0/c27 ;
  wire \biu/cache_ctrl_logic/add0/c28 ;
  wire \biu/cache_ctrl_logic/add0/c29 ;
  wire \biu/cache_ctrl_logic/add0/c3 ;
  wire \biu/cache_ctrl_logic/add0/c30 ;
  wire \biu/cache_ctrl_logic/add0/c31 ;
  wire \biu/cache_ctrl_logic/add0/c32 ;
  wire \biu/cache_ctrl_logic/add0/c33 ;
  wire \biu/cache_ctrl_logic/add0/c34 ;
  wire \biu/cache_ctrl_logic/add0/c35 ;
  wire \biu/cache_ctrl_logic/add0/c36 ;
  wire \biu/cache_ctrl_logic/add0/c37 ;
  wire \biu/cache_ctrl_logic/add0/c38 ;
  wire \biu/cache_ctrl_logic/add0/c39 ;
  wire \biu/cache_ctrl_logic/add0/c4 ;
  wire \biu/cache_ctrl_logic/add0/c40 ;
  wire \biu/cache_ctrl_logic/add0/c41 ;
  wire \biu/cache_ctrl_logic/add0/c42 ;
  wire \biu/cache_ctrl_logic/add0/c43 ;
  wire \biu/cache_ctrl_logic/add0/c44 ;
  wire \biu/cache_ctrl_logic/add0/c45 ;
  wire \biu/cache_ctrl_logic/add0/c46 ;
  wire \biu/cache_ctrl_logic/add0/c47 ;
  wire \biu/cache_ctrl_logic/add0/c48 ;
  wire \biu/cache_ctrl_logic/add0/c49 ;
  wire \biu/cache_ctrl_logic/add0/c5 ;
  wire \biu/cache_ctrl_logic/add0/c50 ;
  wire \biu/cache_ctrl_logic/add0/c51 ;
  wire \biu/cache_ctrl_logic/add0/c52 ;
  wire \biu/cache_ctrl_logic/add0/c53 ;
  wire \biu/cache_ctrl_logic/add0/c54 ;
  wire \biu/cache_ctrl_logic/add0/c55 ;
  wire \biu/cache_ctrl_logic/add0/c56 ;
  wire \biu/cache_ctrl_logic/add0/c57 ;
  wire \biu/cache_ctrl_logic/add0/c58 ;
  wire \biu/cache_ctrl_logic/add0/c59 ;
  wire \biu/cache_ctrl_logic/add0/c6 ;
  wire \biu/cache_ctrl_logic/add0/c60 ;
  wire \biu/cache_ctrl_logic/add0/c61 ;
  wire \biu/cache_ctrl_logic/add0/c62 ;
  wire \biu/cache_ctrl_logic/add0/c63 ;
  wire \biu/cache_ctrl_logic/add0/c7 ;
  wire \biu/cache_ctrl_logic/add0/c8 ;
  wire \biu/cache_ctrl_logic/add0/c9 ;
  wire \biu/cache_ctrl_logic/add1/c0 ;
  wire \biu/cache_ctrl_logic/add1/c1 ;
  wire \biu/cache_ctrl_logic/add1/c10 ;
  wire \biu/cache_ctrl_logic/add1/c11 ;
  wire \biu/cache_ctrl_logic/add1/c12 ;
  wire \biu/cache_ctrl_logic/add1/c13 ;
  wire \biu/cache_ctrl_logic/add1/c14 ;
  wire \biu/cache_ctrl_logic/add1/c15 ;
  wire \biu/cache_ctrl_logic/add1/c16 ;
  wire \biu/cache_ctrl_logic/add1/c17 ;
  wire \biu/cache_ctrl_logic/add1/c18 ;
  wire \biu/cache_ctrl_logic/add1/c19 ;
  wire \biu/cache_ctrl_logic/add1/c2 ;
  wire \biu/cache_ctrl_logic/add1/c20 ;
  wire \biu/cache_ctrl_logic/add1/c21 ;
  wire \biu/cache_ctrl_logic/add1/c22 ;
  wire \biu/cache_ctrl_logic/add1/c23 ;
  wire \biu/cache_ctrl_logic/add1/c24 ;
  wire \biu/cache_ctrl_logic/add1/c25 ;
  wire \biu/cache_ctrl_logic/add1/c26 ;
  wire \biu/cache_ctrl_logic/add1/c27 ;
  wire \biu/cache_ctrl_logic/add1/c28 ;
  wire \biu/cache_ctrl_logic/add1/c29 ;
  wire \biu/cache_ctrl_logic/add1/c3 ;
  wire \biu/cache_ctrl_logic/add1/c30 ;
  wire \biu/cache_ctrl_logic/add1/c31 ;
  wire \biu/cache_ctrl_logic/add1/c32 ;
  wire \biu/cache_ctrl_logic/add1/c33 ;
  wire \biu/cache_ctrl_logic/add1/c34 ;
  wire \biu/cache_ctrl_logic/add1/c35 ;
  wire \biu/cache_ctrl_logic/add1/c36 ;
  wire \biu/cache_ctrl_logic/add1/c37 ;
  wire \biu/cache_ctrl_logic/add1/c38 ;
  wire \biu/cache_ctrl_logic/add1/c39 ;
  wire \biu/cache_ctrl_logic/add1/c4 ;
  wire \biu/cache_ctrl_logic/add1/c40 ;
  wire \biu/cache_ctrl_logic/add1/c41 ;
  wire \biu/cache_ctrl_logic/add1/c42 ;
  wire \biu/cache_ctrl_logic/add1/c43 ;
  wire \biu/cache_ctrl_logic/add1/c44 ;
  wire \biu/cache_ctrl_logic/add1/c45 ;
  wire \biu/cache_ctrl_logic/add1/c46 ;
  wire \biu/cache_ctrl_logic/add1/c47 ;
  wire \biu/cache_ctrl_logic/add1/c48 ;
  wire \biu/cache_ctrl_logic/add1/c49 ;
  wire \biu/cache_ctrl_logic/add1/c5 ;
  wire \biu/cache_ctrl_logic/add1/c50 ;
  wire \biu/cache_ctrl_logic/add1/c51 ;
  wire \biu/cache_ctrl_logic/add1/c52 ;
  wire \biu/cache_ctrl_logic/add1/c53 ;
  wire \biu/cache_ctrl_logic/add1/c54 ;
  wire \biu/cache_ctrl_logic/add1/c55 ;
  wire \biu/cache_ctrl_logic/add1/c56 ;
  wire \biu/cache_ctrl_logic/add1/c57 ;
  wire \biu/cache_ctrl_logic/add1/c58 ;
  wire \biu/cache_ctrl_logic/add1/c59 ;
  wire \biu/cache_ctrl_logic/add1/c6 ;
  wire \biu/cache_ctrl_logic/add1/c60 ;
  wire \biu/cache_ctrl_logic/add1/c61 ;
  wire \biu/cache_ctrl_logic/add1/c62 ;
  wire \biu/cache_ctrl_logic/add1/c63 ;
  wire \biu/cache_ctrl_logic/add1/c7 ;
  wire \biu/cache_ctrl_logic/add1/c8 ;
  wire \biu/cache_ctrl_logic/add1/c9 ;
  wire \biu/cache_ctrl_logic/add2/c0 ;
  wire \biu/cache_ctrl_logic/add2/c1 ;
  wire \biu/cache_ctrl_logic/add2/c10 ;
  wire \biu/cache_ctrl_logic/add2/c11 ;
  wire \biu/cache_ctrl_logic/add2/c12 ;
  wire \biu/cache_ctrl_logic/add2/c13 ;
  wire \biu/cache_ctrl_logic/add2/c14 ;
  wire \biu/cache_ctrl_logic/add2/c15 ;
  wire \biu/cache_ctrl_logic/add2/c16 ;
  wire \biu/cache_ctrl_logic/add2/c17 ;
  wire \biu/cache_ctrl_logic/add2/c18 ;
  wire \biu/cache_ctrl_logic/add2/c19 ;
  wire \biu/cache_ctrl_logic/add2/c2 ;
  wire \biu/cache_ctrl_logic/add2/c20 ;
  wire \biu/cache_ctrl_logic/add2/c21 ;
  wire \biu/cache_ctrl_logic/add2/c22 ;
  wire \biu/cache_ctrl_logic/add2/c23 ;
  wire \biu/cache_ctrl_logic/add2/c24 ;
  wire \biu/cache_ctrl_logic/add2/c25 ;
  wire \biu/cache_ctrl_logic/add2/c26 ;
  wire \biu/cache_ctrl_logic/add2/c27 ;
  wire \biu/cache_ctrl_logic/add2/c28 ;
  wire \biu/cache_ctrl_logic/add2/c29 ;
  wire \biu/cache_ctrl_logic/add2/c3 ;
  wire \biu/cache_ctrl_logic/add2/c30 ;
  wire \biu/cache_ctrl_logic/add2/c31 ;
  wire \biu/cache_ctrl_logic/add2/c32 ;
  wire \biu/cache_ctrl_logic/add2/c33 ;
  wire \biu/cache_ctrl_logic/add2/c34 ;
  wire \biu/cache_ctrl_logic/add2/c35 ;
  wire \biu/cache_ctrl_logic/add2/c36 ;
  wire \biu/cache_ctrl_logic/add2/c37 ;
  wire \biu/cache_ctrl_logic/add2/c38 ;
  wire \biu/cache_ctrl_logic/add2/c39 ;
  wire \biu/cache_ctrl_logic/add2/c4 ;
  wire \biu/cache_ctrl_logic/add2/c40 ;
  wire \biu/cache_ctrl_logic/add2/c41 ;
  wire \biu/cache_ctrl_logic/add2/c42 ;
  wire \biu/cache_ctrl_logic/add2/c43 ;
  wire \biu/cache_ctrl_logic/add2/c44 ;
  wire \biu/cache_ctrl_logic/add2/c45 ;
  wire \biu/cache_ctrl_logic/add2/c46 ;
  wire \biu/cache_ctrl_logic/add2/c47 ;
  wire \biu/cache_ctrl_logic/add2/c48 ;
  wire \biu/cache_ctrl_logic/add2/c49 ;
  wire \biu/cache_ctrl_logic/add2/c5 ;
  wire \biu/cache_ctrl_logic/add2/c50 ;
  wire \biu/cache_ctrl_logic/add2/c51 ;
  wire \biu/cache_ctrl_logic/add2/c52 ;
  wire \biu/cache_ctrl_logic/add2/c53 ;
  wire \biu/cache_ctrl_logic/add2/c54 ;
  wire \biu/cache_ctrl_logic/add2/c55 ;
  wire \biu/cache_ctrl_logic/add2/c56 ;
  wire \biu/cache_ctrl_logic/add2/c57 ;
  wire \biu/cache_ctrl_logic/add2/c58 ;
  wire \biu/cache_ctrl_logic/add2/c59 ;
  wire \biu/cache_ctrl_logic/add2/c6 ;
  wire \biu/cache_ctrl_logic/add2/c60 ;
  wire \biu/cache_ctrl_logic/add2/c61 ;
  wire \biu/cache_ctrl_logic/add2/c62 ;
  wire \biu/cache_ctrl_logic/add2/c63 ;
  wire \biu/cache_ctrl_logic/add2/c7 ;
  wire \biu/cache_ctrl_logic/add2/c8 ;
  wire \biu/cache_ctrl_logic/add2/c9 ;
  wire \biu/cache_ctrl_logic/eq1/xor_i0[4]_i1[4]_o_lutinv ;
  wire \biu/cache_ctrl_logic/ex_l1i_hit ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(155)
  wire \biu/cache_ctrl_logic/l1d_value ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(138)
  wire \biu/cache_ctrl_logic/l1d_value_d ;
  wire \biu/cache_ctrl_logic/l1d_wr_sel_lutinv ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(435)
  wire \biu/cache_ctrl_logic/l1i_value ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(137)
  wire \biu/cache_ctrl_logic/l1i_value_d ;
  wire \biu/cache_ctrl_logic/mux31_b4_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux44_b4_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/n127[4]_d ;
  wire \biu/cache_ctrl_logic/n131[1]_d ;
  wire \biu/cache_ctrl_logic/n132[0]_d ;
  wire \biu/cache_ctrl_logic/n135 ;
  wire \biu/cache_ctrl_logic/n140 ;
  wire \biu/cache_ctrl_logic/n149 ;
  wire \biu/cache_ctrl_logic/n17 ;
  wire \biu/cache_ctrl_logic/n172_lutinv ;
  wire \biu/cache_ctrl_logic/n173_lutinv ;
  wire \biu/cache_ctrl_logic/n174_lutinv ;
  wire \biu/cache_ctrl_logic/n176_lutinv ;
  wire \biu/cache_ctrl_logic/n204_lutinv ;
  wire \biu/cache_ctrl_logic/n26_lutinv ;
  wire \biu/cache_ctrl_logic/n30 ;
  wire \biu/cache_ctrl_logic/n34 ;
  wire \biu/cache_ctrl_logic/n36 ;
  wire \biu/cache_ctrl_logic/n40 ;
  wire \biu/cache_ctrl_logic/n42 ;
  wire \biu/cache_ctrl_logic/n55_lutinv ;
  wire \biu/cache_ctrl_logic/n75_lutinv ;
  wire \biu/cache_ctrl_logic/n97_lutinv ;
  wire \biu/cache_ctrl_logic/u128_sel_is_0_o ;
  wire \biu/cache_write_lutinv ;  // ../../RTL/CPU/BIU/biu.v(115)
  wire \biu/cacheable ;  // ../../RTL/CPU/BIU/biu.v(113)
  wire \biu/l1i_write_lutinv ;  // ../../RTL/CPU/BIU/biu.v(83)
  wire cache_flush;  // ../../RTL/CPU/prv464_top.v(139)
  wire cache_reset;  // ../../RTL/CPU/prv464_top.v(140)
  wire clk_pad;  // ../../RTL/CPU/prv464_top.v(19)
  wire \cu_ru/add0_2/c0 ;
  wire \cu_ru/add0_2/c1 ;
  wire \cu_ru/add0_2/c10 ;
  wire \cu_ru/add0_2/c11 ;
  wire \cu_ru/add0_2/c12 ;
  wire \cu_ru/add0_2/c13 ;
  wire \cu_ru/add0_2/c14 ;
  wire \cu_ru/add0_2/c15 ;
  wire \cu_ru/add0_2/c16 ;
  wire \cu_ru/add0_2/c17 ;
  wire \cu_ru/add0_2/c18 ;
  wire \cu_ru/add0_2/c19 ;
  wire \cu_ru/add0_2/c2 ;
  wire \cu_ru/add0_2/c20 ;
  wire \cu_ru/add0_2/c21 ;
  wire \cu_ru/add0_2/c22 ;
  wire \cu_ru/add0_2/c23 ;
  wire \cu_ru/add0_2/c24 ;
  wire \cu_ru/add0_2/c25 ;
  wire \cu_ru/add0_2/c26 ;
  wire \cu_ru/add0_2/c27 ;
  wire \cu_ru/add0_2/c28 ;
  wire \cu_ru/add0_2/c29 ;
  wire \cu_ru/add0_2/c3 ;
  wire \cu_ru/add0_2/c30 ;
  wire \cu_ru/add0_2/c31 ;
  wire \cu_ru/add0_2/c32 ;
  wire \cu_ru/add0_2/c33 ;
  wire \cu_ru/add0_2/c34 ;
  wire \cu_ru/add0_2/c35 ;
  wire \cu_ru/add0_2/c36 ;
  wire \cu_ru/add0_2/c37 ;
  wire \cu_ru/add0_2/c38 ;
  wire \cu_ru/add0_2/c39 ;
  wire \cu_ru/add0_2/c4 ;
  wire \cu_ru/add0_2/c40 ;
  wire \cu_ru/add0_2/c41 ;
  wire \cu_ru/add0_2/c42 ;
  wire \cu_ru/add0_2/c43 ;
  wire \cu_ru/add0_2/c44 ;
  wire \cu_ru/add0_2/c45 ;
  wire \cu_ru/add0_2/c46 ;
  wire \cu_ru/add0_2/c47 ;
  wire \cu_ru/add0_2/c48 ;
  wire \cu_ru/add0_2/c49 ;
  wire \cu_ru/add0_2/c5 ;
  wire \cu_ru/add0_2/c50 ;
  wire \cu_ru/add0_2/c51 ;
  wire \cu_ru/add0_2/c52 ;
  wire \cu_ru/add0_2/c53 ;
  wire \cu_ru/add0_2/c54 ;
  wire \cu_ru/add0_2/c55 ;
  wire \cu_ru/add0_2/c56 ;
  wire \cu_ru/add0_2/c57 ;
  wire \cu_ru/add0_2/c58 ;
  wire \cu_ru/add0_2/c59 ;
  wire \cu_ru/add0_2/c6 ;
  wire \cu_ru/add0_2/c60 ;
  wire \cu_ru/add0_2/c7 ;
  wire \cu_ru/add0_2/c8 ;
  wire \cu_ru/add0_2/c9 ;
  wire \cu_ru/add0_2_co ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_000 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_001 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_002 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_003 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_004 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_005 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_006 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_007 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_008 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_009 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_010 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_011 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_012 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_013 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_014 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_015 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_016 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_017 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_018 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_019 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_020 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_021 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_022 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_023 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_024 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_025 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_026 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_027 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_028 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_029 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_030 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_031 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_032 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_033 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_034 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_035 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_036 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_037 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_038 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_039 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_040 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_041 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_042 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_043 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_044 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_045 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_046 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_047 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_048 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_049 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_050 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_051 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_052 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_053 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_054 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_055 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_056 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_057 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_058 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_059 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_060 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_061 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_062 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i0_063 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_000 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_001 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_002 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_003 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_004 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_005 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_006 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_007 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_008 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_009 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_010 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_011 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_012 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_013 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_014 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_015 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_016 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_017 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_018 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_019 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_020 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_021 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_022 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_023 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_024 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_025 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_026 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_027 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_028 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_029 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_030 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_031 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_032 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_033 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_034 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_035 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_036 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_037 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_038 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_039 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_040 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_041 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_042 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_043 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_044 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_045 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_046 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_047 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_048 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_049 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_050 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_051 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_052 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_053 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_054 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_055 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_056 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_057 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_058 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_059 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_060 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_061 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_062 ;
  wire \cu_ru/al_ram_gpr_al_u0_do_i1_063 ;
  wire \cu_ru/al_ram_gpr_do_i0_000 ;
  wire \cu_ru/al_ram_gpr_do_i0_001 ;
  wire \cu_ru/al_ram_gpr_do_i0_002 ;
  wire \cu_ru/al_ram_gpr_do_i0_003 ;
  wire \cu_ru/al_ram_gpr_do_i0_004 ;
  wire \cu_ru/al_ram_gpr_do_i0_005 ;
  wire \cu_ru/al_ram_gpr_do_i0_006 ;
  wire \cu_ru/al_ram_gpr_do_i0_007 ;
  wire \cu_ru/al_ram_gpr_do_i0_008 ;
  wire \cu_ru/al_ram_gpr_do_i0_009 ;
  wire \cu_ru/al_ram_gpr_do_i0_010 ;
  wire \cu_ru/al_ram_gpr_do_i0_011 ;
  wire \cu_ru/al_ram_gpr_do_i0_012 ;
  wire \cu_ru/al_ram_gpr_do_i0_013 ;
  wire \cu_ru/al_ram_gpr_do_i0_014 ;
  wire \cu_ru/al_ram_gpr_do_i0_015 ;
  wire \cu_ru/al_ram_gpr_do_i0_016 ;
  wire \cu_ru/al_ram_gpr_do_i0_017 ;
  wire \cu_ru/al_ram_gpr_do_i0_018 ;
  wire \cu_ru/al_ram_gpr_do_i0_019 ;
  wire \cu_ru/al_ram_gpr_do_i0_020 ;
  wire \cu_ru/al_ram_gpr_do_i0_021 ;
  wire \cu_ru/al_ram_gpr_do_i0_022 ;
  wire \cu_ru/al_ram_gpr_do_i0_023 ;
  wire \cu_ru/al_ram_gpr_do_i0_024 ;
  wire \cu_ru/al_ram_gpr_do_i0_025 ;
  wire \cu_ru/al_ram_gpr_do_i0_026 ;
  wire \cu_ru/al_ram_gpr_do_i0_027 ;
  wire \cu_ru/al_ram_gpr_do_i0_028 ;
  wire \cu_ru/al_ram_gpr_do_i0_029 ;
  wire \cu_ru/al_ram_gpr_do_i0_030 ;
  wire \cu_ru/al_ram_gpr_do_i0_031 ;
  wire \cu_ru/al_ram_gpr_do_i0_032 ;
  wire \cu_ru/al_ram_gpr_do_i0_033 ;
  wire \cu_ru/al_ram_gpr_do_i0_034 ;
  wire \cu_ru/al_ram_gpr_do_i0_035 ;
  wire \cu_ru/al_ram_gpr_do_i0_036 ;
  wire \cu_ru/al_ram_gpr_do_i0_037 ;
  wire \cu_ru/al_ram_gpr_do_i0_038 ;
  wire \cu_ru/al_ram_gpr_do_i0_039 ;
  wire \cu_ru/al_ram_gpr_do_i0_040 ;
  wire \cu_ru/al_ram_gpr_do_i0_041 ;
  wire \cu_ru/al_ram_gpr_do_i0_042 ;
  wire \cu_ru/al_ram_gpr_do_i0_043 ;
  wire \cu_ru/al_ram_gpr_do_i0_044 ;
  wire \cu_ru/al_ram_gpr_do_i0_045 ;
  wire \cu_ru/al_ram_gpr_do_i0_046 ;
  wire \cu_ru/al_ram_gpr_do_i0_047 ;
  wire \cu_ru/al_ram_gpr_do_i0_048 ;
  wire \cu_ru/al_ram_gpr_do_i0_049 ;
  wire \cu_ru/al_ram_gpr_do_i0_050 ;
  wire \cu_ru/al_ram_gpr_do_i0_051 ;
  wire \cu_ru/al_ram_gpr_do_i0_052 ;
  wire \cu_ru/al_ram_gpr_do_i0_053 ;
  wire \cu_ru/al_ram_gpr_do_i0_054 ;
  wire \cu_ru/al_ram_gpr_do_i0_055 ;
  wire \cu_ru/al_ram_gpr_do_i0_056 ;
  wire \cu_ru/al_ram_gpr_do_i0_057 ;
  wire \cu_ru/al_ram_gpr_do_i0_058 ;
  wire \cu_ru/al_ram_gpr_do_i0_059 ;
  wire \cu_ru/al_ram_gpr_do_i0_060 ;
  wire \cu_ru/al_ram_gpr_do_i0_061 ;
  wire \cu_ru/al_ram_gpr_do_i0_062 ;
  wire \cu_ru/al_ram_gpr_do_i0_063 ;
  wire \cu_ru/al_ram_gpr_do_i1_000 ;
  wire \cu_ru/al_ram_gpr_do_i1_001 ;
  wire \cu_ru/al_ram_gpr_do_i1_002 ;
  wire \cu_ru/al_ram_gpr_do_i1_003 ;
  wire \cu_ru/al_ram_gpr_do_i1_004 ;
  wire \cu_ru/al_ram_gpr_do_i1_005 ;
  wire \cu_ru/al_ram_gpr_do_i1_006 ;
  wire \cu_ru/al_ram_gpr_do_i1_007 ;
  wire \cu_ru/al_ram_gpr_do_i1_008 ;
  wire \cu_ru/al_ram_gpr_do_i1_009 ;
  wire \cu_ru/al_ram_gpr_do_i1_010 ;
  wire \cu_ru/al_ram_gpr_do_i1_011 ;
  wire \cu_ru/al_ram_gpr_do_i1_012 ;
  wire \cu_ru/al_ram_gpr_do_i1_013 ;
  wire \cu_ru/al_ram_gpr_do_i1_014 ;
  wire \cu_ru/al_ram_gpr_do_i1_015 ;
  wire \cu_ru/al_ram_gpr_do_i1_016 ;
  wire \cu_ru/al_ram_gpr_do_i1_017 ;
  wire \cu_ru/al_ram_gpr_do_i1_018 ;
  wire \cu_ru/al_ram_gpr_do_i1_019 ;
  wire \cu_ru/al_ram_gpr_do_i1_020 ;
  wire \cu_ru/al_ram_gpr_do_i1_021 ;
  wire \cu_ru/al_ram_gpr_do_i1_022 ;
  wire \cu_ru/al_ram_gpr_do_i1_023 ;
  wire \cu_ru/al_ram_gpr_do_i1_024 ;
  wire \cu_ru/al_ram_gpr_do_i1_025 ;
  wire \cu_ru/al_ram_gpr_do_i1_026 ;
  wire \cu_ru/al_ram_gpr_do_i1_027 ;
  wire \cu_ru/al_ram_gpr_do_i1_028 ;
  wire \cu_ru/al_ram_gpr_do_i1_029 ;
  wire \cu_ru/al_ram_gpr_do_i1_030 ;
  wire \cu_ru/al_ram_gpr_do_i1_031 ;
  wire \cu_ru/al_ram_gpr_do_i1_032 ;
  wire \cu_ru/al_ram_gpr_do_i1_033 ;
  wire \cu_ru/al_ram_gpr_do_i1_034 ;
  wire \cu_ru/al_ram_gpr_do_i1_035 ;
  wire \cu_ru/al_ram_gpr_do_i1_036 ;
  wire \cu_ru/al_ram_gpr_do_i1_037 ;
  wire \cu_ru/al_ram_gpr_do_i1_038 ;
  wire \cu_ru/al_ram_gpr_do_i1_039 ;
  wire \cu_ru/al_ram_gpr_do_i1_040 ;
  wire \cu_ru/al_ram_gpr_do_i1_041 ;
  wire \cu_ru/al_ram_gpr_do_i1_042 ;
  wire \cu_ru/al_ram_gpr_do_i1_043 ;
  wire \cu_ru/al_ram_gpr_do_i1_044 ;
  wire \cu_ru/al_ram_gpr_do_i1_045 ;
  wire \cu_ru/al_ram_gpr_do_i1_046 ;
  wire \cu_ru/al_ram_gpr_do_i1_047 ;
  wire \cu_ru/al_ram_gpr_do_i1_048 ;
  wire \cu_ru/al_ram_gpr_do_i1_049 ;
  wire \cu_ru/al_ram_gpr_do_i1_050 ;
  wire \cu_ru/al_ram_gpr_do_i1_051 ;
  wire \cu_ru/al_ram_gpr_do_i1_052 ;
  wire \cu_ru/al_ram_gpr_do_i1_053 ;
  wire \cu_ru/al_ram_gpr_do_i1_054 ;
  wire \cu_ru/al_ram_gpr_do_i1_055 ;
  wire \cu_ru/al_ram_gpr_do_i1_056 ;
  wire \cu_ru/al_ram_gpr_do_i1_057 ;
  wire \cu_ru/al_ram_gpr_do_i1_058 ;
  wire \cu_ru/al_ram_gpr_do_i1_059 ;
  wire \cu_ru/al_ram_gpr_do_i1_060 ;
  wire \cu_ru/al_ram_gpr_do_i1_061 ;
  wire \cu_ru/al_ram_gpr_do_i1_062 ;
  wire \cu_ru/al_ram_gpr_do_i1_063 ;
  wire \cu_ru/csr_satp/n0 ;
  wire \cu_ru/m_cycle_event/add0/c0 ;
  wire \cu_ru/m_cycle_event/add0/c1 ;
  wire \cu_ru/m_cycle_event/add0/c10 ;
  wire \cu_ru/m_cycle_event/add0/c11 ;
  wire \cu_ru/m_cycle_event/add0/c12 ;
  wire \cu_ru/m_cycle_event/add0/c13 ;
  wire \cu_ru/m_cycle_event/add0/c14 ;
  wire \cu_ru/m_cycle_event/add0/c15 ;
  wire \cu_ru/m_cycle_event/add0/c16 ;
  wire \cu_ru/m_cycle_event/add0/c17 ;
  wire \cu_ru/m_cycle_event/add0/c18 ;
  wire \cu_ru/m_cycle_event/add0/c19 ;
  wire \cu_ru/m_cycle_event/add0/c2 ;
  wire \cu_ru/m_cycle_event/add0/c20 ;
  wire \cu_ru/m_cycle_event/add0/c21 ;
  wire \cu_ru/m_cycle_event/add0/c22 ;
  wire \cu_ru/m_cycle_event/add0/c23 ;
  wire \cu_ru/m_cycle_event/add0/c24 ;
  wire \cu_ru/m_cycle_event/add0/c25 ;
  wire \cu_ru/m_cycle_event/add0/c26 ;
  wire \cu_ru/m_cycle_event/add0/c27 ;
  wire \cu_ru/m_cycle_event/add0/c28 ;
  wire \cu_ru/m_cycle_event/add0/c29 ;
  wire \cu_ru/m_cycle_event/add0/c3 ;
  wire \cu_ru/m_cycle_event/add0/c30 ;
  wire \cu_ru/m_cycle_event/add0/c31 ;
  wire \cu_ru/m_cycle_event/add0/c32 ;
  wire \cu_ru/m_cycle_event/add0/c33 ;
  wire \cu_ru/m_cycle_event/add0/c34 ;
  wire \cu_ru/m_cycle_event/add0/c35 ;
  wire \cu_ru/m_cycle_event/add0/c36 ;
  wire \cu_ru/m_cycle_event/add0/c37 ;
  wire \cu_ru/m_cycle_event/add0/c38 ;
  wire \cu_ru/m_cycle_event/add0/c39 ;
  wire \cu_ru/m_cycle_event/add0/c4 ;
  wire \cu_ru/m_cycle_event/add0/c40 ;
  wire \cu_ru/m_cycle_event/add0/c41 ;
  wire \cu_ru/m_cycle_event/add0/c42 ;
  wire \cu_ru/m_cycle_event/add0/c43 ;
  wire \cu_ru/m_cycle_event/add0/c44 ;
  wire \cu_ru/m_cycle_event/add0/c45 ;
  wire \cu_ru/m_cycle_event/add0/c46 ;
  wire \cu_ru/m_cycle_event/add0/c47 ;
  wire \cu_ru/m_cycle_event/add0/c48 ;
  wire \cu_ru/m_cycle_event/add0/c49 ;
  wire \cu_ru/m_cycle_event/add0/c5 ;
  wire \cu_ru/m_cycle_event/add0/c50 ;
  wire \cu_ru/m_cycle_event/add0/c51 ;
  wire \cu_ru/m_cycle_event/add0/c52 ;
  wire \cu_ru/m_cycle_event/add0/c53 ;
  wire \cu_ru/m_cycle_event/add0/c54 ;
  wire \cu_ru/m_cycle_event/add0/c55 ;
  wire \cu_ru/m_cycle_event/add0/c56 ;
  wire \cu_ru/m_cycle_event/add0/c57 ;
  wire \cu_ru/m_cycle_event/add0/c58 ;
  wire \cu_ru/m_cycle_event/add0/c59 ;
  wire \cu_ru/m_cycle_event/add0/c6 ;
  wire \cu_ru/m_cycle_event/add0/c60 ;
  wire \cu_ru/m_cycle_event/add0/c61 ;
  wire \cu_ru/m_cycle_event/add0/c62 ;
  wire \cu_ru/m_cycle_event/add0/c63 ;
  wire \cu_ru/m_cycle_event/add0/c7 ;
  wire \cu_ru/m_cycle_event/add0/c8 ;
  wire \cu_ru/m_cycle_event/add0/c9 ;
  wire \cu_ru/m_cycle_event/add1/c0 ;
  wire \cu_ru/m_cycle_event/add1/c1 ;
  wire \cu_ru/m_cycle_event/add1/c10 ;
  wire \cu_ru/m_cycle_event/add1/c11 ;
  wire \cu_ru/m_cycle_event/add1/c12 ;
  wire \cu_ru/m_cycle_event/add1/c13 ;
  wire \cu_ru/m_cycle_event/add1/c14 ;
  wire \cu_ru/m_cycle_event/add1/c15 ;
  wire \cu_ru/m_cycle_event/add1/c16 ;
  wire \cu_ru/m_cycle_event/add1/c17 ;
  wire \cu_ru/m_cycle_event/add1/c18 ;
  wire \cu_ru/m_cycle_event/add1/c19 ;
  wire \cu_ru/m_cycle_event/add1/c2 ;
  wire \cu_ru/m_cycle_event/add1/c20 ;
  wire \cu_ru/m_cycle_event/add1/c21 ;
  wire \cu_ru/m_cycle_event/add1/c22 ;
  wire \cu_ru/m_cycle_event/add1/c23 ;
  wire \cu_ru/m_cycle_event/add1/c24 ;
  wire \cu_ru/m_cycle_event/add1/c25 ;
  wire \cu_ru/m_cycle_event/add1/c26 ;
  wire \cu_ru/m_cycle_event/add1/c27 ;
  wire \cu_ru/m_cycle_event/add1/c28 ;
  wire \cu_ru/m_cycle_event/add1/c29 ;
  wire \cu_ru/m_cycle_event/add1/c3 ;
  wire \cu_ru/m_cycle_event/add1/c30 ;
  wire \cu_ru/m_cycle_event/add1/c31 ;
  wire \cu_ru/m_cycle_event/add1/c32 ;
  wire \cu_ru/m_cycle_event/add1/c33 ;
  wire \cu_ru/m_cycle_event/add1/c34 ;
  wire \cu_ru/m_cycle_event/add1/c35 ;
  wire \cu_ru/m_cycle_event/add1/c36 ;
  wire \cu_ru/m_cycle_event/add1/c37 ;
  wire \cu_ru/m_cycle_event/add1/c38 ;
  wire \cu_ru/m_cycle_event/add1/c39 ;
  wire \cu_ru/m_cycle_event/add1/c4 ;
  wire \cu_ru/m_cycle_event/add1/c40 ;
  wire \cu_ru/m_cycle_event/add1/c41 ;
  wire \cu_ru/m_cycle_event/add1/c42 ;
  wire \cu_ru/m_cycle_event/add1/c43 ;
  wire \cu_ru/m_cycle_event/add1/c44 ;
  wire \cu_ru/m_cycle_event/add1/c45 ;
  wire \cu_ru/m_cycle_event/add1/c46 ;
  wire \cu_ru/m_cycle_event/add1/c47 ;
  wire \cu_ru/m_cycle_event/add1/c48 ;
  wire \cu_ru/m_cycle_event/add1/c49 ;
  wire \cu_ru/m_cycle_event/add1/c5 ;
  wire \cu_ru/m_cycle_event/add1/c50 ;
  wire \cu_ru/m_cycle_event/add1/c51 ;
  wire \cu_ru/m_cycle_event/add1/c52 ;
  wire \cu_ru/m_cycle_event/add1/c53 ;
  wire \cu_ru/m_cycle_event/add1/c54 ;
  wire \cu_ru/m_cycle_event/add1/c55 ;
  wire \cu_ru/m_cycle_event/add1/c56 ;
  wire \cu_ru/m_cycle_event/add1/c57 ;
  wire \cu_ru/m_cycle_event/add1/c58 ;
  wire \cu_ru/m_cycle_event/add1/c59 ;
  wire \cu_ru/m_cycle_event/add1/c6 ;
  wire \cu_ru/m_cycle_event/add1/c60 ;
  wire \cu_ru/m_cycle_event/add1/c61 ;
  wire \cu_ru/m_cycle_event/add1/c62 ;
  wire \cu_ru/m_cycle_event/add1/c63 ;
  wire \cu_ru/m_cycle_event/add1/c7 ;
  wire \cu_ru/m_cycle_event/add1/c8 ;
  wire \cu_ru/m_cycle_event/add1/c9 ;
  wire \cu_ru/m_cycle_event/mcountinhibit[2] ;  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(16)
  wire \cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ;
  wire \cu_ru/m_cycle_event/n13 ;
  wire \cu_ru/m_s_cause/mux2_b0_sel_is_2_o ;
  wire \cu_ru/m_s_cause/mux4_b0_sel_is_2_o ;
  wire \cu_ru/m_s_cause/mux7_b10_sel_is_0_o ;
  wire \cu_ru/m_s_epc/add0/c0 ;
  wire \cu_ru/m_s_epc/add0/c1 ;
  wire \cu_ru/m_s_epc/add0/c10 ;
  wire \cu_ru/m_s_epc/add0/c11 ;
  wire \cu_ru/m_s_epc/add0/c12 ;
  wire \cu_ru/m_s_epc/add0/c13 ;
  wire \cu_ru/m_s_epc/add0/c14 ;
  wire \cu_ru/m_s_epc/add0/c15 ;
  wire \cu_ru/m_s_epc/add0/c16 ;
  wire \cu_ru/m_s_epc/add0/c17 ;
  wire \cu_ru/m_s_epc/add0/c18 ;
  wire \cu_ru/m_s_epc/add0/c19 ;
  wire \cu_ru/m_s_epc/add0/c2 ;
  wire \cu_ru/m_s_epc/add0/c20 ;
  wire \cu_ru/m_s_epc/add0/c21 ;
  wire \cu_ru/m_s_epc/add0/c22 ;
  wire \cu_ru/m_s_epc/add0/c23 ;
  wire \cu_ru/m_s_epc/add0/c24 ;
  wire \cu_ru/m_s_epc/add0/c25 ;
  wire \cu_ru/m_s_epc/add0/c26 ;
  wire \cu_ru/m_s_epc/add0/c27 ;
  wire \cu_ru/m_s_epc/add0/c28 ;
  wire \cu_ru/m_s_epc/add0/c29 ;
  wire \cu_ru/m_s_epc/add0/c3 ;
  wire \cu_ru/m_s_epc/add0/c30 ;
  wire \cu_ru/m_s_epc/add0/c31 ;
  wire \cu_ru/m_s_epc/add0/c32 ;
  wire \cu_ru/m_s_epc/add0/c33 ;
  wire \cu_ru/m_s_epc/add0/c34 ;
  wire \cu_ru/m_s_epc/add0/c35 ;
  wire \cu_ru/m_s_epc/add0/c36 ;
  wire \cu_ru/m_s_epc/add0/c37 ;
  wire \cu_ru/m_s_epc/add0/c38 ;
  wire \cu_ru/m_s_epc/add0/c39 ;
  wire \cu_ru/m_s_epc/add0/c4 ;
  wire \cu_ru/m_s_epc/add0/c40 ;
  wire \cu_ru/m_s_epc/add0/c41 ;
  wire \cu_ru/m_s_epc/add0/c42 ;
  wire \cu_ru/m_s_epc/add0/c43 ;
  wire \cu_ru/m_s_epc/add0/c44 ;
  wire \cu_ru/m_s_epc/add0/c45 ;
  wire \cu_ru/m_s_epc/add0/c46 ;
  wire \cu_ru/m_s_epc/add0/c47 ;
  wire \cu_ru/m_s_epc/add0/c48 ;
  wire \cu_ru/m_s_epc/add0/c49 ;
  wire \cu_ru/m_s_epc/add0/c5 ;
  wire \cu_ru/m_s_epc/add0/c50 ;
  wire \cu_ru/m_s_epc/add0/c51 ;
  wire \cu_ru/m_s_epc/add0/c52 ;
  wire \cu_ru/m_s_epc/add0/c53 ;
  wire \cu_ru/m_s_epc/add0/c54 ;
  wire \cu_ru/m_s_epc/add0/c55 ;
  wire \cu_ru/m_s_epc/add0/c56 ;
  wire \cu_ru/m_s_epc/add0/c57 ;
  wire \cu_ru/m_s_epc/add0/c58 ;
  wire \cu_ru/m_s_epc/add0/c59 ;
  wire \cu_ru/m_s_epc/add0/c6 ;
  wire \cu_ru/m_s_epc/add0/c60 ;
  wire \cu_ru/m_s_epc/add0/c61 ;
  wire \cu_ru/m_s_epc/add0/c7 ;
  wire \cu_ru/m_s_epc/add0/c8 ;
  wire \cu_ru/m_s_epc/add0/c9 ;
  wire \cu_ru/m_s_epc/mux4_b0_sel_is_2_o ;
  wire \cu_ru/m_s_epc/mux6_b0_sel_is_2_o ;
  wire \cu_ru/m_s_ie/n0 ;
  wire \cu_ru/m_s_ie/u11_sel_is_0_o ;
  wire \cu_ru/m_s_ip/n0 ;
  wire \cu_ru/m_s_ip/n1 ;
  wire \cu_ru/m_s_ip/seip ;  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(28)
  wire \cu_ru/m_s_ip/u11_sel_is_0_o ;
  wire \cu_ru/m_s_ip/u12_sel_is_2_o ;
  wire \cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ;
  wire \cu_ru/m_s_scratch/n0 ;
  wire \cu_ru/m_s_status/mux3_b0_sel_is_2_o ;
  wire \cu_ru/m_s_status/n0 ;
  wire \cu_ru/m_s_status/n2 ;
  wire \cu_ru/m_s_status/n36 ;
  wire \cu_ru/m_s_status/n37 ;
  wire \cu_ru/m_s_status/n44 ;
  wire \cu_ru/m_s_status/n45 ;
  wire \cu_ru/m_s_status/n46 ;
  wire \cu_ru/m_s_status/u14_sel_is_2_o ;
  wire \cu_ru/m_s_status/u34_sel_is_0_o ;
  wire \cu_ru/m_s_tval/mux3_b0_sel_is_2_o ;
  wire \cu_ru/m_s_tval/mux5_b0_sel_is_2_o ;
  wire \cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ;
  wire \cu_ru/m_s_tvec/n0 ;
  wire \cu_ru/mcountinhibit ;  // ../../RTL/CPU/CU&RU/cu_ru.v(639)
  wire \cu_ru/medeleg_exc_ctrl/ecu_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(78)
  wire \cu_ru/medeleg_exc_ctrl/ecu_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(92)
  wire \cu_ru/medeleg_exc_ctrl/iaf_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(71)
  wire \cu_ru/medeleg_exc_ctrl/iam_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(70)
  wire \cu_ru/medeleg_exc_ctrl/iam_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(84)
  wire \cu_ru/medeleg_exc_ctrl/ii_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(86)
  wire \cu_ru/medeleg_exc_ctrl/laf_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(75)
  wire \cu_ru/medeleg_exc_ctrl/laf_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(89)
  wire \cu_ru/medeleg_exc_ctrl/lam_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(74)
  wire \cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/n0 ;
  wire \cu_ru/medeleg_exc_ctrl/n80_neg_lutinv ;
  wire \cu_ru/medeleg_exc_ctrl/n84_neg_lutinv ;
  wire \cu_ru/medeleg_exc_ctrl/n85_neg_lutinv ;
  wire \cu_ru/medeleg_exc_ctrl/n87_neg_lutinv ;
  wire \cu_ru/medeleg_exc_ctrl/saf_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(77)
  wire \cu_ru/medeleg_exc_ctrl/sam_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(90)
  wire \cu_ru/medeleg_exc_ctrl/spf_target_m_lutinv ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(82)
  wire \cu_ru/medeleg_exc_ctrl/spf_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(96)
  wire \cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o ;
  wire \cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ;
  wire \cu_ru/mideleg_int_ctrl/n0 ;
  wire \cu_ru/mideleg_int_ctrl/n28_lutinv ;
  wire \cu_ru/mideleg_int_ctrl/n29_lutinv ;
  wire \cu_ru/mideleg_int_ctrl/n33_neg_lutinv ;
  wire \cu_ru/mideleg_int_ctrl/sei_ack_m ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(61)
  wire \cu_ru/mideleg_int_ctrl/sti_ack_s ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(67)
  wire \cu_ru/mie ;  // ../../RTL/CPU/CU&RU/cu_ru.v(381)
  wire \cu_ru/mux34_b0_sel_is_2_o ;
  wire \cu_ru/n41 ;
  wire \cu_ru/n45_lutinv ;
  wire \cu_ru/n53_0_al_n1985 ;
  wire \cu_ru/n53_1_al_n1986 ;
  wire \cu_ru/n53_lutinv ;
  wire \cu_ru/n66_lutinv ;
  wire \cu_ru/read_cycle_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(220)
  wire \cu_ru/read_instret_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(222)
  wire \cu_ru/read_mcause_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(248)
  wire \cu_ru/read_mcycle_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(254)
  wire \cu_ru/read_medeleg_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(241)
  wire \cu_ru/read_mepc_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(247)
  wire \cu_ru/read_mideleg_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(242)
  wire \cu_ru/read_minstret_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(255)
  wire \cu_ru/read_mip_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(250)
  wire \cu_ru/read_mscratch_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(246)
  wire \cu_ru/read_mtval_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(249)
  wire \cu_ru/read_mtvec_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(244)
  wire \cu_ru/read_satp_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(234)
  wire \cu_ru/read_scause_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(231)
  wire \cu_ru/read_sepc_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(230)
  wire \cu_ru/read_sscratch_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(229)
  wire \cu_ru/read_stval_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(232)
  wire \cu_ru/read_stvec_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(227)
  wire \cu_ru/read_time_sel_lutinv ;  // ../../RTL/CPU/CU&RU/cu_ru.v(221)
  wire \cu_ru/sub0/c0 ;
  wire \cu_ru/sub0/c1 ;
  wire \cu_ru/sub0/c2 ;
  wire \cu_ru/sub0/c3 ;
  wire \cu_ru/sub0/c4 ;
  wire \cu_ru/sub1/c0 ;
  wire \cu_ru/sub1/c1 ;
  wire \cu_ru/sub1/c2 ;
  wire \cu_ru/sub1/c3 ;
  wire \cu_ru/sub1/c4 ;
  wire \cu_ru/sub2/c0 ;
  wire \cu_ru/sub2/c1 ;
  wire \cu_ru/sub2/c2 ;
  wire \cu_ru/sub2/c3 ;
  wire \cu_ru/sub2/c4 ;
  wire \cu_ru/trap_target_m ;  // ../../RTL/CPU/CU&RU/cu_ru.v(148)
  wire ex_csr_write;  // ../../RTL/CPU/prv464_top.v(145)
  wire ex_ebreak;  // ../../RTL/CPU/prv464_top.v(171)
  wire ex_ecall;  // ../../RTL/CPU/prv464_top.v(170)
  wire ex_gpr_write;  // ../../RTL/CPU/prv464_top.v(146)
  wire ex_ill_ins;  // ../../RTL/CPU/prv464_top.v(167)
  wire ex_ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(162)
  wire ex_ins_addr_mis;  // ../../RTL/CPU/prv464_top.v(163)
  wire ex_ins_page_fault;  // ../../RTL/CPU/prv464_top.v(164)
  wire ex_int_acc;  // ../../RTL/CPU/prv464_top.v(165)
  wire ex_jmp;  // ../../RTL/CPU/prv464_top.v(161)
  wire ex_m_ret;  // ../../RTL/CPU/prv464_top.v(168)
  wire ex_more_exception_neg_lutinv;
  wire ex_nop;  // ../../RTL/CPU/prv464_top.v(580)
  wire ex_s_ret;  // ../../RTL/CPU/prv464_top.v(169)
  wire ex_system;  // ../../RTL/CPU/prv464_top.v(160)
  wire ex_valid;  // ../../RTL/CPU/prv464_top.v(166)
  wire \exu/alu_au/add0/c0 ;
  wire \exu/alu_au/add0/c1 ;
  wire \exu/alu_au/add0/c10 ;
  wire \exu/alu_au/add0/c11 ;
  wire \exu/alu_au/add0/c12 ;
  wire \exu/alu_au/add0/c13 ;
  wire \exu/alu_au/add0/c14 ;
  wire \exu/alu_au/add0/c15 ;
  wire \exu/alu_au/add0/c16 ;
  wire \exu/alu_au/add0/c17 ;
  wire \exu/alu_au/add0/c18 ;
  wire \exu/alu_au/add0/c19 ;
  wire \exu/alu_au/add0/c2 ;
  wire \exu/alu_au/add0/c20 ;
  wire \exu/alu_au/add0/c21 ;
  wire \exu/alu_au/add0/c22 ;
  wire \exu/alu_au/add0/c23 ;
  wire \exu/alu_au/add0/c24 ;
  wire \exu/alu_au/add0/c25 ;
  wire \exu/alu_au/add0/c26 ;
  wire \exu/alu_au/add0/c27 ;
  wire \exu/alu_au/add0/c28 ;
  wire \exu/alu_au/add0/c29 ;
  wire \exu/alu_au/add0/c3 ;
  wire \exu/alu_au/add0/c30 ;
  wire \exu/alu_au/add0/c31 ;
  wire \exu/alu_au/add0/c32 ;
  wire \exu/alu_au/add0/c33 ;
  wire \exu/alu_au/add0/c34 ;
  wire \exu/alu_au/add0/c35 ;
  wire \exu/alu_au/add0/c36 ;
  wire \exu/alu_au/add0/c37 ;
  wire \exu/alu_au/add0/c38 ;
  wire \exu/alu_au/add0/c39 ;
  wire \exu/alu_au/add0/c4 ;
  wire \exu/alu_au/add0/c40 ;
  wire \exu/alu_au/add0/c41 ;
  wire \exu/alu_au/add0/c42 ;
  wire \exu/alu_au/add0/c43 ;
  wire \exu/alu_au/add0/c44 ;
  wire \exu/alu_au/add0/c45 ;
  wire \exu/alu_au/add0/c46 ;
  wire \exu/alu_au/add0/c47 ;
  wire \exu/alu_au/add0/c48 ;
  wire \exu/alu_au/add0/c49 ;
  wire \exu/alu_au/add0/c5 ;
  wire \exu/alu_au/add0/c50 ;
  wire \exu/alu_au/add0/c51 ;
  wire \exu/alu_au/add0/c52 ;
  wire \exu/alu_au/add0/c53 ;
  wire \exu/alu_au/add0/c54 ;
  wire \exu/alu_au/add0/c55 ;
  wire \exu/alu_au/add0/c56 ;
  wire \exu/alu_au/add0/c57 ;
  wire \exu/alu_au/add0/c58 ;
  wire \exu/alu_au/add0/c59 ;
  wire \exu/alu_au/add0/c6 ;
  wire \exu/alu_au/add0/c60 ;
  wire \exu/alu_au/add0/c61 ;
  wire \exu/alu_au/add0/c62 ;
  wire \exu/alu_au/add0/c63 ;
  wire \exu/alu_au/add0/c7 ;
  wire \exu/alu_au/add0/c8 ;
  wire \exu/alu_au/add0/c9 ;
  wire \exu/alu_au/add1/c0 ;
  wire \exu/alu_au/add1/c1 ;
  wire \exu/alu_au/add1/c10 ;
  wire \exu/alu_au/add1/c11 ;
  wire \exu/alu_au/add1/c12 ;
  wire \exu/alu_au/add1/c13 ;
  wire \exu/alu_au/add1/c14 ;
  wire \exu/alu_au/add1/c15 ;
  wire \exu/alu_au/add1/c16 ;
  wire \exu/alu_au/add1/c17 ;
  wire \exu/alu_au/add1/c18 ;
  wire \exu/alu_au/add1/c19 ;
  wire \exu/alu_au/add1/c2 ;
  wire \exu/alu_au/add1/c20 ;
  wire \exu/alu_au/add1/c21 ;
  wire \exu/alu_au/add1/c22 ;
  wire \exu/alu_au/add1/c23 ;
  wire \exu/alu_au/add1/c24 ;
  wire \exu/alu_au/add1/c25 ;
  wire \exu/alu_au/add1/c26 ;
  wire \exu/alu_au/add1/c27 ;
  wire \exu/alu_au/add1/c28 ;
  wire \exu/alu_au/add1/c29 ;
  wire \exu/alu_au/add1/c3 ;
  wire \exu/alu_au/add1/c30 ;
  wire \exu/alu_au/add1/c31 ;
  wire \exu/alu_au/add1/c4 ;
  wire \exu/alu_au/add1/c5 ;
  wire \exu/alu_au/add1/c6 ;
  wire \exu/alu_au/add1/c7 ;
  wire \exu/alu_au/add1/c8 ;
  wire \exu/alu_au/add1/c9 ;
  wire \exu/alu_au/add2/c0 ;
  wire \exu/alu_au/add2/c1 ;
  wire \exu/alu_au/add2/c10 ;
  wire \exu/alu_au/add2/c11 ;
  wire \exu/alu_au/add2/c12 ;
  wire \exu/alu_au/add2/c13 ;
  wire \exu/alu_au/add2/c14 ;
  wire \exu/alu_au/add2/c15 ;
  wire \exu/alu_au/add2/c16 ;
  wire \exu/alu_au/add2/c17 ;
  wire \exu/alu_au/add2/c18 ;
  wire \exu/alu_au/add2/c19 ;
  wire \exu/alu_au/add2/c2 ;
  wire \exu/alu_au/add2/c20 ;
  wire \exu/alu_au/add2/c21 ;
  wire \exu/alu_au/add2/c22 ;
  wire \exu/alu_au/add2/c23 ;
  wire \exu/alu_au/add2/c24 ;
  wire \exu/alu_au/add2/c25 ;
  wire \exu/alu_au/add2/c26 ;
  wire \exu/alu_au/add2/c27 ;
  wire \exu/alu_au/add2/c28 ;
  wire \exu/alu_au/add2/c29 ;
  wire \exu/alu_au/add2/c3 ;
  wire \exu/alu_au/add2/c30 ;
  wire \exu/alu_au/add2/c31 ;
  wire \exu/alu_au/add2/c32 ;
  wire \exu/alu_au/add2/c33 ;
  wire \exu/alu_au/add2/c34 ;
  wire \exu/alu_au/add2/c35 ;
  wire \exu/alu_au/add2/c36 ;
  wire \exu/alu_au/add2/c37 ;
  wire \exu/alu_au/add2/c38 ;
  wire \exu/alu_au/add2/c39 ;
  wire \exu/alu_au/add2/c4 ;
  wire \exu/alu_au/add2/c40 ;
  wire \exu/alu_au/add2/c41 ;
  wire \exu/alu_au/add2/c42 ;
  wire \exu/alu_au/add2/c43 ;
  wire \exu/alu_au/add2/c44 ;
  wire \exu/alu_au/add2/c45 ;
  wire \exu/alu_au/add2/c46 ;
  wire \exu/alu_au/add2/c47 ;
  wire \exu/alu_au/add2/c48 ;
  wire \exu/alu_au/add2/c49 ;
  wire \exu/alu_au/add2/c5 ;
  wire \exu/alu_au/add2/c50 ;
  wire \exu/alu_au/add2/c51 ;
  wire \exu/alu_au/add2/c52 ;
  wire \exu/alu_au/add2/c53 ;
  wire \exu/alu_au/add2/c54 ;
  wire \exu/alu_au/add2/c55 ;
  wire \exu/alu_au/add2/c56 ;
  wire \exu/alu_au/add2/c57 ;
  wire \exu/alu_au/add2/c58 ;
  wire \exu/alu_au/add2/c59 ;
  wire \exu/alu_au/add2/c6 ;
  wire \exu/alu_au/add2/c60 ;
  wire \exu/alu_au/add2/c61 ;
  wire \exu/alu_au/add2/c62 ;
  wire \exu/alu_au/add2/c63 ;
  wire \exu/alu_au/add2/c7 ;
  wire \exu/alu_au/add2/c8 ;
  wire \exu/alu_au/add2/c9 ;
  wire \exu/alu_au/ds1_light_than_ds2_lutinv ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(67)
  wire \exu/alu_au/lt0_c0 ;
  wire \exu/alu_au/lt0_c1 ;
  wire \exu/alu_au/lt0_c10 ;
  wire \exu/alu_au/lt0_c11 ;
  wire \exu/alu_au/lt0_c12 ;
  wire \exu/alu_au/lt0_c13 ;
  wire \exu/alu_au/lt0_c14 ;
  wire \exu/alu_au/lt0_c15 ;
  wire \exu/alu_au/lt0_c16 ;
  wire \exu/alu_au/lt0_c17 ;
  wire \exu/alu_au/lt0_c18 ;
  wire \exu/alu_au/lt0_c19 ;
  wire \exu/alu_au/lt0_c2 ;
  wire \exu/alu_au/lt0_c20 ;
  wire \exu/alu_au/lt0_c21 ;
  wire \exu/alu_au/lt0_c22 ;
  wire \exu/alu_au/lt0_c23 ;
  wire \exu/alu_au/lt0_c24 ;
  wire \exu/alu_au/lt0_c25 ;
  wire \exu/alu_au/lt0_c26 ;
  wire \exu/alu_au/lt0_c27 ;
  wire \exu/alu_au/lt0_c28 ;
  wire \exu/alu_au/lt0_c29 ;
  wire \exu/alu_au/lt0_c3 ;
  wire \exu/alu_au/lt0_c30 ;
  wire \exu/alu_au/lt0_c31 ;
  wire \exu/alu_au/lt0_c32 ;
  wire \exu/alu_au/lt0_c33 ;
  wire \exu/alu_au/lt0_c34 ;
  wire \exu/alu_au/lt0_c35 ;
  wire \exu/alu_au/lt0_c36 ;
  wire \exu/alu_au/lt0_c37 ;
  wire \exu/alu_au/lt0_c38 ;
  wire \exu/alu_au/lt0_c39 ;
  wire \exu/alu_au/lt0_c4 ;
  wire \exu/alu_au/lt0_c40 ;
  wire \exu/alu_au/lt0_c41 ;
  wire \exu/alu_au/lt0_c42 ;
  wire \exu/alu_au/lt0_c43 ;
  wire \exu/alu_au/lt0_c44 ;
  wire \exu/alu_au/lt0_c45 ;
  wire \exu/alu_au/lt0_c46 ;
  wire \exu/alu_au/lt0_c47 ;
  wire \exu/alu_au/lt0_c48 ;
  wire \exu/alu_au/lt0_c49 ;
  wire \exu/alu_au/lt0_c5 ;
  wire \exu/alu_au/lt0_c50 ;
  wire \exu/alu_au/lt0_c51 ;
  wire \exu/alu_au/lt0_c52 ;
  wire \exu/alu_au/lt0_c53 ;
  wire \exu/alu_au/lt0_c54 ;
  wire \exu/alu_au/lt0_c55 ;
  wire \exu/alu_au/lt0_c56 ;
  wire \exu/alu_au/lt0_c57 ;
  wire \exu/alu_au/lt0_c58 ;
  wire \exu/alu_au/lt0_c59 ;
  wire \exu/alu_au/lt0_c6 ;
  wire \exu/alu_au/lt0_c60 ;
  wire \exu/alu_au/lt0_c61 ;
  wire \exu/alu_au/lt0_c62 ;
  wire \exu/alu_au/lt0_c63 ;
  wire \exu/alu_au/lt0_c64 ;
  wire \exu/alu_au/lt0_c7 ;
  wire \exu/alu_au/lt0_c8 ;
  wire \exu/alu_au/lt0_c9 ;
  wire \exu/alu_au/lt1_c0 ;
  wire \exu/alu_au/lt1_c1 ;
  wire \exu/alu_au/lt1_c10 ;
  wire \exu/alu_au/lt1_c11 ;
  wire \exu/alu_au/lt1_c12 ;
  wire \exu/alu_au/lt1_c13 ;
  wire \exu/alu_au/lt1_c14 ;
  wire \exu/alu_au/lt1_c15 ;
  wire \exu/alu_au/lt1_c16 ;
  wire \exu/alu_au/lt1_c17 ;
  wire \exu/alu_au/lt1_c18 ;
  wire \exu/alu_au/lt1_c19 ;
  wire \exu/alu_au/lt1_c2 ;
  wire \exu/alu_au/lt1_c20 ;
  wire \exu/alu_au/lt1_c21 ;
  wire \exu/alu_au/lt1_c22 ;
  wire \exu/alu_au/lt1_c23 ;
  wire \exu/alu_au/lt1_c24 ;
  wire \exu/alu_au/lt1_c25 ;
  wire \exu/alu_au/lt1_c26 ;
  wire \exu/alu_au/lt1_c27 ;
  wire \exu/alu_au/lt1_c28 ;
  wire \exu/alu_au/lt1_c29 ;
  wire \exu/alu_au/lt1_c3 ;
  wire \exu/alu_au/lt1_c30 ;
  wire \exu/alu_au/lt1_c31 ;
  wire \exu/alu_au/lt1_c32 ;
  wire \exu/alu_au/lt1_c33 ;
  wire \exu/alu_au/lt1_c34 ;
  wire \exu/alu_au/lt1_c35 ;
  wire \exu/alu_au/lt1_c36 ;
  wire \exu/alu_au/lt1_c37 ;
  wire \exu/alu_au/lt1_c38 ;
  wire \exu/alu_au/lt1_c39 ;
  wire \exu/alu_au/lt1_c4 ;
  wire \exu/alu_au/lt1_c40 ;
  wire \exu/alu_au/lt1_c41 ;
  wire \exu/alu_au/lt1_c42 ;
  wire \exu/alu_au/lt1_c43 ;
  wire \exu/alu_au/lt1_c44 ;
  wire \exu/alu_au/lt1_c45 ;
  wire \exu/alu_au/lt1_c46 ;
  wire \exu/alu_au/lt1_c47 ;
  wire \exu/alu_au/lt1_c48 ;
  wire \exu/alu_au/lt1_c49 ;
  wire \exu/alu_au/lt1_c5 ;
  wire \exu/alu_au/lt1_c50 ;
  wire \exu/alu_au/lt1_c51 ;
  wire \exu/alu_au/lt1_c52 ;
  wire \exu/alu_au/lt1_c53 ;
  wire \exu/alu_au/lt1_c54 ;
  wire \exu/alu_au/lt1_c55 ;
  wire \exu/alu_au/lt1_c56 ;
  wire \exu/alu_au/lt1_c57 ;
  wire \exu/alu_au/lt1_c58 ;
  wire \exu/alu_au/lt1_c59 ;
  wire \exu/alu_au/lt1_c6 ;
  wire \exu/alu_au/lt1_c60 ;
  wire \exu/alu_au/lt1_c61 ;
  wire \exu/alu_au/lt1_c62 ;
  wire \exu/alu_au/lt1_c63 ;
  wire \exu/alu_au/lt1_c64 ;
  wire \exu/alu_au/lt1_c7 ;
  wire \exu/alu_au/lt1_c8 ;
  wire \exu/alu_au/lt1_c9 ;
  wire \exu/alu_au/n12 ;
  wire \exu/alu_au/n15 ;
  wire \exu/alu_au/n5 ;
  wire \exu/c_fence_lutinv ;  // ../../RTL/CPU/EX/exu.v(182)
  wire \exu/c_load_1_lutinv ;  // ../../RTL/CPU/EX/exu.v(176)
  wire \exu/c_stb_lutinv ;  // ../../RTL/CPU/EX/exu.v(173)
  wire \exu/load_addr_mis ;  // ../../RTL/CPU/EX/exu.v(202)
  wire \exu/lsu/mux27_b56_sel_is_3_o ;
  wire \exu/lsu/n0_lutinv ;
  wire \exu/lsu/n2_lutinv ;
  wire \exu/lsu/n51 ;
  wire \exu/lsu/n53 ;
  wire \exu/lsu/n56 ;
  wire \exu/lsu/n5_lutinv ;
  wire \exu/lsu/n8_lutinv ;
  wire \exu/mux27_b32_sel_is_1_o ;
  wire \exu/n10 ;
  wire \exu/n138_lutinv ;
  wire \exu/n17_lutinv ;
  wire \exu/n19 ;
  wire \exu/n49 ;
  wire \exu/n59_lutinv ;
  wire \exu/n60_lutinv ;
  wire \exu/n86 ;
  wire \exu/n88 ;
  wire \exu/n90 ;
  wire \exu/n92 ;
  wire \exu/n95 ;
  wire \exu/shift_multi_ready ;  // ../../RTL/CPU/EX/exu.v(209)
  wire \exu/store_addr_mis ;  // ../../RTL/CPU/EX/exu.v(203)
  wire \exu/sub0/c0 ;
  wire \exu/sub0/c1 ;
  wire \exu/sub0/c2 ;
  wire \exu/sub0/c3 ;
  wire \exu/sub0/c4 ;
  wire \exu/sub0/c5 ;
  wire \exu/sub0/c6 ;
  wire \exu/sub0/c7 ;
  wire hready_pad;  // ../../RTL/CPU/prv464_top.v(31)
  wire hresp_pad;  // ../../RTL/CPU/prv464_top.v(32)
  wire hwrite_pad;  // ../../RTL/CPU/prv464_top.v(23)
  wire id_hold;  // ../../RTL/CPU/prv464_top.v(177)
  wire id_ill_ins;  // ../../RTL/CPU/prv464_top.v(176)
  wire id_ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(92)
  wire id_ins_addr_mis;  // ../../RTL/CPU/prv464_top.v(93)
  wire id_ins_page_fault;  // ../../RTL/CPU/prv464_top.v(94)
  wire id_int_acc;  // ../../RTL/CPU/prv464_top.v(95)
  wire id_nop_neg_lutinv;
  wire id_system;  // ../../RTL/CPU/prv464_top.v(175)
  wire id_valid;  // ../../RTL/CPU/prv464_top.v(96)
  wire if_hold;  // ../../RTL/CPU/prv464_top.v(263)
  wire ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(68)
  wire \ins_dec/dbyte ;  // ../../RTL/CPU/ID/ins_dec.v(235)
  wire \ins_dec/dec_gpr_write ;  // ../../RTL/CPU/ID/ins_dec.v(119)
  wire \ins_dec/dec_ins_dec_fault_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(336)
  wire \ins_dec/funct3_0_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(172)
  wire \ins_dec/funct5_8_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(189)
  wire \ins_dec/funct6_0_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(214)
  wire \ins_dec/funct7_0_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(220)
  wire \ins_dec/funct7_32_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(217)
  wire \ins_dec/funct7_8_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(219)
  wire \ins_dec/ins_addw ;  // ../../RTL/CPU/ID/ins_dec.v(299)
  wire \ins_dec/ins_ebreak ;  // ../../RTL/CPU/ID/ins_dec.v(284)
  wire \ins_dec/ins_ecall ;  // ../../RTL/CPU/ID/ins_dec.v(283)
  wire \ins_dec/ins_fence ;  // ../../RTL/CPU/ID/ins_dec.v(282)
  wire \ins_dec/ins_sfencevma ;  // ../../RTL/CPU/ID/ins_dec.v(331)
  wire \ins_dec/ins_slli ;  // ../../RTL/CPU/ID/ins_dec.v(269)
  wire \ins_dec/ins_srai ;  // ../../RTL/CPU/ID/ins_dec.v(271)
  wire \ins_dec/ins_srli ;  // ../../RTL/CPU/ID/ins_dec.v(270)
  wire \ins_dec/mux13_b0_sel_is_0_o ;
  wire \ins_dec/mux19_b10_sel_is_2_o ;
  wire \ins_dec/mux24_b10_sel_is_0_o ;
  wire \ins_dec/mux27_b12_sel_is_0_o ;
  wire \ins_dec/mux27_b56_sel_is_0_o ;
  wire \ins_dec/n107 ;
  wire \ins_dec/n126 ;
  wire \ins_dec/n132 ;
  wire \ins_dec/n133 ;
  wire \ins_dec/n134 ;
  wire \ins_dec/n135 ;
  wire \ins_dec/n136 ;
  wire \ins_dec/n139 ;
  wire \ins_dec/n141_lutinv ;
  wire \ins_dec/n145 ;
  wire \ins_dec/n146 ;
  wire \ins_dec/n148 ;
  wire \ins_dec/n149_lutinv ;
  wire \ins_dec/n151 ;
  wire \ins_dec/n152 ;
  wire \ins_dec/n155 ;
  wire \ins_dec/n158 ;
  wire \ins_dec/n198_lutinv ;
  wire \ins_dec/n206 ;
  wire \ins_dec/n225 ;
  wire \ins_dec/n232 ;
  wire \ins_dec/n235 ;
  wire \ins_dec/n239 ;
  wire \ins_dec/n302 ;
  wire \ins_dec/n35_lutinv ;
  wire \ins_dec/n38 ;
  wire \ins_dec/n48_lutinv ;
  wire \ins_dec/n57_neg_lutinv ;
  wire \ins_dec/n59 ;
  wire \ins_dec/n71 ;
  wire \ins_dec/n80_lutinv ;
  wire \ins_dec/obyte ;  // ../../RTL/CPU/ID/ins_dec.v(237)
  wire \ins_dec/op_32_imm_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(158)
  wire \ins_dec/op_32_reg_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(167)
  wire \ins_dec/op_amo ;  // ../../RTL/CPU/ID/ins_dec.v(168)
  wire \ins_dec/op_load ;  // ../../RTL/CPU/ID/ins_dec.v(165)
  wire \ins_dec/op_lui_lutinv ;  // ../../RTL/CPU/ID/ins_dec.v(159)
  wire \ins_dec/op_store ;  // ../../RTL/CPU/ID/ins_dec.v(164)
  wire \ins_dec/qbyte ;  // ../../RTL/CPU/ID/ins_dec.v(236)
  wire \ins_dec/sbyte ;  // ../../RTL/CPU/ID/ins_dec.v(234)
  wire \ins_dec/u461_sel_is_0_o ;
  wire \ins_dec/u478_sel_is_0_o ;
  wire \ins_fetch/add0/c0 ;
  wire \ins_fetch/add0/c1 ;
  wire \ins_fetch/add0/c10 ;
  wire \ins_fetch/add0/c11 ;
  wire \ins_fetch/add0/c12 ;
  wire \ins_fetch/add0/c13 ;
  wire \ins_fetch/add0/c14 ;
  wire \ins_fetch/add0/c15 ;
  wire \ins_fetch/add0/c16 ;
  wire \ins_fetch/add0/c17 ;
  wire \ins_fetch/add0/c18 ;
  wire \ins_fetch/add0/c19 ;
  wire \ins_fetch/add0/c2 ;
  wire \ins_fetch/add0/c20 ;
  wire \ins_fetch/add0/c21 ;
  wire \ins_fetch/add0/c22 ;
  wire \ins_fetch/add0/c23 ;
  wire \ins_fetch/add0/c24 ;
  wire \ins_fetch/add0/c25 ;
  wire \ins_fetch/add0/c26 ;
  wire \ins_fetch/add0/c27 ;
  wire \ins_fetch/add0/c28 ;
  wire \ins_fetch/add0/c29 ;
  wire \ins_fetch/add0/c3 ;
  wire \ins_fetch/add0/c30 ;
  wire \ins_fetch/add0/c31 ;
  wire \ins_fetch/add0/c32 ;
  wire \ins_fetch/add0/c33 ;
  wire \ins_fetch/add0/c34 ;
  wire \ins_fetch/add0/c35 ;
  wire \ins_fetch/add0/c36 ;
  wire \ins_fetch/add0/c37 ;
  wire \ins_fetch/add0/c38 ;
  wire \ins_fetch/add0/c39 ;
  wire \ins_fetch/add0/c4 ;
  wire \ins_fetch/add0/c40 ;
  wire \ins_fetch/add0/c41 ;
  wire \ins_fetch/add0/c42 ;
  wire \ins_fetch/add0/c43 ;
  wire \ins_fetch/add0/c44 ;
  wire \ins_fetch/add0/c45 ;
  wire \ins_fetch/add0/c46 ;
  wire \ins_fetch/add0/c47 ;
  wire \ins_fetch/add0/c48 ;
  wire \ins_fetch/add0/c49 ;
  wire \ins_fetch/add0/c5 ;
  wire \ins_fetch/add0/c50 ;
  wire \ins_fetch/add0/c51 ;
  wire \ins_fetch/add0/c52 ;
  wire \ins_fetch/add0/c53 ;
  wire \ins_fetch/add0/c54 ;
  wire \ins_fetch/add0/c55 ;
  wire \ins_fetch/add0/c56 ;
  wire \ins_fetch/add0/c57 ;
  wire \ins_fetch/add0/c58 ;
  wire \ins_fetch/add0/c59 ;
  wire \ins_fetch/add0/c6 ;
  wire \ins_fetch/add0/c60 ;
  wire \ins_fetch/add0/c61 ;
  wire \ins_fetch/add0/c7 ;
  wire \ins_fetch/add0/c8 ;
  wire \ins_fetch/add0/c9 ;
  wire \ins_fetch/addr_mis ;  // ../../RTL/CPU/IF/ins_fetch.v(57)
  wire \ins_fetch/hold ;  // ../../RTL/CPU/IF/ins_fetch.v(53)
  wire \ins_fetch/n25 ;
  wire \ins_fetch/n27 ;
  wire \ins_fetch/n9 ;
  wire ins_page_fault;  // ../../RTL/CPU/prv464_top.v(69)
  wire int_req;  // ../../RTL/CPU/prv464_top.v(259)
  wire jmp;  // ../../RTL/CPU/prv464_top.v(127)
  wire load;  // ../../RTL/CPU/prv464_top.v(136)
  wire load_acc_fault;  // ../../RTL/CPU/prv464_top.v(83)
  wire load_page_fault;  // ../../RTL/CPU/prv464_top.v(84)
  wire mem_csr_data_add;  // ../../RTL/CPU/prv464_top.v(116)
  wire mem_csr_data_and;  // ../../RTL/CPU/prv464_top.v(117)
  wire mem_csr_data_ds2;  // ../../RTL/CPU/prv464_top.v(115)
  wire mem_csr_data_max;  // ../../RTL/CPU/prv464_top.v(120)
  wire mem_csr_data_min;  // ../../RTL/CPU/prv464_top.v(121)
  wire mem_csr_data_or;  // ../../RTL/CPU/prv464_top.v(118)
  wire mem_csr_data_xor;  // ../../RTL/CPU/prv464_top.v(119)
  wire mprv;  // ../../RTL/CPU/prv464_top.v(53)
  wire mxr;  // ../../RTL/CPU/prv464_top.v(52)
  wire pc_jmp;  // ../../RTL/CPU/prv464_top.v(522)
  wire \pip_ctrl/eq2/xor_i0[1]_i1[1]_o_lutinv ;
  wire \pip_ctrl/ex_exception ;  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(80)
  wire \pip_ctrl/id_ex_war_lutinv ;  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(83)
  wire \pip_ctrl/id_exception ;  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(79)
  wire \pip_ctrl/n34 ;
  wire \pip_ctrl/n36_lutinv ;
  wire pip_flush;  // ../../RTL/CPU/prv464_top.v(265)
  wire rd_data_add;  // ../../RTL/CPU/prv464_top.v(104)
  wire rd_data_and;  // ../../RTL/CPU/prv464_top.v(106)
  wire rd_data_ds1;  // ../../RTL/CPU/prv464_top.v(103)
  wire rd_data_or;  // ../../RTL/CPU/prv464_top.v(107)
  wire rd_data_slt;  // ../../RTL/CPU/prv464_top.v(109)
  wire rd_data_sub;  // ../../RTL/CPU/prv464_top.v(105)
  wire rd_data_xor;  // ../../RTL/CPU/prv464_top.v(108)
  wire read;  // ../../RTL/CPU/prv464_top.v(81)
  wire rst_pad;  // ../../RTL/CPU/prv464_top.v(20)
  wire s_ext_int_pad;  // ../../RTL/CPU/prv464_top.v(40)
  wire shift_l;  // ../../RTL/CPU/prv464_top.v(142)
  wire shift_r;  // ../../RTL/CPU/prv464_top.v(141)
  wire store;  // ../../RTL/CPU/prv464_top.v(137)
  wire sum;  // ../../RTL/CPU/prv464_top.v(51)
  wire tsr;  // ../../RTL/CPU/prv464_top.v(50)
  wire tvm;  // ../../RTL/CPU/prv464_top.v(49)
  wire tw;  // ../../RTL/CPU/prv464_top.v(309)
  wire unsign;  // ../../RTL/CPU/prv464_top.v(128)
  wire wb_csr_write;  // ../../RTL/CPU/prv464_top.v(520)
  wire wb_ebreak;  // ../../RTL/CPU/prv464_top.v(547)
  wire wb_ecall;  // ../../RTL/CPU/prv464_top.v(546)
  wire wb_gpr_write;  // ../../RTL/CPU/prv464_top.v(521)
  wire wb_ill_ins;  // ../../RTL/CPU/prv464_top.v(543)
  wire wb_ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(532)
  wire wb_ins_addr_mis;  // ../../RTL/CPU/prv464_top.v(533)
  wire wb_ins_page_fault;  // ../../RTL/CPU/prv464_top.v(534)
  wire wb_int_acc;  // ../../RTL/CPU/prv464_top.v(541)
  wire wb_jmp;  // ../../RTL/CPU/prv464_top.v(531)
  wire wb_ld_acc_fault;  // ../../RTL/CPU/prv464_top.v(537)
  wire wb_ld_addr_mis;  // ../../RTL/CPU/prv464_top.v(535)
  wire wb_ld_page_fault;  // ../../RTL/CPU/prv464_top.v(539)
  wire wb_m_ret;  // ../../RTL/CPU/prv464_top.v(544)
  wire wb_s_ret;  // ../../RTL/CPU/prv464_top.v(545)
  wire wb_st_acc_fault;  // ../../RTL/CPU/prv464_top.v(538)
  wire wb_st_addr_mis;  // ../../RTL/CPU/prv464_top.v(536)
  wire wb_st_page_fault;  // ../../RTL/CPU/prv464_top.v(540)
  wire wb_system;  // ../../RTL/CPU/prv464_top.v(530)
  wire wb_valid;  // ../../RTL/CPU/prv464_top.v(542)
  wire write;  // ../../RTL/CPU/prv464_top.v(82)

  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1926 (
    .ipad(cacheability_block[31]),
    .di(cacheability_block_pad[31]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1927 (
    .ipad(cacheability_block[30]),
    .di(cacheability_block_pad[30]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1928 (
    .ipad(cacheability_block[29]),
    .di(cacheability_block_pad[29]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1929 (
    .ipad(cacheability_block[28]),
    .di(cacheability_block_pad[28]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1930 (
    .ipad(cacheability_block[27]),
    .di(cacheability_block_pad[27]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1931 (
    .ipad(cacheability_block[26]),
    .di(cacheability_block_pad[26]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1932 (
    .ipad(cacheability_block[25]),
    .di(cacheability_block_pad[25]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1933 (
    .ipad(cacheability_block[24]),
    .di(cacheability_block_pad[24]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1934 (
    .ipad(cacheability_block[23]),
    .di(cacheability_block_pad[23]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1935 (
    .ipad(cacheability_block[22]),
    .di(cacheability_block_pad[22]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1936 (
    .ipad(cacheability_block[21]),
    .di(cacheability_block_pad[21]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1937 (
    .ipad(cacheability_block[20]),
    .di(cacheability_block_pad[20]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1938 (
    .ipad(cacheability_block[19]),
    .di(cacheability_block_pad[19]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1939 (
    .ipad(cacheability_block[18]),
    .di(cacheability_block_pad[18]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1940 (
    .ipad(cacheability_block[17]),
    .di(cacheability_block_pad[17]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1941 (
    .ipad(cacheability_block[16]),
    .di(cacheability_block_pad[16]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1942 (
    .ipad(cacheability_block[15]),
    .di(cacheability_block_pad[15]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1943 (
    .ipad(cacheability_block[14]),
    .di(cacheability_block_pad[14]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1944 (
    .ipad(cacheability_block[13]),
    .di(cacheability_block_pad[13]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1945 (
    .ipad(cacheability_block[12]),
    .di(cacheability_block_pad[12]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1946 (
    .ipad(cacheability_block[11]),
    .di(cacheability_block_pad[11]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1947 (
    .ipad(cacheability_block[10]),
    .di(cacheability_block_pad[10]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1948 (
    .ipad(cacheability_block[9]),
    .di(cacheability_block_pad[9]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1949 (
    .ipad(cacheability_block[8]),
    .di(cacheability_block_pad[8]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1950 (
    .ipad(cacheability_block[7]),
    .di(cacheability_block_pad[7]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1951 (
    .ipad(cacheability_block[6]),
    .di(cacheability_block_pad[6]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1952 (
    .ipad(cacheability_block[5]),
    .di(cacheability_block_pad[5]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1953 (
    .ipad(cacheability_block[4]),
    .di(cacheability_block_pad[4]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1954 (
    .ipad(cacheability_block[3]),
    .di(cacheability_block_pad[3]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1955 (
    .ipad(cacheability_block[2]),
    .di(cacheability_block_pad[2]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1956 (
    .ipad(cacheability_block[1]),
    .di(cacheability_block_pad[1]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1957 (
    .ipad(cacheability_block[0]),
    .di(cacheability_block_pad[0]));  // ../../RTL/CPU/prv464_top.v(17)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u1958 (
    .ipad(clk),
    .di(clk_pad));  // ../../RTL/CPU/prv464_top.v(19)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1959 (
    .do({open_n562,open_n563,open_n564,haddr_pad[63]}),
    .opad(haddr[63]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1960 (
    .do({open_n579,open_n580,open_n581,haddr_pad[62]}),
    .opad(haddr[62]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1961 (
    .do({open_n596,open_n597,open_n598,haddr_pad[61]}),
    .opad(haddr[61]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1962 (
    .do({open_n613,open_n614,open_n615,haddr_pad[60]}),
    .opad(haddr[60]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1963 (
    .do({open_n630,open_n631,open_n632,haddr_pad[59]}),
    .opad(haddr[59]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1964 (
    .do({open_n647,open_n648,open_n649,haddr_pad[58]}),
    .opad(haddr[58]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1965 (
    .do({open_n664,open_n665,open_n666,haddr_pad[57]}),
    .opad(haddr[57]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1966 (
    .do({open_n681,open_n682,open_n683,haddr_pad[56]}),
    .opad(haddr[56]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1967 (
    .do({open_n698,open_n699,open_n700,haddr_pad[55]}),
    .opad(haddr[55]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1968 (
    .do({open_n715,open_n716,open_n717,haddr_pad[54]}),
    .opad(haddr[54]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1969 (
    .do({open_n732,open_n733,open_n734,haddr_pad[53]}),
    .opad(haddr[53]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1970 (
    .do({open_n749,open_n750,open_n751,haddr_pad[52]}),
    .opad(haddr[52]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1971 (
    .do({open_n766,open_n767,open_n768,haddr_pad[51]}),
    .opad(haddr[51]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1972 (
    .do({open_n783,open_n784,open_n785,haddr_pad[50]}),
    .opad(haddr[50]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1973 (
    .do({open_n800,open_n801,open_n802,haddr_pad[49]}),
    .opad(haddr[49]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1974 (
    .do({open_n817,open_n818,open_n819,haddr_pad[48]}),
    .opad(haddr[48]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1975 (
    .do({open_n834,open_n835,open_n836,haddr_pad[47]}),
    .opad(haddr[47]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1976 (
    .do({open_n851,open_n852,open_n853,haddr_pad[46]}),
    .opad(haddr[46]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1977 (
    .do({open_n868,open_n869,open_n870,haddr_pad[45]}),
    .opad(haddr[45]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1978 (
    .do({open_n885,open_n886,open_n887,haddr_pad[44]}),
    .opad(haddr[44]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1979 (
    .do({open_n902,open_n903,open_n904,haddr_pad[43]}),
    .opad(haddr[43]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1980 (
    .do({open_n919,open_n920,open_n921,haddr_pad[42]}),
    .opad(haddr[42]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1981 (
    .do({open_n936,open_n937,open_n938,haddr_pad[41]}),
    .opad(haddr[41]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1982 (
    .do({open_n953,open_n954,open_n955,haddr_pad[40]}),
    .opad(haddr[40]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1983 (
    .do({open_n970,open_n971,open_n972,haddr_pad[39]}),
    .opad(haddr[39]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1984 (
    .do({open_n987,open_n988,open_n989,haddr_pad[38]}),
    .opad(haddr[38]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1985 (
    .do({open_n1004,open_n1005,open_n1006,haddr_pad[37]}),
    .opad(haddr[37]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1986 (
    .do({open_n1021,open_n1022,open_n1023,haddr_pad[36]}),
    .opad(haddr[36]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1987 (
    .do({open_n1038,open_n1039,open_n1040,haddr_pad[35]}),
    .opad(haddr[35]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1988 (
    .do({open_n1055,open_n1056,open_n1057,haddr_pad[34]}),
    .opad(haddr[34]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1989 (
    .do({open_n1072,open_n1073,open_n1074,haddr_pad[33]}),
    .opad(haddr[33]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1990 (
    .do({open_n1089,open_n1090,open_n1091,haddr_pad[32]}),
    .opad(haddr[32]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1991 (
    .do({open_n1106,open_n1107,open_n1108,haddr_pad[31]}),
    .opad(haddr[31]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1992 (
    .do({open_n1123,open_n1124,open_n1125,haddr_pad[30]}),
    .opad(haddr[30]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1993 (
    .do({open_n1140,open_n1141,open_n1142,haddr_pad[29]}),
    .opad(haddr[29]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1994 (
    .do({open_n1157,open_n1158,open_n1159,haddr_pad[28]}),
    .opad(haddr[28]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1995 (
    .do({open_n1174,open_n1175,open_n1176,haddr_pad[27]}),
    .opad(haddr[27]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1996 (
    .do({open_n1191,open_n1192,open_n1193,haddr_pad[26]}),
    .opad(haddr[26]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1997 (
    .do({open_n1208,open_n1209,open_n1210,haddr_pad[25]}),
    .opad(haddr[25]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1998 (
    .do({open_n1225,open_n1226,open_n1227,haddr_pad[24]}),
    .opad(haddr[24]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u1999 (
    .do({open_n1242,open_n1243,open_n1244,haddr_pad[23]}),
    .opad(haddr[23]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2000 (
    .do({open_n1259,open_n1260,open_n1261,haddr_pad[22]}),
    .opad(haddr[22]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2001 (
    .do({open_n1276,open_n1277,open_n1278,haddr_pad[21]}),
    .opad(haddr[21]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2002 (
    .do({open_n1293,open_n1294,open_n1295,haddr_pad[20]}),
    .opad(haddr[20]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2003 (
    .do({open_n1310,open_n1311,open_n1312,haddr_pad[19]}),
    .opad(haddr[19]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2004 (
    .do({open_n1327,open_n1328,open_n1329,haddr_pad[18]}),
    .opad(haddr[18]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2005 (
    .do({open_n1344,open_n1345,open_n1346,haddr_pad[17]}),
    .opad(haddr[17]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2006 (
    .do({open_n1361,open_n1362,open_n1363,haddr_pad[16]}),
    .opad(haddr[16]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2007 (
    .do({open_n1378,open_n1379,open_n1380,haddr_pad[15]}),
    .opad(haddr[15]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2008 (
    .do({open_n1395,open_n1396,open_n1397,haddr_pad[14]}),
    .opad(haddr[14]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2009 (
    .do({open_n1412,open_n1413,open_n1414,haddr_pad[13]}),
    .opad(haddr[13]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2010 (
    .do({open_n1429,open_n1430,open_n1431,haddr_pad[12]}),
    .opad(haddr[12]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2011 (
    .do({open_n1446,open_n1447,open_n1448,haddr_pad[11]}),
    .opad(haddr[11]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2012 (
    .do({open_n1463,open_n1464,open_n1465,haddr_pad[10]}),
    .opad(haddr[10]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2013 (
    .do({open_n1480,open_n1481,open_n1482,haddr_pad[9]}),
    .opad(haddr[9]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2014 (
    .do({open_n1497,open_n1498,open_n1499,haddr_pad[8]}),
    .opad(haddr[8]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2015 (
    .do({open_n1514,open_n1515,open_n1516,haddr_pad[7]}),
    .opad(haddr[7]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2016 (
    .do({open_n1531,open_n1532,open_n1533,haddr_pad[6]}),
    .opad(haddr[6]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2017 (
    .do({open_n1548,open_n1549,open_n1550,haddr_pad[5]}),
    .opad(haddr[5]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2018 (
    .do({open_n1565,open_n1566,open_n1567,haddr_pad[4]}),
    .opad(haddr[4]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2019 (
    .do({open_n1582,open_n1583,open_n1584,haddr_pad[3]}),
    .opad(haddr[3]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2020 (
    .do({open_n1599,open_n1600,open_n1601,haddr_pad[2]}),
    .opad(haddr[2]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2021 (
    .do({open_n1616,open_n1617,open_n1618,haddr_pad[1]}),
    .opad(haddr[1]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2022 (
    .do({open_n1633,open_n1634,open_n1635,haddr_pad[0]}),
    .opad(haddr[0]));  // ../../RTL/CPU/prv464_top.v(22)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2023 (
    .do({open_n1650,open_n1651,open_n1652,1'b0}),
    .opad(hburst[2]));  // ../../RTL/CPU/prv464_top.v(25)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2024 (
    .do({open_n1667,open_n1668,open_n1669,1'b0}),
    .opad(hburst[1]));  // ../../RTL/CPU/prv464_top.v(25)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2025 (
    .do({open_n1684,open_n1685,open_n1686,hburst_pad[0]}),
    .opad(hburst[0]));  // ../../RTL/CPU/prv464_top.v(25)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2026 (
    .do({open_n1701,open_n1702,open_n1703,1'b0}),
    .opad(hmastlock));  // ../../RTL/CPU/prv464_top.v(28)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2027 (
    .do({open_n1718,open_n1719,open_n1720,1'b0}),
    .opad(hprot[3]));  // ../../RTL/CPU/prv464_top.v(26)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2028 (
    .do({open_n1735,open_n1736,open_n1737,1'b0}),
    .opad(hprot[2]));  // ../../RTL/CPU/prv464_top.v(26)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2029 (
    .do({open_n1752,open_n1753,open_n1754,1'b1}),
    .opad(hprot[1]));  // ../../RTL/CPU/prv464_top.v(26)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2030 (
    .do({open_n1769,open_n1770,open_n1771,1'b1}),
    .opad(hprot[0]));  // ../../RTL/CPU/prv464_top.v(26)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2031 (
    .ipad(hrdata[63]),
    .di(hrdata_pad[63]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2032 (
    .ipad(hrdata[62]),
    .di(hrdata_pad[62]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2033 (
    .ipad(hrdata[61]),
    .di(hrdata_pad[61]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2034 (
    .ipad(hrdata[60]),
    .di(hrdata_pad[60]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2035 (
    .ipad(hrdata[59]),
    .di(hrdata_pad[59]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2036 (
    .ipad(hrdata[58]),
    .di(hrdata_pad[58]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2037 (
    .ipad(hrdata[57]),
    .di(hrdata_pad[57]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2038 (
    .ipad(hrdata[56]),
    .di(hrdata_pad[56]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2039 (
    .ipad(hrdata[55]),
    .di(hrdata_pad[55]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2040 (
    .ipad(hrdata[54]),
    .di(hrdata_pad[54]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2041 (
    .ipad(hrdata[53]),
    .di(hrdata_pad[53]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2042 (
    .ipad(hrdata[52]),
    .di(hrdata_pad[52]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2043 (
    .ipad(hrdata[51]),
    .di(hrdata_pad[51]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2044 (
    .ipad(hrdata[50]),
    .di(hrdata_pad[50]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2045 (
    .ipad(hrdata[49]),
    .di(hrdata_pad[49]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2046 (
    .ipad(hrdata[48]),
    .di(hrdata_pad[48]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2047 (
    .ipad(hrdata[47]),
    .di(hrdata_pad[47]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2048 (
    .ipad(hrdata[46]),
    .di(hrdata_pad[46]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2049 (
    .ipad(hrdata[45]),
    .di(hrdata_pad[45]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2050 (
    .ipad(hrdata[44]),
    .di(hrdata_pad[44]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2051 (
    .ipad(hrdata[43]),
    .di(hrdata_pad[43]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2052 (
    .ipad(hrdata[42]),
    .di(hrdata_pad[42]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2053 (
    .ipad(hrdata[41]),
    .di(hrdata_pad[41]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2054 (
    .ipad(hrdata[40]),
    .di(hrdata_pad[40]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2055 (
    .ipad(hrdata[39]),
    .di(hrdata_pad[39]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2056 (
    .ipad(hrdata[38]),
    .di(hrdata_pad[38]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2057 (
    .ipad(hrdata[37]),
    .di(hrdata_pad[37]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2058 (
    .ipad(hrdata[36]),
    .di(hrdata_pad[36]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2059 (
    .ipad(hrdata[35]),
    .di(hrdata_pad[35]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2060 (
    .ipad(hrdata[34]),
    .di(hrdata_pad[34]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2061 (
    .ipad(hrdata[33]),
    .di(hrdata_pad[33]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2062 (
    .ipad(hrdata[32]),
    .di(hrdata_pad[32]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2063 (
    .ipad(hrdata[31]),
    .di(hrdata_pad[31]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2064 (
    .ipad(hrdata[30]),
    .di(hrdata_pad[30]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2065 (
    .ipad(hrdata[29]),
    .di(hrdata_pad[29]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2066 (
    .ipad(hrdata[28]),
    .di(hrdata_pad[28]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2067 (
    .ipad(hrdata[27]),
    .di(hrdata_pad[27]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2068 (
    .ipad(hrdata[26]),
    .di(hrdata_pad[26]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2069 (
    .ipad(hrdata[25]),
    .di(hrdata_pad[25]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2070 (
    .ipad(hrdata[24]),
    .di(hrdata_pad[24]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2071 (
    .ipad(hrdata[23]),
    .di(hrdata_pad[23]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2072 (
    .ipad(hrdata[22]),
    .di(hrdata_pad[22]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2073 (
    .ipad(hrdata[21]),
    .di(hrdata_pad[21]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2074 (
    .ipad(hrdata[20]),
    .di(hrdata_pad[20]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2075 (
    .ipad(hrdata[19]),
    .di(hrdata_pad[19]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2076 (
    .ipad(hrdata[18]),
    .di(hrdata_pad[18]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2077 (
    .ipad(hrdata[17]),
    .di(hrdata_pad[17]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2078 (
    .ipad(hrdata[16]),
    .di(hrdata_pad[16]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2079 (
    .ipad(hrdata[15]),
    .di(hrdata_pad[15]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2080 (
    .ipad(hrdata[14]),
    .di(hrdata_pad[14]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2081 (
    .ipad(hrdata[13]),
    .di(hrdata_pad[13]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2082 (
    .ipad(hrdata[12]),
    .di(hrdata_pad[12]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2083 (
    .ipad(hrdata[11]),
    .di(hrdata_pad[11]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2084 (
    .ipad(hrdata[10]),
    .di(hrdata_pad[10]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2085 (
    .ipad(hrdata[9]),
    .di(hrdata_pad[9]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2086 (
    .ipad(hrdata[8]),
    .di(hrdata_pad[8]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2087 (
    .ipad(hrdata[7]),
    .di(hrdata_pad[7]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2088 (
    .ipad(hrdata[6]),
    .di(hrdata_pad[6]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2089 (
    .ipad(hrdata[5]),
    .di(hrdata_pad[5]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2090 (
    .ipad(hrdata[4]),
    .di(hrdata_pad[4]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2091 (
    .ipad(hrdata[3]),
    .di(hrdata_pad[3]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2092 (
    .ipad(hrdata[2]),
    .di(hrdata_pad[2]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2093 (
    .ipad(hrdata[1]),
    .di(hrdata_pad[1]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2094 (
    .ipad(hrdata[0]),
    .di(hrdata_pad[0]));  // ../../RTL/CPU/prv464_top.v(34)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2095 (
    .ipad(hready),
    .di(hready_pad));  // ../../RTL/CPU/prv464_top.v(31)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2096 (
    .ipad(hreset_n));  // ../../RTL/CPU/prv464_top.v(33)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2097 (
    .ipad(hresp),
    .di(hresp_pad));  // ../../RTL/CPU/prv464_top.v(32)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2098 (
    .do({open_n2926,open_n2927,open_n2928,1'b0}),
    .opad(hsize[2]));  // ../../RTL/CPU/prv464_top.v(24)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2099 (
    .do({open_n2943,open_n2944,open_n2945,hsize_pad[1]}),
    .opad(hsize[1]));  // ../../RTL/CPU/prv464_top.v(24)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2100 (
    .do({open_n2960,open_n2961,open_n2962,hsize_pad[0]}),
    .opad(hsize[0]));  // ../../RTL/CPU/prv464_top.v(24)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2101 (
    .do({open_n2977,open_n2978,open_n2979,htrans_pad[1]}),
    .opad(htrans[1]));  // ../../RTL/CPU/prv464_top.v(27)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2102 (
    .do({open_n2994,open_n2995,open_n2996,htrans_pad[0]}),
    .opad(htrans[0]));  // ../../RTL/CPU/prv464_top.v(27)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2103 (
    .do({open_n3011,open_n3012,open_n3013,hwdata_pad[63]}),
    .opad(hwdata[63]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2104 (
    .do({open_n3028,open_n3029,open_n3030,hwdata_pad[62]}),
    .opad(hwdata[62]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2105 (
    .do({open_n3045,open_n3046,open_n3047,hwdata_pad[61]}),
    .opad(hwdata[61]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2106 (
    .do({open_n3062,open_n3063,open_n3064,hwdata_pad[60]}),
    .opad(hwdata[60]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2107 (
    .do({open_n3079,open_n3080,open_n3081,hwdata_pad[59]}),
    .opad(hwdata[59]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2108 (
    .do({open_n3096,open_n3097,open_n3098,hwdata_pad[58]}),
    .opad(hwdata[58]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2109 (
    .do({open_n3113,open_n3114,open_n3115,hwdata_pad[57]}),
    .opad(hwdata[57]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2110 (
    .do({open_n3130,open_n3131,open_n3132,hwdata_pad[56]}),
    .opad(hwdata[56]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2111 (
    .do({open_n3147,open_n3148,open_n3149,hwdata_pad[55]}),
    .opad(hwdata[55]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2112 (
    .do({open_n3164,open_n3165,open_n3166,hwdata_pad[54]}),
    .opad(hwdata[54]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2113 (
    .do({open_n3181,open_n3182,open_n3183,hwdata_pad[53]}),
    .opad(hwdata[53]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2114 (
    .do({open_n3198,open_n3199,open_n3200,hwdata_pad[52]}),
    .opad(hwdata[52]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2115 (
    .do({open_n3215,open_n3216,open_n3217,hwdata_pad[51]}),
    .opad(hwdata[51]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2116 (
    .do({open_n3232,open_n3233,open_n3234,hwdata_pad[50]}),
    .opad(hwdata[50]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2117 (
    .do({open_n3249,open_n3250,open_n3251,hwdata_pad[49]}),
    .opad(hwdata[49]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2118 (
    .do({open_n3266,open_n3267,open_n3268,hwdata_pad[48]}),
    .opad(hwdata[48]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2119 (
    .do({open_n3283,open_n3284,open_n3285,hwdata_pad[47]}),
    .opad(hwdata[47]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2120 (
    .do({open_n3300,open_n3301,open_n3302,hwdata_pad[46]}),
    .opad(hwdata[46]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2121 (
    .do({open_n3317,open_n3318,open_n3319,hwdata_pad[45]}),
    .opad(hwdata[45]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2122 (
    .do({open_n3334,open_n3335,open_n3336,hwdata_pad[44]}),
    .opad(hwdata[44]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2123 (
    .do({open_n3351,open_n3352,open_n3353,hwdata_pad[43]}),
    .opad(hwdata[43]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2124 (
    .do({open_n3368,open_n3369,open_n3370,hwdata_pad[42]}),
    .opad(hwdata[42]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2125 (
    .do({open_n3385,open_n3386,open_n3387,hwdata_pad[41]}),
    .opad(hwdata[41]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2126 (
    .do({open_n3402,open_n3403,open_n3404,hwdata_pad[40]}),
    .opad(hwdata[40]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2127 (
    .do({open_n3419,open_n3420,open_n3421,hwdata_pad[39]}),
    .opad(hwdata[39]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2128 (
    .do({open_n3436,open_n3437,open_n3438,hwdata_pad[38]}),
    .opad(hwdata[38]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2129 (
    .do({open_n3453,open_n3454,open_n3455,hwdata_pad[37]}),
    .opad(hwdata[37]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2130 (
    .do({open_n3470,open_n3471,open_n3472,hwdata_pad[36]}),
    .opad(hwdata[36]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2131 (
    .do({open_n3487,open_n3488,open_n3489,hwdata_pad[35]}),
    .opad(hwdata[35]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2132 (
    .do({open_n3504,open_n3505,open_n3506,hwdata_pad[34]}),
    .opad(hwdata[34]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2133 (
    .do({open_n3521,open_n3522,open_n3523,hwdata_pad[33]}),
    .opad(hwdata[33]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2134 (
    .do({open_n3538,open_n3539,open_n3540,hwdata_pad[32]}),
    .opad(hwdata[32]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2135 (
    .do({open_n3555,open_n3556,open_n3557,hwdata_pad[31]}),
    .opad(hwdata[31]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2136 (
    .do({open_n3572,open_n3573,open_n3574,hwdata_pad[30]}),
    .opad(hwdata[30]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2137 (
    .do({open_n3589,open_n3590,open_n3591,hwdata_pad[29]}),
    .opad(hwdata[29]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2138 (
    .do({open_n3606,open_n3607,open_n3608,hwdata_pad[28]}),
    .opad(hwdata[28]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2139 (
    .do({open_n3623,open_n3624,open_n3625,hwdata_pad[27]}),
    .opad(hwdata[27]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2140 (
    .do({open_n3640,open_n3641,open_n3642,hwdata_pad[26]}),
    .opad(hwdata[26]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2141 (
    .do({open_n3657,open_n3658,open_n3659,hwdata_pad[25]}),
    .opad(hwdata[25]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2142 (
    .do({open_n3674,open_n3675,open_n3676,hwdata_pad[24]}),
    .opad(hwdata[24]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2143 (
    .do({open_n3691,open_n3692,open_n3693,hwdata_pad[23]}),
    .opad(hwdata[23]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2144 (
    .do({open_n3708,open_n3709,open_n3710,hwdata_pad[22]}),
    .opad(hwdata[22]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2145 (
    .do({open_n3725,open_n3726,open_n3727,hwdata_pad[21]}),
    .opad(hwdata[21]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2146 (
    .do({open_n3742,open_n3743,open_n3744,hwdata_pad[20]}),
    .opad(hwdata[20]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2147 (
    .do({open_n3759,open_n3760,open_n3761,hwdata_pad[19]}),
    .opad(hwdata[19]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2148 (
    .do({open_n3776,open_n3777,open_n3778,hwdata_pad[18]}),
    .opad(hwdata[18]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2149 (
    .do({open_n3793,open_n3794,open_n3795,hwdata_pad[17]}),
    .opad(hwdata[17]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2150 (
    .do({open_n3810,open_n3811,open_n3812,hwdata_pad[16]}),
    .opad(hwdata[16]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2151 (
    .do({open_n3827,open_n3828,open_n3829,hwdata_pad[15]}),
    .opad(hwdata[15]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2152 (
    .do({open_n3844,open_n3845,open_n3846,hwdata_pad[14]}),
    .opad(hwdata[14]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2153 (
    .do({open_n3861,open_n3862,open_n3863,hwdata_pad[13]}),
    .opad(hwdata[13]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2154 (
    .do({open_n3878,open_n3879,open_n3880,hwdata_pad[12]}),
    .opad(hwdata[12]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2155 (
    .do({open_n3895,open_n3896,open_n3897,hwdata_pad[11]}),
    .opad(hwdata[11]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2156 (
    .do({open_n3912,open_n3913,open_n3914,hwdata_pad[10]}),
    .opad(hwdata[10]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2157 (
    .do({open_n3929,open_n3930,open_n3931,hwdata_pad[9]}),
    .opad(hwdata[9]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2158 (
    .do({open_n3946,open_n3947,open_n3948,hwdata_pad[8]}),
    .opad(hwdata[8]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2159 (
    .do({open_n3963,open_n3964,open_n3965,hwdata_pad[7]}),
    .opad(hwdata[7]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2160 (
    .do({open_n3980,open_n3981,open_n3982,hwdata_pad[6]}),
    .opad(hwdata[6]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2161 (
    .do({open_n3997,open_n3998,open_n3999,hwdata_pad[5]}),
    .opad(hwdata[5]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2162 (
    .do({open_n4014,open_n4015,open_n4016,hwdata_pad[4]}),
    .opad(hwdata[4]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2163 (
    .do({open_n4031,open_n4032,open_n4033,hwdata_pad[3]}),
    .opad(hwdata[3]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2164 (
    .do({open_n4048,open_n4049,open_n4050,hwdata_pad[2]}),
    .opad(hwdata[2]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2165 (
    .do({open_n4065,open_n4066,open_n4067,hwdata_pad[1]}),
    .opad(hwdata[1]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2166 (
    .do({open_n4082,open_n4083,open_n4084,hwdata_pad[0]}),
    .opad(hwdata[0]));  // ../../RTL/CPU/prv464_top.v(29)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u2167 (
    .do({open_n4099,open_n4100,open_n4101,hwrite_pad}),
    .opad(hwrite));  // ../../RTL/CPU/prv464_top.v(23)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2168 (
    .ipad(mtime[63]),
    .di(mtime_pad[63]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2169 (
    .ipad(mtime[62]),
    .di(mtime_pad[62]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2170 (
    .ipad(mtime[61]),
    .di(mtime_pad[61]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2171 (
    .ipad(mtime[60]),
    .di(mtime_pad[60]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2172 (
    .ipad(mtime[59]),
    .di(mtime_pad[59]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2173 (
    .ipad(mtime[58]),
    .di(mtime_pad[58]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2174 (
    .ipad(mtime[57]),
    .di(mtime_pad[57]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2175 (
    .ipad(mtime[56]),
    .di(mtime_pad[56]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2176 (
    .ipad(mtime[55]),
    .di(mtime_pad[55]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2177 (
    .ipad(mtime[54]),
    .di(mtime_pad[54]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2178 (
    .ipad(mtime[53]),
    .di(mtime_pad[53]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2179 (
    .ipad(mtime[52]),
    .di(mtime_pad[52]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2180 (
    .ipad(mtime[51]),
    .di(mtime_pad[51]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2181 (
    .ipad(mtime[50]),
    .di(mtime_pad[50]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2182 (
    .ipad(mtime[49]),
    .di(mtime_pad[49]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2183 (
    .ipad(mtime[48]),
    .di(mtime_pad[48]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2184 (
    .ipad(mtime[47]),
    .di(mtime_pad[47]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2185 (
    .ipad(mtime[46]),
    .di(mtime_pad[46]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2186 (
    .ipad(mtime[45]),
    .di(mtime_pad[45]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2187 (
    .ipad(mtime[44]),
    .di(mtime_pad[44]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2188 (
    .ipad(mtime[43]),
    .di(mtime_pad[43]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2189 (
    .ipad(mtime[42]),
    .di(mtime_pad[42]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2190 (
    .ipad(mtime[41]),
    .di(mtime_pad[41]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2191 (
    .ipad(mtime[40]),
    .di(mtime_pad[40]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2192 (
    .ipad(mtime[39]),
    .di(mtime_pad[39]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2193 (
    .ipad(mtime[38]),
    .di(mtime_pad[38]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2194 (
    .ipad(mtime[37]),
    .di(mtime_pad[37]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2195 (
    .ipad(mtime[36]),
    .di(mtime_pad[36]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2196 (
    .ipad(mtime[35]),
    .di(mtime_pad[35]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2197 (
    .ipad(mtime[34]),
    .di(mtime_pad[34]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2198 (
    .ipad(mtime[33]),
    .di(mtime_pad[33]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2199 (
    .ipad(mtime[32]),
    .di(mtime_pad[32]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2200 (
    .ipad(mtime[31]),
    .di(mtime_pad[31]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2201 (
    .ipad(mtime[30]),
    .di(mtime_pad[30]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2202 (
    .ipad(mtime[29]),
    .di(mtime_pad[29]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2203 (
    .ipad(mtime[28]),
    .di(mtime_pad[28]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2204 (
    .ipad(mtime[27]),
    .di(mtime_pad[27]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2205 (
    .ipad(mtime[26]),
    .di(mtime_pad[26]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2206 (
    .ipad(mtime[25]),
    .di(mtime_pad[25]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2207 (
    .ipad(mtime[24]),
    .di(mtime_pad[24]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2208 (
    .ipad(mtime[23]),
    .di(mtime_pad[23]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2209 (
    .ipad(mtime[22]),
    .di(mtime_pad[22]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2210 (
    .ipad(mtime[21]),
    .di(mtime_pad[21]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2211 (
    .ipad(mtime[20]),
    .di(mtime_pad[20]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2212 (
    .ipad(mtime[19]),
    .di(mtime_pad[19]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2213 (
    .ipad(mtime[18]),
    .di(mtime_pad[18]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2214 (
    .ipad(mtime[17]),
    .di(mtime_pad[17]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2215 (
    .ipad(mtime[16]),
    .di(mtime_pad[16]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2216 (
    .ipad(mtime[15]),
    .di(mtime_pad[15]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2217 (
    .ipad(mtime[14]),
    .di(mtime_pad[14]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2218 (
    .ipad(mtime[13]),
    .di(mtime_pad[13]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2219 (
    .ipad(mtime[12]),
    .di(mtime_pad[12]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2220 (
    .ipad(mtime[11]),
    .di(mtime_pad[11]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2221 (
    .ipad(mtime[10]),
    .di(mtime_pad[10]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2222 (
    .ipad(mtime[9]),
    .di(mtime_pad[9]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2223 (
    .ipad(mtime[8]),
    .di(mtime_pad[8]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2224 (
    .ipad(mtime[7]),
    .di(mtime_pad[7]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2225 (
    .ipad(mtime[6]),
    .di(mtime_pad[6]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2226 (
    .ipad(mtime[5]),
    .di(mtime_pad[5]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2227 (
    .ipad(mtime[4]),
    .di(mtime_pad[4]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2228 (
    .ipad(mtime[3]),
    .di(mtime_pad[3]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2229 (
    .ipad(mtime[2]),
    .di(mtime_pad[2]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2230 (
    .ipad(mtime[1]),
    .di(mtime_pad[1]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2231 (
    .ipad(mtime[0]),
    .di(mtime_pad[0]));  // ../../RTL/CPU/prv464_top.v(42)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2232 (
    .ipad(rst),
    .di(rst_pad));  // ../../RTL/CPU/prv464_top.v(20)
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u2233 (
    .ipad(s_ext_int),
    .di(s_ext_int_pad));  // ../../RTL/CPU/prv464_top.v(40)
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2558 (
    .a(s_ext_int_pad),
    .b(data_csr[9]),
    .o(\cu_ru/m_s_ip/n1 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2559 (
    .a(ins_read[9]),
    .b(ins_read[41]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [9]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2560 (
    .a(ins_read[8]),
    .b(ins_read[40]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2561 (
    .a(ins_read[7]),
    .b(ins_read[39]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2562 (
    .a(ins_read[6]),
    .b(ins_read[38]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2563 (
    .a(ins_read[5]),
    .b(ins_read[37]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2564 (
    .a(ins_read[4]),
    .b(ins_read[36]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2565 (
    .a(ins_read[31]),
    .b(ins_read[63]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2566 (
    .a(ins_read[30]),
    .b(ins_read[62]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2567 (
    .a(ins_read[3]),
    .b(ins_read[35]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2568 (
    .a(ins_read[29]),
    .b(ins_read[61]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2569 (
    .a(ins_read[28]),
    .b(ins_read[60]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2570 (
    .a(ins_read[27]),
    .b(ins_read[59]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2571 (
    .a(ins_read[26]),
    .b(ins_read[58]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2572 (
    .a(ins_read[25]),
    .b(ins_read[57]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2573 (
    .a(ins_read[24]),
    .b(ins_read[56]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2574 (
    .a(ins_read[23]),
    .b(ins_read[55]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2575 (
    .a(ins_read[22]),
    .b(ins_read[54]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2576 (
    .a(ins_read[21]),
    .b(ins_read[53]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2577 (
    .a(ins_read[20]),
    .b(ins_read[52]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2578 (
    .a(ins_read[2]),
    .b(ins_read[34]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2579 (
    .a(ins_read[19]),
    .b(ins_read[51]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2580 (
    .a(ins_read[18]),
    .b(ins_read[50]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2581 (
    .a(ins_read[17]),
    .b(ins_read[49]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2582 (
    .a(ins_read[16]),
    .b(ins_read[48]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2583 (
    .a(ins_read[15]),
    .b(ins_read[47]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2584 (
    .a(ins_read[14]),
    .b(ins_read[46]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2585 (
    .a(ins_read[13]),
    .b(ins_read[45]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2586 (
    .a(ins_read[12]),
    .b(ins_read[44]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2587 (
    .a(ins_read[11]),
    .b(ins_read[43]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2588 (
    .a(ins_read[10]),
    .b(ins_read[42]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2589 (
    .a(ins_read[1]),
    .b(ins_read[33]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u2590 (
    .a(ins_read[0]),
    .b(ins_read[32]),
    .c(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [0]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2591 (
    .a(addr_if[0]),
    .b(addr_if[1]),
    .o(\ins_fetch/addr_mis ));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2592 (
    .a(rd_data_sub),
    .b(ds2[0]),
    .o(\exu/alu_au/n17 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2593 (
    .a(rd_data_sub),
    .b(ds2[1]),
    .o(\exu/alu_au/n17 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2594 (
    .a(rd_data_sub),
    .b(ds2[10]),
    .o(\exu/alu_au/n17 [10]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2595 (
    .a(rd_data_sub),
    .b(ds2[11]),
    .o(\exu/alu_au/n17 [11]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2596 (
    .a(rd_data_sub),
    .b(ds2[12]),
    .o(\exu/alu_au/n17 [12]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2597 (
    .a(rd_data_sub),
    .b(ds2[13]),
    .o(\exu/alu_au/n17 [13]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2598 (
    .a(rd_data_sub),
    .b(ds2[14]),
    .o(\exu/alu_au/n17 [14]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2599 (
    .a(rd_data_sub),
    .b(ds2[15]),
    .o(\exu/alu_au/n17 [15]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2600 (
    .a(rd_data_sub),
    .b(ds2[16]),
    .o(\exu/alu_au/n17 [16]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2601 (
    .a(rd_data_sub),
    .b(ds2[17]),
    .o(\exu/alu_au/n17 [17]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2602 (
    .a(rd_data_sub),
    .b(ds2[18]),
    .o(\exu/alu_au/n17 [18]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2603 (
    .a(rd_data_sub),
    .b(ds2[19]),
    .o(\exu/alu_au/n17 [19]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2604 (
    .a(rd_data_sub),
    .b(ds2[2]),
    .o(\exu/alu_au/n17 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2605 (
    .a(rd_data_sub),
    .b(ds2[20]),
    .o(\exu/alu_au/n17 [20]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2606 (
    .a(rd_data_sub),
    .b(ds2[21]),
    .o(\exu/alu_au/n17 [21]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2607 (
    .a(rd_data_sub),
    .b(ds2[22]),
    .o(\exu/alu_au/n17 [22]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2608 (
    .a(rd_data_sub),
    .b(ds2[23]),
    .o(\exu/alu_au/n17 [23]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2609 (
    .a(rd_data_sub),
    .b(ds2[24]),
    .o(\exu/alu_au/n17 [24]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2610 (
    .a(rd_data_sub),
    .b(ds2[25]),
    .o(\exu/alu_au/n17 [25]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2611 (
    .a(rd_data_sub),
    .b(ds2[26]),
    .o(\exu/alu_au/n17 [26]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2612 (
    .a(rd_data_sub),
    .b(ds2[27]),
    .o(\exu/alu_au/n17 [27]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2613 (
    .a(rd_data_sub),
    .b(ds2[28]),
    .o(\exu/alu_au/n17 [28]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2614 (
    .a(rd_data_sub),
    .b(ds2[29]),
    .o(\exu/alu_au/n17 [29]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2615 (
    .a(rd_data_sub),
    .b(ds2[3]),
    .o(\exu/alu_au/n17 [3]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2616 (
    .a(rd_data_sub),
    .b(ds2[30]),
    .o(\exu/alu_au/n17 [30]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2617 (
    .a(rd_data_sub),
    .b(ds2[31]),
    .o(\exu/alu_au/n17 [31]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2618 (
    .a(rd_data_sub),
    .b(ds2[32]),
    .o(\exu/alu_au/n17 [32]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2619 (
    .a(rd_data_sub),
    .b(ds2[33]),
    .o(\exu/alu_au/n17 [33]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2620 (
    .a(rd_data_sub),
    .b(ds2[34]),
    .o(\exu/alu_au/n17 [34]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2621 (
    .a(rd_data_sub),
    .b(ds2[35]),
    .o(\exu/alu_au/n17 [35]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2622 (
    .a(rd_data_sub),
    .b(ds2[36]),
    .o(\exu/alu_au/n17 [36]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2623 (
    .a(rd_data_sub),
    .b(ds2[37]),
    .o(\exu/alu_au/n17 [37]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2624 (
    .a(rd_data_sub),
    .b(ds2[38]),
    .o(\exu/alu_au/n17 [38]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2625 (
    .a(rd_data_sub),
    .b(ds2[39]),
    .o(\exu/alu_au/n17 [39]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2626 (
    .a(rd_data_sub),
    .b(ds2[4]),
    .o(\exu/alu_au/n17 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2627 (
    .a(rd_data_sub),
    .b(ds2[40]),
    .o(\exu/alu_au/n17 [40]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2628 (
    .a(rd_data_sub),
    .b(ds2[41]),
    .o(\exu/alu_au/n17 [41]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2629 (
    .a(rd_data_sub),
    .b(ds2[42]),
    .o(\exu/alu_au/n17 [42]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2630 (
    .a(rd_data_sub),
    .b(ds2[43]),
    .o(\exu/alu_au/n17 [43]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2631 (
    .a(rd_data_sub),
    .b(ds2[44]),
    .o(\exu/alu_au/n17 [44]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2632 (
    .a(rd_data_sub),
    .b(ds2[45]),
    .o(\exu/alu_au/n17 [45]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2633 (
    .a(rd_data_sub),
    .b(ds2[46]),
    .o(\exu/alu_au/n17 [46]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2634 (
    .a(rd_data_sub),
    .b(ds2[47]),
    .o(\exu/alu_au/n17 [47]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2635 (
    .a(rd_data_sub),
    .b(ds2[48]),
    .o(\exu/alu_au/n17 [48]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2636 (
    .a(rd_data_sub),
    .b(ds2[49]),
    .o(\exu/alu_au/n17 [49]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2637 (
    .a(rd_data_sub),
    .b(ds2[5]),
    .o(\exu/alu_au/n17 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2638 (
    .a(rd_data_sub),
    .b(ds2[50]),
    .o(\exu/alu_au/n17 [50]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2639 (
    .a(rd_data_sub),
    .b(ds2[51]),
    .o(\exu/alu_au/n17 [51]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2640 (
    .a(rd_data_sub),
    .b(ds2[52]),
    .o(\exu/alu_au/n17 [52]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2641 (
    .a(rd_data_sub),
    .b(ds2[53]),
    .o(\exu/alu_au/n17 [53]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2642 (
    .a(rd_data_sub),
    .b(ds2[54]),
    .o(\exu/alu_au/n17 [54]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2643 (
    .a(rd_data_sub),
    .b(ds2[55]),
    .o(\exu/alu_au/n17 [55]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2644 (
    .a(rd_data_sub),
    .b(ds2[56]),
    .o(\exu/alu_au/n17 [56]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2645 (
    .a(rd_data_sub),
    .b(ds2[57]),
    .o(\exu/alu_au/n17 [57]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2646 (
    .a(rd_data_sub),
    .b(ds2[58]),
    .o(\exu/alu_au/n17 [58]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2647 (
    .a(rd_data_sub),
    .b(ds2[59]),
    .o(\exu/alu_au/n17 [59]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2648 (
    .a(rd_data_sub),
    .b(ds2[6]),
    .o(\exu/alu_au/n17 [6]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2649 (
    .a(rd_data_sub),
    .b(ds2[60]),
    .o(\exu/alu_au/n17 [60]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2650 (
    .a(rd_data_sub),
    .b(ds2[61]),
    .o(\exu/alu_au/n17 [61]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2651 (
    .a(rd_data_sub),
    .b(ds2[62]),
    .o(\exu/alu_au/n17 [62]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2652 (
    .a(rd_data_sub),
    .b(ds2[63]),
    .o(\exu/alu_au/n17 [63]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2653 (
    .a(rd_data_sub),
    .b(ds2[7]),
    .o(\exu/alu_au/n17 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2654 (
    .a(rd_data_sub),
    .b(ds2[8]),
    .o(\exu/alu_au/n17 [8]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u2655 (
    .a(rd_data_sub),
    .b(ds2[9]),
    .o(\exu/alu_au/n17 [9]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u2656 (
    .a(\ins_fetch/ins_shift [9]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [9]),
    .o(id_ins[9]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u2657 (
    .a(\ins_fetch/ins_shift [8]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [8]),
    .o(id_ins[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u2658 (
    .a(\ins_fetch/ins_shift [7]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [7]),
    .o(id_ins[7]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2659 (
    .a(ins_read[31]),
    .b(ins_read[63]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2659_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2660 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [31]),
    .o(_al_u2660_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2661 (
    .a(_al_u2659_o),
    .b(_al_u2660_o),
    .o(id_ins[31]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2662 (
    .a(ins_read[30]),
    .b(ins_read[62]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2662_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2663 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [30]),
    .o(_al_u2663_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2664 (
    .a(_al_u2662_o),
    .b(_al_u2663_o),
    .o(id_ins[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u2665 (
    .a(\ins_fetch/ins_shift [29]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [29]),
    .o(id_ins[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u2666 (
    .a(\ins_fetch/ins_shift [28]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [28]),
    .o(id_ins[28]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2667 (
    .a(ins_read[27]),
    .b(ins_read[59]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2667_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2668 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [27]),
    .o(_al_u2668_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2669 (
    .a(_al_u2667_o),
    .b(_al_u2668_o),
    .o(id_ins[27]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2670 (
    .a(ins_read[26]),
    .b(ins_read[58]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2670_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2671 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [26]),
    .o(_al_u2671_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2672 (
    .a(_al_u2670_o),
    .b(_al_u2671_o),
    .o(id_ins[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u2673 (
    .a(\ins_fetch/ins_shift [25]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [25]),
    .o(id_ins[25]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2674 (
    .a(ins_read[24]),
    .b(ins_read[56]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2674_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2675 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [24]),
    .o(_al_u2675_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2676 (
    .a(_al_u2674_o),
    .b(_al_u2675_o),
    .o(id_ins[24]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2677 (
    .a(ins_read[23]),
    .b(ins_read[55]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2677_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2678 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [23]),
    .o(_al_u2678_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2679 (
    .a(_al_u2677_o),
    .b(_al_u2678_o),
    .o(id_ins[23]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2680 (
    .a(ins_read[22]),
    .b(ins_read[54]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2680_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2681 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [22]),
    .o(_al_u2681_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2682 (
    .a(_al_u2680_o),
    .b(_al_u2681_o),
    .o(id_ins[22]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2683 (
    .a(ins_read[21]),
    .b(ins_read[53]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2683_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2684 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [21]),
    .o(_al_u2684_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2685 (
    .a(_al_u2683_o),
    .b(_al_u2684_o),
    .o(id_ins[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u2686 (
    .a(\ins_fetch/ins_shift [20]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [20]),
    .o(id_ins[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u2687 (
    .a(\ins_fetch/ins_shift [11]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [11]),
    .o(id_ins[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u2688 (
    .a(\ins_fetch/ins_shift [10]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [10]),
    .o(id_ins[10]));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u2689 (
    .a(rst_pad),
    .b(id_valid),
    .o(\ins_dec/n107 ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u2690 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .o(\biu/bus_unit/mmu/n59 [1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2691 (
    .a(wb_rd_index[2]),
    .b(wb_rd_index[3]),
    .c(wb_rd_index[4]),
    .o(_al_u2691_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u2692 (
    .a(_al_u2691_o),
    .b(wb_gpr_write),
    .c(wb_rd_index[0]),
    .d(wb_rd_index[1]),
    .o(\cu_ru/n53_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2693 (
    .a(\cu_ru/n53_lutinv ),
    .b(\cu_ru/n52 [4]),
    .o(\cu_ru/n53_1_al_n1986 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2694 (
    .a(\cu_ru/n53_lutinv ),
    .b(\cu_ru/n52 [4]),
    .o(\cu_ru/n53_0_al_n1985 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2695 (
    .a(id_ins_acc_fault),
    .b(id_ins_addr_mis),
    .c(id_ins_page_fault),
    .o(_al_u2695_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u2696 (
    .a(_al_u2695_o),
    .b(rst_pad),
    .o(\ins_fetch/n25 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2697 (
    .a(\biu/bus_unit/mmu/statu [1]),
    .b(\biu/bus_unit/mmu/statu [2]),
    .c(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u2697_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2698 (
    .a(_al_u2697_o),
    .b(\biu/bus_unit/mmu/statu [0]),
    .o(_al_u2698_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2699 (
    .a(_al_u2698_o),
    .b(rst_pad),
    .o(\biu/bus_unit/mmu/n58 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2700 (
    .a(\biu/bus_unit/mmu/statu [0]),
    .b(\biu/bus_unit/mmu/statu [1]),
    .c(\biu/bus_unit/mmu/statu [2]),
    .d(\biu/bus_unit/mmu/statu [3]),
    .o(\biu/bus_unit/mmu/n37_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2701 (
    .a(\biu/bus_unit/mmu_hwdata [1]),
    .b(\biu/bus_unit/mmu_hwdata [3]),
    .o(\biu/bus_unit/mmu/n39 [0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2702 (
    .a(\biu/bus_unit/mmu/n37_lutinv ),
    .b(\biu/bus_unit/mmu/n39 [0]),
    .c(\biu/bus_unit/mmu_hwdata [2]),
    .o(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2703 (
    .a(\biu/bus_unit/statu [2]),
    .b(\biu/bus_unit/statu [4]),
    .o(_al_u2703_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2704 (
    .a(_al_u2703_o),
    .b(\biu/bus_unit/statu [1]),
    .c(\biu/bus_unit/statu [3]),
    .o(_al_u2704_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2705 (
    .a(_al_u2704_o),
    .b(\biu/bus_unit/statu [0]),
    .o(_al_u2705_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u2706 (
    .a(_al_u2703_o),
    .b(\biu/bus_unit/statu [0]),
    .c(\biu/bus_unit/statu [1]),
    .d(\biu/bus_unit/statu [3]),
    .o(_al_u2706_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u2707 (
    .a(\biu/bus_unit/mmu/statu [0]),
    .b(\biu/bus_unit/mmu/statu [1]),
    .c(\biu/bus_unit/mmu/statu [2]),
    .d(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u2707_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u2708 (
    .a(_al_u2705_o),
    .b(_al_u2706_o),
    .c(_al_u2707_o),
    .o(hwrite_pad));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2709 (
    .a(_al_u2705_o),
    .b(hrdata_pad[9]),
    .o(uncache_data[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2710 (
    .a(_al_u2705_o),
    .b(hrdata_pad[8]),
    .o(uncache_data[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2711 (
    .a(_al_u2705_o),
    .b(hrdata_pad[63]),
    .o(uncache_data[63]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2712 (
    .a(_al_u2705_o),
    .b(hrdata_pad[62]),
    .o(uncache_data[62]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2713 (
    .a(_al_u2705_o),
    .b(hrdata_pad[61]),
    .o(uncache_data[61]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2714 (
    .a(_al_u2705_o),
    .b(hrdata_pad[60]),
    .o(uncache_data[60]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2715 (
    .a(_al_u2705_o),
    .b(hrdata_pad[6]),
    .o(uncache_data[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2716 (
    .a(_al_u2705_o),
    .b(hrdata_pad[59]),
    .o(uncache_data[59]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2717 (
    .a(_al_u2705_o),
    .b(hrdata_pad[58]),
    .o(uncache_data[58]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2718 (
    .a(_al_u2705_o),
    .b(hrdata_pad[57]),
    .o(uncache_data[57]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2719 (
    .a(_al_u2705_o),
    .b(hrdata_pad[56]),
    .o(uncache_data[56]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2720 (
    .a(_al_u2705_o),
    .b(hrdata_pad[55]),
    .o(uncache_data[55]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2721 (
    .a(_al_u2705_o),
    .b(hrdata_pad[54]),
    .o(uncache_data[54]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2722 (
    .a(_al_u2705_o),
    .b(hrdata_pad[53]),
    .o(uncache_data[53]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2723 (
    .a(_al_u2705_o),
    .b(hrdata_pad[52]),
    .o(uncache_data[52]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2724 (
    .a(_al_u2705_o),
    .b(hrdata_pad[51]),
    .o(uncache_data[51]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2725 (
    .a(_al_u2705_o),
    .b(hrdata_pad[50]),
    .o(uncache_data[50]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2726 (
    .a(_al_u2705_o),
    .b(hrdata_pad[5]),
    .o(uncache_data[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2727 (
    .a(_al_u2705_o),
    .b(hrdata_pad[49]),
    .o(uncache_data[49]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2728 (
    .a(_al_u2705_o),
    .b(hrdata_pad[48]),
    .o(uncache_data[48]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2729 (
    .a(_al_u2705_o),
    .b(hrdata_pad[47]),
    .o(uncache_data[47]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2730 (
    .a(_al_u2705_o),
    .b(hrdata_pad[46]),
    .o(uncache_data[46]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2731 (
    .a(_al_u2705_o),
    .b(hrdata_pad[45]),
    .o(uncache_data[45]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2732 (
    .a(_al_u2705_o),
    .b(hrdata_pad[44]),
    .o(uncache_data[44]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2733 (
    .a(_al_u2705_o),
    .b(hrdata_pad[43]),
    .o(uncache_data[43]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2734 (
    .a(_al_u2705_o),
    .b(hrdata_pad[42]),
    .o(uncache_data[42]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2735 (
    .a(_al_u2705_o),
    .b(hrdata_pad[41]),
    .o(uncache_data[41]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2736 (
    .a(_al_u2705_o),
    .b(hrdata_pad[40]),
    .o(uncache_data[40]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2737 (
    .a(_al_u2705_o),
    .b(hrdata_pad[4]),
    .o(uncache_data[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2738 (
    .a(_al_u2705_o),
    .b(hrdata_pad[39]),
    .o(uncache_data[39]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2739 (
    .a(_al_u2705_o),
    .b(hrdata_pad[38]),
    .o(uncache_data[38]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2740 (
    .a(_al_u2705_o),
    .b(hrdata_pad[37]),
    .o(uncache_data[37]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2741 (
    .a(_al_u2705_o),
    .b(hrdata_pad[36]),
    .o(uncache_data[36]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2742 (
    .a(_al_u2705_o),
    .b(hrdata_pad[35]),
    .o(uncache_data[35]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2743 (
    .a(_al_u2705_o),
    .b(hrdata_pad[34]),
    .o(uncache_data[34]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2744 (
    .a(_al_u2705_o),
    .b(hrdata_pad[33]),
    .o(uncache_data[33]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2745 (
    .a(_al_u2705_o),
    .b(hrdata_pad[32]),
    .o(uncache_data[32]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2746 (
    .a(_al_u2705_o),
    .b(hrdata_pad[31]),
    .o(uncache_data[31]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2747 (
    .a(_al_u2705_o),
    .b(hrdata_pad[30]),
    .o(uncache_data[30]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2748 (
    .a(_al_u2705_o),
    .b(hrdata_pad[3]),
    .o(uncache_data[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2749 (
    .a(_al_u2705_o),
    .b(hrdata_pad[29]),
    .o(uncache_data[29]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2750 (
    .a(_al_u2705_o),
    .b(hrdata_pad[28]),
    .o(uncache_data[28]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2751 (
    .a(_al_u2705_o),
    .b(hrdata_pad[27]),
    .o(uncache_data[27]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2752 (
    .a(_al_u2705_o),
    .b(hrdata_pad[26]),
    .o(uncache_data[26]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2753 (
    .a(_al_u2705_o),
    .b(hrdata_pad[25]),
    .o(uncache_data[25]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2754 (
    .a(_al_u2705_o),
    .b(hrdata_pad[24]),
    .o(uncache_data[24]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2755 (
    .a(_al_u2705_o),
    .b(hrdata_pad[23]),
    .o(uncache_data[23]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2756 (
    .a(_al_u2705_o),
    .b(hrdata_pad[22]),
    .o(uncache_data[22]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2757 (
    .a(_al_u2705_o),
    .b(hrdata_pad[21]),
    .o(uncache_data[21]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2758 (
    .a(_al_u2705_o),
    .b(hrdata_pad[20]),
    .o(uncache_data[20]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2759 (
    .a(_al_u2705_o),
    .b(hrdata_pad[2]),
    .o(uncache_data[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2760 (
    .a(_al_u2705_o),
    .b(hrdata_pad[19]),
    .o(uncache_data[19]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2761 (
    .a(_al_u2705_o),
    .b(hrdata_pad[18]),
    .o(uncache_data[18]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2762 (
    .a(_al_u2705_o),
    .b(hrdata_pad[17]),
    .o(uncache_data[17]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2763 (
    .a(_al_u2705_o),
    .b(hrdata_pad[16]),
    .o(uncache_data[16]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2764 (
    .a(_al_u2705_o),
    .b(hrdata_pad[15]),
    .o(uncache_data[15]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2765 (
    .a(_al_u2705_o),
    .b(hrdata_pad[14]),
    .o(uncache_data[14]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2766 (
    .a(_al_u2705_o),
    .b(hrdata_pad[13]),
    .o(uncache_data[13]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2767 (
    .a(_al_u2705_o),
    .b(hrdata_pad[12]),
    .o(uncache_data[12]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2768 (
    .a(_al_u2705_o),
    .b(hrdata_pad[11]),
    .o(uncache_data[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2769 (
    .a(_al_u2705_o),
    .b(hrdata_pad[10]),
    .o(uncache_data[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2770 (
    .a(_al_u2705_o),
    .b(hrdata_pad[1]),
    .o(uncache_data[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2771 (
    .a(_al_u2705_o),
    .b(hrdata_pad[0]),
    .c(\biu/bus_unit/mmu_hwdata [0]),
    .o(uncache_data[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2772 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [6]),
    .c(\biu/paddress [73]),
    .o(haddr_pad[9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2773 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [5]),
    .c(\biu/paddress [72]),
    .o(haddr_pad[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2774 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [4]),
    .c(\biu/paddress [71]),
    .o(haddr_pad[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2775 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [60]),
    .c(\biu/paddress [127]),
    .o(haddr_pad[63]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2776 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [59]),
    .c(\biu/paddress [126]),
    .o(haddr_pad[62]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2777 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [58]),
    .c(\biu/paddress [125]),
    .o(haddr_pad[61]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2778 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [57]),
    .c(\biu/paddress [124]),
    .o(haddr_pad[60]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2779 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [3]),
    .c(\biu/paddress [70]),
    .o(haddr_pad[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2780 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [56]),
    .c(\biu/paddress [123]),
    .o(haddr_pad[59]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2781 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [55]),
    .c(\biu/paddress [122]),
    .o(haddr_pad[58]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2782 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [54]),
    .c(\biu/paddress [121]),
    .o(haddr_pad[57]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2783 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [53]),
    .c(\biu/paddress [120]),
    .o(haddr_pad[56]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2784 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [52]),
    .c(\biu/paddress [119]),
    .o(haddr_pad[55]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2785 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [51]),
    .c(\biu/paddress [118]),
    .o(haddr_pad[54]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2786 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [50]),
    .c(\biu/paddress [117]),
    .o(haddr_pad[53]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2787 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [49]),
    .c(\biu/paddress [116]),
    .o(haddr_pad[52]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2788 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [48]),
    .c(\biu/paddress [115]),
    .o(haddr_pad[51]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2789 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [47]),
    .c(\biu/paddress [114]),
    .o(haddr_pad[50]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2790 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [2]),
    .c(\biu/paddress [69]),
    .o(haddr_pad[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2791 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [46]),
    .c(\biu/paddress [113]),
    .o(haddr_pad[49]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2792 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [45]),
    .c(\biu/paddress [112]),
    .o(haddr_pad[48]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2793 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [44]),
    .c(\biu/paddress [111]),
    .o(haddr_pad[47]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2794 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [43]),
    .c(\biu/paddress [110]),
    .o(haddr_pad[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2795 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [42]),
    .c(\biu/paddress [109]),
    .o(haddr_pad[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2796 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [41]),
    .c(\biu/paddress [108]),
    .o(haddr_pad[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2797 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [40]),
    .c(\biu/paddress [107]),
    .o(haddr_pad[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2798 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [39]),
    .c(\biu/paddress [106]),
    .o(haddr_pad[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2799 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [38]),
    .c(\biu/paddress [105]),
    .o(haddr_pad[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2800 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [37]),
    .c(\biu/paddress [104]),
    .o(haddr_pad[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2801 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [1]),
    .c(\biu/paddress [68]),
    .o(haddr_pad[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2802 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [36]),
    .c(\biu/paddress [103]),
    .o(haddr_pad[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2803 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [35]),
    .c(\biu/paddress [102]),
    .o(haddr_pad[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2804 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [34]),
    .c(\biu/paddress [101]),
    .o(haddr_pad[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2805 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [33]),
    .c(\biu/paddress [100]),
    .o(haddr_pad[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2806 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [32]),
    .c(\biu/paddress [99]),
    .o(haddr_pad[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2807 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [31]),
    .c(\biu/paddress [98]),
    .o(haddr_pad[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2808 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [30]),
    .c(\biu/paddress [97]),
    .o(haddr_pad[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2809 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [29]),
    .c(\biu/paddress [96]),
    .o(haddr_pad[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2810 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [28]),
    .c(\biu/paddress [95]),
    .o(haddr_pad[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2811 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [27]),
    .c(\biu/paddress [94]),
    .o(haddr_pad[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2812 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [0]),
    .c(\biu/paddress [67]),
    .o(haddr_pad[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2813 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [26]),
    .c(\biu/paddress [93]),
    .o(haddr_pad[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2814 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [25]),
    .c(\biu/paddress [92]),
    .o(haddr_pad[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2815 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [24]),
    .c(\biu/paddress [91]),
    .o(haddr_pad[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2816 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [23]),
    .c(\biu/paddress [90]),
    .o(haddr_pad[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2817 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [22]),
    .c(\biu/paddress [89]),
    .o(haddr_pad[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2818 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [21]),
    .c(\biu/paddress [88]),
    .o(haddr_pad[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2819 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [20]),
    .c(\biu/paddress [87]),
    .o(haddr_pad[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2820 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [19]),
    .c(\biu/paddress [86]),
    .o(haddr_pad[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2821 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [18]),
    .c(\biu/paddress [85]),
    .o(haddr_pad[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2822 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [17]),
    .c(\biu/paddress [84]),
    .o(haddr_pad[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2823 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [16]),
    .c(\biu/paddress [83]),
    .o(haddr_pad[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2824 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [15]),
    .c(\biu/paddress [82]),
    .o(haddr_pad[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2825 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [14]),
    .c(\biu/paddress [81]),
    .o(haddr_pad[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2826 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [13]),
    .c(\biu/paddress [80]),
    .o(haddr_pad[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2827 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [12]),
    .c(\biu/paddress [79]),
    .o(haddr_pad[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2828 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [11]),
    .c(\biu/paddress [78]),
    .o(haddr_pad[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2829 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [10]),
    .c(\biu/paddress [77]),
    .o(haddr_pad[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2830 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [9]),
    .c(\biu/paddress [76]),
    .o(haddr_pad[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2831 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [8]),
    .c(\biu/paddress [75]),
    .o(haddr_pad[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2832 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/n49 [7]),
    .c(\biu/paddress [74]),
    .o(haddr_pad[10]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2833 (
    .a(_al_u2704_o),
    .b(\biu/bus_unit/statu [0]),
    .o(_al_u2833_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2834 (
    .a(_al_u2833_o),
    .b(rst_pad),
    .o(\biu/bus_unit/n37 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2835 (
    .a(\biu/cache_ctrl_logic/statu [2]),
    .b(\biu/cache_ctrl_logic/statu [3]),
    .c(\biu/cache_ctrl_logic/statu [4]),
    .o(_al_u2835_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u2836 (
    .a(_al_u2835_o),
    .b(\biu/cache_ctrl_logic/statu [0]),
    .c(\biu/cache_ctrl_logic/statu [1]),
    .o(load_acc_fault));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2837 (
    .a(\biu/cache_ctrl_logic/statu [0]),
    .b(\biu/cache_ctrl_logic/statu [1]),
    .o(_al_u2837_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u2838 (
    .a(\biu/cache_ctrl_logic/statu [2]),
    .b(\biu/cache_ctrl_logic/statu [3]),
    .c(\biu/cache_ctrl_logic/statu [4]),
    .o(_al_u2838_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2839 (
    .a(_al_u2837_o),
    .b(_al_u2838_o),
    .o(ins_acc_fault));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2840 (
    .a(wb_m_ret),
    .b(wb_valid),
    .o(\cu_ru/m_s_status/n2 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2841 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mstatus [11]),
    .o(_al_u2841_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u2842 (
    .a(wb_m_ret),
    .b(wb_s_ret),
    .c(wb_valid),
    .o(_al_u2842_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~B)*~(C*A))"),
    .INIT(16'hb3a0))
    _al_u2843 (
    .a(_al_u2841_o),
    .b(_al_u2842_o),
    .c(\cu_ru/mstatus [12]),
    .d(priv[3]),
    .o(\cu_ru/m_s_status/n64 [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2844 (
    .a(wb_s_ret),
    .b(wb_valid),
    .o(_al_u2844_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u2845 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(priv[1]),
    .d(\cu_ru/mstatus [8]),
    .o(_al_u2845_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(~C*A))"),
    .INIT(8'hce))
    _al_u2846 (
    .a(_al_u2841_o),
    .b(_al_u2845_o),
    .c(\cu_ru/mstatus [12]),
    .o(\cu_ru/m_s_status/n64 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2847 (
    .a(\biu/cache_ctrl_logic/statu [0]),
    .b(\biu/cache_ctrl_logic/statu [1]),
    .o(_al_u2847_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u2848 (
    .a(_al_u2847_o),
    .b(\biu/cache_ctrl_logic/statu [2]),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(_al_u2848_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2849 (
    .a(_al_u2848_o),
    .b(rst_pad),
    .o(\biu/cache_ctrl_logic/u128_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(~A*(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B))"),
    .INIT(16'h4501))
    _al_u2850 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(priv[0]),
    .d(\cu_ru/mstatus [8]),
    .o(_al_u2850_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2851 (
    .a(_al_u2841_o),
    .b(_al_u2850_o),
    .o(\cu_ru/m_s_status/n64 [0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2852 (
    .a(shift_l),
    .b(shift_r),
    .o(_al_u2852_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2853 (
    .a(\exu/main_state [0]),
    .b(\exu/main_state [1]),
    .c(\exu/main_state [2]),
    .d(\exu/main_state [3]),
    .o(\exu/c_stb_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u2854 (
    .a(_al_u2852_o),
    .b(\exu/c_stb_lutinv ),
    .c(ex_valid),
    .o(\exu/n49 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u2855 (
    .a(\exu/main_state [0]),
    .b(\exu/main_state [1]),
    .c(\exu/main_state [2]),
    .d(\exu/main_state [3]),
    .o(_al_u2855_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u2856 (
    .a(_al_u2855_o),
    .b(\exu/shift_count [7]),
    .c(\exu/n50 [7]),
    .o(_al_u2856_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u2857 (
    .a(\exu/n49 ),
    .b(_al_u2856_o),
    .c(op_count[7]),
    .o(\exu/n52 [7]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u2858 (
    .a(_al_u2855_o),
    .b(\exu/shift_count [6]),
    .c(\exu/n50 [6]),
    .o(_al_u2858_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u2859 (
    .a(\exu/n49 ),
    .b(_al_u2858_o),
    .c(op_count[6]),
    .o(\exu/n52 [6]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u2860 (
    .a(_al_u2855_o),
    .b(\exu/shift_count [5]),
    .c(\exu/n50 [5]),
    .o(_al_u2860_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u2861 (
    .a(\exu/n49 ),
    .b(_al_u2860_o),
    .c(op_count[5]),
    .o(\exu/n52 [5]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u2862 (
    .a(_al_u2855_o),
    .b(\exu/shift_count [4]),
    .c(\exu/n50 [4]),
    .o(_al_u2862_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u2863 (
    .a(\exu/n49 ),
    .b(_al_u2862_o),
    .c(op_count[4]),
    .o(\exu/n52 [4]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u2864 (
    .a(_al_u2855_o),
    .b(\exu/shift_count [3]),
    .c(\exu/n50 [3]),
    .o(_al_u2864_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u2865 (
    .a(\exu/n49 ),
    .b(_al_u2864_o),
    .c(op_count[3]),
    .o(\exu/n52 [3]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u2866 (
    .a(_al_u2855_o),
    .b(\exu/shift_count [2]),
    .c(\exu/n50 [2]),
    .o(_al_u2866_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u2867 (
    .a(\exu/n49 ),
    .b(_al_u2866_o),
    .c(op_count[2]),
    .o(\exu/n52 [2]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u2868 (
    .a(_al_u2855_o),
    .b(\exu/shift_count [1]),
    .c(\exu/n50 [1]),
    .o(_al_u2868_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u2869 (
    .a(\exu/n49 ),
    .b(_al_u2868_o),
    .c(op_count[1]),
    .o(\exu/n52 [1]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u2870 (
    .a(_al_u2855_o),
    .b(\exu/shift_count [0]),
    .c(\exu/n50 [0]),
    .o(_al_u2870_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u2871 (
    .a(\exu/n49 ),
    .b(_al_u2870_o),
    .c(op_count[0]),
    .o(\exu/n52 [0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2872 (
    .a(_al_u2697_o),
    .b(rst_pad),
    .o(\biu/bus_unit/mmu/mux18_b3_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2873 (
    .a(\biu/bus_unit/addr_counter [6]),
    .b(\biu/bus_unit/addr_counter [7]),
    .c(\biu/bus_unit/addr_counter [8]),
    .o(_al_u2873_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2874 (
    .a(\biu/bus_unit/addr_counter [2]),
    .b(\biu/bus_unit/addr_counter [3]),
    .c(\biu/bus_unit/addr_counter [4]),
    .d(\biu/bus_unit/addr_counter [5]),
    .o(_al_u2874_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2875 (
    .a(_al_u2873_o),
    .b(_al_u2874_o),
    .c(\biu/bus_unit/addr_counter [0]),
    .d(\biu/bus_unit/addr_counter [1]),
    .o(\biu/bus_unit/n15_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2876 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(\biu/bus_unit/n39 [8]),
    .o(\biu/bus_unit/n39[8]_d ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2877 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(\biu/bus_unit/n39 [7]),
    .o(\biu/bus_unit/n39[7]_d ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2878 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(\biu/bus_unit/n39 [6]),
    .o(\biu/bus_unit/n39[6]_d ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2879 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(\biu/bus_unit/n39 [5]),
    .o(\biu/bus_unit/n39[5]_d ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2880 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(\biu/bus_unit/n39 [4]),
    .o(\biu/bus_unit/n39[4]_d ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2881 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(\biu/bus_unit/n39 [3]),
    .o(\biu/bus_unit/n39[3]_d ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2882 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(\biu/bus_unit/n39 [2]),
    .o(\biu/bus_unit/n39[2]_d ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2883 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(\biu/bus_unit/n39 [1]),
    .o(\biu/bus_unit/n39[1]_d ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2884 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(\biu/bus_unit/n39 [0]),
    .o(\biu/bus_unit/n39[0]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u2885 (
    .a(\biu/cache_ctrl_logic/statu [0]),
    .b(\biu/cache_ctrl_logic/statu [2]),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(_al_u2885_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2886 (
    .a(_al_u2885_o),
    .b(\biu/cache_ctrl_logic/statu [1]),
    .o(_al_u2886_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u2887 (
    .a(_al_u2837_o),
    .b(\biu/cache_ctrl_logic/statu [2]),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2888 (
    .a(_al_u2886_o),
    .b(\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ),
    .o(\biu/bus_unit/mux1_b1_sel_is_0_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2889 (
    .a(\biu/bus_unit/statu [0]),
    .b(\biu/bus_unit/statu [1]),
    .c(\biu/bus_unit/statu [3]),
    .o(_al_u2889_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2890 (
    .a(_al_u2703_o),
    .b(_al_u2889_o),
    .o(_al_u2890_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u2891 (
    .a(_al_u2890_o),
    .b(\biu/bus_unit/addr_counter [8]),
    .c(\biu/bus_unit/last_addr [8]),
    .o(_al_u2891_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2892 (
    .a(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .b(_al_u2891_o),
    .c(addr_ex[8]),
    .o(\biu/l1d_addr [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u2893 (
    .a(_al_u2890_o),
    .b(\biu/bus_unit/addr_counter [7]),
    .c(\biu/bus_unit/last_addr [7]),
    .o(_al_u2893_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2894 (
    .a(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .b(_al_u2893_o),
    .c(addr_ex[7]),
    .o(\biu/l1d_addr [7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u2895 (
    .a(_al_u2890_o),
    .b(\biu/bus_unit/addr_counter [6]),
    .c(\biu/bus_unit/last_addr [6]),
    .o(_al_u2895_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2896 (
    .a(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .b(_al_u2895_o),
    .c(addr_ex[6]),
    .o(\biu/l1d_addr [6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u2897 (
    .a(_al_u2890_o),
    .b(\biu/bus_unit/addr_counter [5]),
    .c(\biu/bus_unit/last_addr [5]),
    .o(_al_u2897_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2898 (
    .a(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .b(_al_u2897_o),
    .c(addr_ex[5]),
    .o(\biu/l1d_addr [5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u2899 (
    .a(_al_u2890_o),
    .b(\biu/bus_unit/addr_counter [4]),
    .c(\biu/bus_unit/last_addr [4]),
    .o(_al_u2899_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2900 (
    .a(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .b(_al_u2899_o),
    .c(addr_ex[4]),
    .o(\biu/l1d_addr [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u2901 (
    .a(_al_u2890_o),
    .b(\biu/bus_unit/addr_counter [3]),
    .c(\biu/bus_unit/last_addr [3]),
    .o(_al_u2901_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2902 (
    .a(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .b(_al_u2901_o),
    .c(addr_ex[3]),
    .o(\biu/l1d_addr [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u2903 (
    .a(_al_u2890_o),
    .b(\biu/bus_unit/addr_counter [2]),
    .c(\biu/bus_unit/last_addr [2]),
    .o(_al_u2903_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2904 (
    .a(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .b(_al_u2903_o),
    .c(addr_ex[2]),
    .o(\biu/l1d_addr [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u2905 (
    .a(_al_u2890_o),
    .b(\biu/bus_unit/addr_counter [1]),
    .c(\biu/bus_unit/last_addr [1]),
    .o(_al_u2905_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2906 (
    .a(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .b(_al_u2905_o),
    .c(addr_ex[1]),
    .o(\biu/l1d_addr [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u2907 (
    .a(_al_u2890_o),
    .b(\biu/bus_unit/addr_counter [0]),
    .c(\biu/bus_unit/last_addr [0]),
    .o(_al_u2907_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u2908 (
    .a(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .b(_al_u2907_o),
    .c(addr_ex[0]),
    .o(\biu/l1d_addr [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u2909 (
    .a(\exu/main_state [0]),
    .b(\exu/main_state [1]),
    .c(\exu/main_state [3]),
    .o(_al_u2909_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2910 (
    .a(_al_u2909_o),
    .b(\exu/main_state [2]),
    .o(_al_u2910_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*C)*~(B*A))"),
    .INIT(16'hf888))
    _al_u2911 (
    .a(load_acc_fault),
    .b(_al_u2910_o),
    .c(_al_u2838_o),
    .d(_al_u2847_o),
    .o(\exu/n90 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u2912 (
    .a(_al_u2847_o),
    .b(\biu/cache_ctrl_logic/statu [2]),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(\biu/cache_ctrl_logic/n75_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2913 (
    .a(_al_u2885_o),
    .b(\biu/cache_ctrl_logic/statu [1]),
    .o(\biu/bus_unit/mmu/n19_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2914 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .o(_al_u2914_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u2915 (
    .a(\biu/bus_unit/mmu/statu [0]),
    .b(\biu/bus_unit/mmu/statu [1]),
    .c(\biu/bus_unit/mmu/statu [2]),
    .d(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u2915_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u2916 (
    .a(_al_u2915_o),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .o(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2917 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [9]),
    .o(\biu/bus_unit/mmu/n66 [9]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2918 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [8]),
    .o(\biu/bus_unit/mmu/n66 [8]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2919 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [7]),
    .o(\biu/bus_unit/mmu/n66 [7]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2920 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [6]),
    .o(\biu/bus_unit/mmu/n66 [6]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2921 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [5]),
    .o(\biu/bus_unit/mmu/n66 [5]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2922 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [4]),
    .o(\biu/bus_unit/mmu/n66 [4]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2923 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [3]),
    .o(\biu/bus_unit/mmu/n66 [3]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2924 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [2]),
    .o(\biu/bus_unit/mmu/n66 [2]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2925 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [11]),
    .o(\biu/bus_unit/mmu/n66 [11]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2926 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [10]),
    .o(\biu/bus_unit/mmu/n66 [10]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2927 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [1]),
    .o(\biu/bus_unit/mmu/n66 [1]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h8b00))
    _al_u2928 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [0]),
    .o(\biu/bus_unit/mmu/n66 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2929 (
    .a(ins_read[4]),
    .b(ins_read[36]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2929_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2930 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [4]),
    .o(_al_u2930_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2931 (
    .a(ins_read[3]),
    .b(ins_read[35]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2931_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2932 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [3]),
    .o(_al_u2932_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(~B*~A))"),
    .INIT(16'heee0))
    _al_u2933 (
    .a(_al_u2929_o),
    .b(_al_u2930_o),
    .c(_al_u2931_o),
    .d(_al_u2932_o),
    .o(_al_u2933_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2934 (
    .a(ins_read[0]),
    .b(ins_read[32]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2934_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2935 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [0]),
    .o(_al_u2935_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2936 (
    .a(ins_read[1]),
    .b(ins_read[33]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2936_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2937 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [1]),
    .o(_al_u2937_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2938 (
    .a(_al_u2934_o),
    .b(_al_u2935_o),
    .c(_al_u2936_o),
    .d(_al_u2937_o),
    .o(_al_u2938_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u2939 (
    .a(\ins_fetch/ins_shift [2]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [2]),
    .o(_al_u2939_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2940 (
    .a(ins_read[6]),
    .b(ins_read[38]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2940_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2941 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [6]),
    .o(_al_u2941_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0305))
    _al_u2942 (
    .a(ins_read[5]),
    .b(ins_read[37]),
    .c(\ins_fetch/hold ),
    .d(id_ins_pc[2]),
    .o(_al_u2942_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2943 (
    .a(\ins_fetch/hold ),
    .b(\ins_fetch/ins_hold [5]),
    .o(_al_u2943_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*~A))"),
    .INIT(16'h000e))
    _al_u2944 (
    .a(_al_u2940_o),
    .b(_al_u2941_o),
    .c(_al_u2942_o),
    .d(_al_u2943_o),
    .o(_al_u2944_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u2945 (
    .a(_al_u2933_o),
    .b(_al_u2938_o),
    .c(_al_u2939_o),
    .d(_al_u2944_o),
    .o(\ins_dec/op_store ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(~B*~A))"),
    .INIT(16'heee0))
    _al_u2946 (
    .a(_al_u2940_o),
    .b(_al_u2941_o),
    .c(_al_u2942_o),
    .d(_al_u2943_o),
    .o(_al_u2946_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u2947 (
    .a(_al_u2933_o),
    .b(_al_u2938_o),
    .c(_al_u2939_o),
    .d(_al_u2946_o),
    .o(\ins_dec/op_load ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(~B*~A))"),
    .INIT(16'h000e))
    _al_u2948 (
    .a(_al_u2929_o),
    .b(_al_u2930_o),
    .c(_al_u2931_o),
    .d(_al_u2932_o),
    .o(_al_u2948_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2949 (
    .a(_al_u2938_o),
    .b(_al_u2939_o),
    .c(_al_u2944_o),
    .d(_al_u2948_o),
    .o(\ins_dec/op_amo ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2950 (
    .a(_al_u2938_o),
    .b(_al_u2939_o),
    .c(_al_u2946_o),
    .d(_al_u2948_o),
    .o(id_system));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u2951 (
    .a(_al_u2703_o),
    .b(\biu/bus_unit/statu [0]),
    .c(\biu/bus_unit/statu [1]),
    .d(\biu/bus_unit/statu [3]),
    .o(htrans_pad[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u2952 (
    .a(_al_u2703_o),
    .b(\biu/bus_unit/statu [0]),
    .c(\biu/bus_unit/statu [1]),
    .d(\biu/bus_unit/statu [3]),
    .o(_al_u2952_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(~C*~B)))"),
    .INIT(16'hfeaa))
    _al_u2953 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(htrans_pad[0]),
    .c(_al_u2952_o),
    .d(hready_pad),
    .o(\biu/bus_unit/n39[0]_en ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*B))"),
    .INIT(16'haaa2))
    _al_u2954 (
    .a(_al_u2705_o),
    .b(\biu/bus_unit/mmu/statu [0]),
    .c(\biu/bus_unit/mmu/statu [1]),
    .d(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u2954_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2955 (
    .a(\biu/bus_unit/statu [2]),
    .b(\biu/bus_unit/statu [3]),
    .c(\biu/bus_unit/statu [4]),
    .o(_al_u2955_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u2956 (
    .a(_al_u2955_o),
    .b(\biu/bus_unit/statu [0]),
    .c(\biu/bus_unit/statu [1]),
    .o(_al_u2956_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u2957 (
    .a(_al_u2706_o),
    .b(_al_u2956_o),
    .o(_al_u2957_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u2958 (
    .a(_al_u2703_o),
    .b(\biu/bus_unit/statu [0]),
    .c(\biu/bus_unit/statu [1]),
    .o(_al_u2958_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2959 (
    .a(_al_u2957_o),
    .b(_al_u2958_o),
    .o(\biu/bus_unit/mux15_b4_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u2960 (
    .a(_al_u2954_o),
    .b(\biu/bus_unit/mux15_b4_sel_is_2_o ),
    .c(htrans_pad[0]),
    .o(htrans_pad[1]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u2961 (
    .a(htrans_pad[0]),
    .b(_al_u2952_o),
    .o(hburst_pad[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u2962 (
    .a(satp[60]),
    .b(satp[61]),
    .c(satp[62]),
    .d(satp[63]),
    .o(\biu/bus_unit/mmu/n31_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u2963 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/n31_lutinv ),
    .o(_al_u2963_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u2964 (
    .a(\biu/bus_unit/mmu/statu [0]),
    .b(\biu/bus_unit/mmu/statu [1]),
    .c(\biu/bus_unit/mmu/statu [2]),
    .d(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u2964_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2965 (
    .a(_al_u2964_o),
    .b(hready_pad),
    .o(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u2966 (
    .a(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .b(hrdata_pad[9]),
    .c(\biu/bus_unit/mmu_hwdata [9]),
    .o(_al_u2966_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u2967 (
    .a(_al_u2963_o),
    .b(_al_u2966_o),
    .o(\biu/bus_unit/mmu/n79 [9]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2968 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [8]),
    .d(hrdata_pad[8]),
    .o(\biu/bus_unit/mmu/n79 [8]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2969 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [7]),
    .d(hrdata_pad[7]),
    .o(\biu/bus_unit/mmu/n79 [7]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2970 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [63]),
    .d(hrdata_pad[63]),
    .o(\biu/bus_unit/mmu/n79 [63]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2971 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [62]),
    .d(hrdata_pad[62]),
    .o(\biu/bus_unit/mmu/n79 [62]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2972 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [61]),
    .d(hrdata_pad[61]),
    .o(\biu/bus_unit/mmu/n79 [61]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2973 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [60]),
    .d(hrdata_pad[60]),
    .o(\biu/bus_unit/mmu/n79 [60]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u2974 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [6]),
    .o(_al_u2974_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u2975 (
    .a(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .b(_al_u2915_o),
    .c(hrdata_pad[6]),
    .o(_al_u2975_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u2976 (
    .a(_al_u2974_o),
    .b(_al_u2975_o),
    .o(\biu/bus_unit/mmu/n79 [6]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2977 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [59]),
    .d(hrdata_pad[59]),
    .o(\biu/bus_unit/mmu/n79 [59]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2978 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [58]),
    .d(hrdata_pad[58]),
    .o(\biu/bus_unit/mmu/n79 [58]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2979 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [57]),
    .d(hrdata_pad[57]),
    .o(\biu/bus_unit/mmu/n79 [57]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2980 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [56]),
    .d(hrdata_pad[56]),
    .o(\biu/bus_unit/mmu/n79 [56]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2981 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [55]),
    .d(hrdata_pad[55]),
    .o(\biu/bus_unit/mmu/n79 [55]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2982 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [54]),
    .d(hrdata_pad[54]),
    .o(\biu/bus_unit/mmu/n79 [54]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2983 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [53]),
    .d(hrdata_pad[53]),
    .o(\biu/bus_unit/mmu/n79 [53]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2984 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [52]),
    .d(hrdata_pad[52]),
    .o(\biu/bus_unit/mmu/n79 [52]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2985 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [51]),
    .d(hrdata_pad[51]),
    .o(\biu/bus_unit/mmu/n79 [51]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2986 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [50]),
    .d(hrdata_pad[50]),
    .o(\biu/bus_unit/mmu/n79 [50]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2987 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [5]),
    .d(hrdata_pad[5]),
    .o(\biu/bus_unit/mmu/n79 [5]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2988 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [49]),
    .d(hrdata_pad[49]),
    .o(\biu/bus_unit/mmu/n79 [49]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2989 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [48]),
    .d(hrdata_pad[48]),
    .o(\biu/bus_unit/mmu/n79 [48]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2990 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [47]),
    .d(hrdata_pad[47]),
    .o(\biu/bus_unit/mmu/n79 [47]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2991 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [46]),
    .d(hrdata_pad[46]),
    .o(\biu/bus_unit/mmu/n79 [46]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2992 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [45]),
    .d(hrdata_pad[45]),
    .o(\biu/bus_unit/mmu/n79 [45]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2993 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [44]),
    .d(hrdata_pad[44]),
    .o(\biu/bus_unit/mmu/n79 [44]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2994 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [43]),
    .d(hrdata_pad[43]),
    .o(\biu/bus_unit/mmu/n79 [43]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2995 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [42]),
    .d(hrdata_pad[42]),
    .o(\biu/bus_unit/mmu/n79 [42]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2996 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [41]),
    .d(hrdata_pad[41]),
    .o(\biu/bus_unit/mmu/n79 [41]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2997 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [40]),
    .d(hrdata_pad[40]),
    .o(\biu/bus_unit/mmu/n79 [40]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2998 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [4]),
    .d(hrdata_pad[4]),
    .o(\biu/bus_unit/mmu/n79 [4]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u2999 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [39]),
    .d(hrdata_pad[39]),
    .o(\biu/bus_unit/mmu/n79 [39]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3000 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [38]),
    .d(hrdata_pad[38]),
    .o(\biu/bus_unit/mmu/n79 [38]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3001 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [37]),
    .d(hrdata_pad[37]),
    .o(\biu/bus_unit/mmu/n79 [37]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3002 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [36]),
    .d(hrdata_pad[36]),
    .o(\biu/bus_unit/mmu/n79 [36]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3003 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [35]),
    .d(hrdata_pad[35]),
    .o(\biu/bus_unit/mmu/n79 [35]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3004 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [34]),
    .d(hrdata_pad[34]),
    .o(\biu/bus_unit/mmu/n79 [34]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3005 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [33]),
    .d(hrdata_pad[33]),
    .o(\biu/bus_unit/mmu/n79 [33]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3006 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [32]),
    .d(hrdata_pad[32]),
    .o(\biu/bus_unit/mmu/n79 [32]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3007 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [31]),
    .d(hrdata_pad[31]),
    .o(\biu/bus_unit/mmu/n79 [31]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3008 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [30]),
    .d(hrdata_pad[30]),
    .o(\biu/bus_unit/mmu/n79 [30]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3009 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [3]),
    .d(hrdata_pad[3]),
    .o(\biu/bus_unit/mmu/n79 [3]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3010 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [29]),
    .d(hrdata_pad[29]),
    .o(\biu/bus_unit/mmu/n79 [29]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3011 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [28]),
    .d(hrdata_pad[28]),
    .o(\biu/bus_unit/mmu/n79 [28]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3012 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [27]),
    .d(hrdata_pad[27]),
    .o(\biu/bus_unit/mmu/n79 [27]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3013 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [26]),
    .d(hrdata_pad[26]),
    .o(\biu/bus_unit/mmu/n79 [26]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3014 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [25]),
    .d(hrdata_pad[25]),
    .o(\biu/bus_unit/mmu/n79 [25]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3015 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [24]),
    .d(hrdata_pad[24]),
    .o(\biu/bus_unit/mmu/n79 [24]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3016 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [23]),
    .d(hrdata_pad[23]),
    .o(\biu/bus_unit/mmu/n79 [23]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3017 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [22]),
    .d(hrdata_pad[22]),
    .o(\biu/bus_unit/mmu/n79 [22]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3018 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [21]),
    .d(hrdata_pad[21]),
    .o(\biu/bus_unit/mmu/n79 [21]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3019 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [20]),
    .d(hrdata_pad[20]),
    .o(\biu/bus_unit/mmu/n79 [20]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3020 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [2]),
    .d(hrdata_pad[2]),
    .o(\biu/bus_unit/mmu/n79 [2]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3021 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [19]),
    .d(hrdata_pad[19]),
    .o(\biu/bus_unit/mmu/n79 [19]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3022 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [18]),
    .d(hrdata_pad[18]),
    .o(\biu/bus_unit/mmu/n79 [18]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3023 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [17]),
    .d(hrdata_pad[17]),
    .o(\biu/bus_unit/mmu/n79 [17]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3024 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [16]),
    .d(hrdata_pad[16]),
    .o(\biu/bus_unit/mmu/n79 [16]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3025 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [15]),
    .d(hrdata_pad[15]),
    .o(\biu/bus_unit/mmu/n79 [15]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3026 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [14]),
    .d(hrdata_pad[14]),
    .o(\biu/bus_unit/mmu/n79 [14]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3027 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [13]),
    .d(hrdata_pad[13]),
    .o(\biu/bus_unit/mmu/n79 [13]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3028 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [12]),
    .d(hrdata_pad[12]),
    .o(\biu/bus_unit/mmu/n79 [12]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3029 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [11]),
    .d(hrdata_pad[11]),
    .o(\biu/bus_unit/mmu/n79 [11]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3030 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [10]),
    .d(hrdata_pad[10]),
    .o(\biu/bus_unit/mmu/n79 [10]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3031 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [1]),
    .d(hrdata_pad[1]),
    .o(\biu/bus_unit/mmu/n79 [1]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'hfeba))
    _al_u3032 (
    .a(_al_u2963_o),
    .b(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .c(\biu/bus_unit/mmu_hwdata [0]),
    .d(hrdata_pad[0]),
    .o(\biu/bus_unit/mmu/n79 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3033 (
    .a(_al_u2914_o),
    .b(\biu/bus_unit/mmu/n31_lutinv ),
    .o(_al_u3033_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u3034 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(_al_u3034_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3035 (
    .a(_al_u3034_o),
    .b(\biu/paddress [127]),
    .o(\biu/bus_unit/mmu/n71 [63]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3036 (
    .a(_al_u3034_o),
    .b(\biu/paddress [126]),
    .o(\biu/bus_unit/mmu/n71 [62]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3037 (
    .a(_al_u3034_o),
    .b(\biu/paddress [125]),
    .o(\biu/bus_unit/mmu/n71 [61]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3038 (
    .a(_al_u3034_o),
    .b(\biu/paddress [124]),
    .o(\biu/bus_unit/mmu/n71 [60]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3039 (
    .a(_al_u3034_o),
    .b(\biu/paddress [123]),
    .o(\biu/bus_unit/mmu/n71 [59]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3040 (
    .a(_al_u3034_o),
    .b(\biu/paddress [122]),
    .o(\biu/bus_unit/mmu/n71 [58]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3041 (
    .a(_al_u3034_o),
    .b(\biu/paddress [121]),
    .o(\biu/bus_unit/mmu/n71 [57]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3042 (
    .a(_al_u3034_o),
    .b(\biu/paddress [120]),
    .o(\biu/bus_unit/mmu/n71 [56]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3043 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [119]),
    .d(satp[43]),
    .o(_al_u3043_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3044 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [119]),
    .d(\biu/bus_unit/mmu_hwdata [53]),
    .o(_al_u3044_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3045 (
    .a(_al_u3043_o),
    .b(_al_u3044_o),
    .o(\biu/bus_unit/mmu/n71 [55]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3046 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [118]),
    .d(satp[42]),
    .o(_al_u3046_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3047 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [118]),
    .d(\biu/bus_unit/mmu_hwdata [52]),
    .o(_al_u3047_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3048 (
    .a(_al_u3046_o),
    .b(_al_u3047_o),
    .o(\biu/bus_unit/mmu/n71 [54]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3049 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [117]),
    .d(satp[41]),
    .o(_al_u3049_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3050 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [117]),
    .d(\biu/bus_unit/mmu_hwdata [51]),
    .o(_al_u3050_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3051 (
    .a(_al_u3049_o),
    .b(_al_u3050_o),
    .o(\biu/bus_unit/mmu/n71 [53]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3052 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [116]),
    .d(satp[40]),
    .o(_al_u3052_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3053 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [116]),
    .d(\biu/bus_unit/mmu_hwdata [50]),
    .o(_al_u3053_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3054 (
    .a(_al_u3052_o),
    .b(_al_u3053_o),
    .o(\biu/bus_unit/mmu/n71 [52]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3055 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [115]),
    .d(satp[39]),
    .o(_al_u3055_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3056 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [115]),
    .d(\biu/bus_unit/mmu_hwdata [49]),
    .o(_al_u3056_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3057 (
    .a(_al_u3055_o),
    .b(_al_u3056_o),
    .o(\biu/bus_unit/mmu/n71 [51]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3058 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [114]),
    .d(satp[38]),
    .o(_al_u3058_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3059 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [114]),
    .d(\biu/bus_unit/mmu_hwdata [48]),
    .o(_al_u3059_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3060 (
    .a(_al_u3058_o),
    .b(_al_u3059_o),
    .o(\biu/bus_unit/mmu/n71 [50]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3061 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [113]),
    .d(satp[37]),
    .o(_al_u3061_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3062 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [113]),
    .d(\biu/bus_unit/mmu_hwdata [47]),
    .o(_al_u3062_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3063 (
    .a(_al_u3061_o),
    .b(_al_u3062_o),
    .o(\biu/bus_unit/mmu/n71 [49]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3064 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [112]),
    .d(satp[36]),
    .o(_al_u3064_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3065 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [112]),
    .d(\biu/bus_unit/mmu_hwdata [46]),
    .o(_al_u3065_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3066 (
    .a(_al_u3064_o),
    .b(_al_u3065_o),
    .o(\biu/bus_unit/mmu/n71 [48]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3067 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [111]),
    .d(satp[35]),
    .o(_al_u3067_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3068 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [111]),
    .d(\biu/bus_unit/mmu_hwdata [45]),
    .o(_al_u3068_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3069 (
    .a(_al_u3067_o),
    .b(_al_u3068_o),
    .o(\biu/bus_unit/mmu/n71 [47]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3070 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [110]),
    .d(satp[34]),
    .o(_al_u3070_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3071 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [110]),
    .d(\biu/bus_unit/mmu_hwdata [44]),
    .o(_al_u3071_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3072 (
    .a(_al_u3070_o),
    .b(_al_u3071_o),
    .o(\biu/bus_unit/mmu/n71 [46]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3073 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [109]),
    .d(satp[33]),
    .o(_al_u3073_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3074 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [109]),
    .d(\biu/bus_unit/mmu_hwdata [43]),
    .o(_al_u3074_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3075 (
    .a(_al_u3073_o),
    .b(_al_u3074_o),
    .o(\biu/bus_unit/mmu/n71 [45]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3076 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [108]),
    .d(satp[32]),
    .o(_al_u3076_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3077 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [108]),
    .d(\biu/bus_unit/mmu_hwdata [42]),
    .o(_al_u3077_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3078 (
    .a(_al_u3076_o),
    .b(_al_u3077_o),
    .o(\biu/bus_unit/mmu/n71 [44]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3079 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [107]),
    .d(satp[31]),
    .o(_al_u3079_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3080 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [107]),
    .d(\biu/bus_unit/mmu_hwdata [41]),
    .o(_al_u3080_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3081 (
    .a(_al_u3079_o),
    .b(_al_u3080_o),
    .o(\biu/bus_unit/mmu/n71 [43]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3082 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [106]),
    .d(satp[30]),
    .o(_al_u3082_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3083 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [106]),
    .d(\biu/bus_unit/mmu_hwdata [40]),
    .o(_al_u3083_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3084 (
    .a(_al_u3082_o),
    .b(_al_u3083_o),
    .o(\biu/bus_unit/mmu/n71 [42]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3085 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [105]),
    .d(satp[29]),
    .o(_al_u3085_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3086 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [105]),
    .d(\biu/bus_unit/mmu_hwdata [39]),
    .o(_al_u3086_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3087 (
    .a(_al_u3085_o),
    .b(_al_u3086_o),
    .o(\biu/bus_unit/mmu/n71 [41]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3088 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [104]),
    .d(satp[28]),
    .o(_al_u3088_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3089 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [104]),
    .d(\biu/bus_unit/mmu_hwdata [38]),
    .o(_al_u3089_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3090 (
    .a(_al_u3088_o),
    .b(_al_u3089_o),
    .o(\biu/bus_unit/mmu/n71 [40]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3091 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [103]),
    .d(satp[27]),
    .o(_al_u3091_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3092 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [103]),
    .d(\biu/bus_unit/mmu_hwdata [37]),
    .o(_al_u3092_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3093 (
    .a(_al_u3091_o),
    .b(_al_u3092_o),
    .o(\biu/bus_unit/mmu/n71 [39]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3094 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [102]),
    .d(satp[26]),
    .o(_al_u3094_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3095 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [102]),
    .d(\biu/bus_unit/mmu_hwdata [36]),
    .o(_al_u3095_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3096 (
    .a(_al_u3094_o),
    .b(_al_u3095_o),
    .o(\biu/bus_unit/mmu/n71 [38]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3097 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [101]),
    .d(satp[25]),
    .o(_al_u3097_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3098 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [101]),
    .d(\biu/bus_unit/mmu_hwdata [35]),
    .o(_al_u3098_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3099 (
    .a(_al_u3097_o),
    .b(_al_u3098_o),
    .o(\biu/bus_unit/mmu/n71 [37]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3100 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [100]),
    .d(satp[24]),
    .o(_al_u3100_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3101 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [100]),
    .d(\biu/bus_unit/mmu_hwdata [34]),
    .o(_al_u3101_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3102 (
    .a(_al_u3100_o),
    .b(_al_u3101_o),
    .o(\biu/bus_unit/mmu/n71 [36]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3103 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [99]),
    .d(satp[23]),
    .o(_al_u3103_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3104 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [99]),
    .d(\biu/bus_unit/mmu_hwdata [33]),
    .o(_al_u3104_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3105 (
    .a(_al_u3103_o),
    .b(_al_u3104_o),
    .o(\biu/bus_unit/mmu/n71 [35]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3106 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [98]),
    .d(satp[22]),
    .o(_al_u3106_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3107 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [98]),
    .d(\biu/bus_unit/mmu_hwdata [32]),
    .o(_al_u3107_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3108 (
    .a(_al_u3106_o),
    .b(_al_u3107_o),
    .o(\biu/bus_unit/mmu/n71 [34]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3109 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [97]),
    .d(satp[21]),
    .o(_al_u3109_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3110 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [97]),
    .d(\biu/bus_unit/mmu_hwdata [31]),
    .o(_al_u3110_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3111 (
    .a(_al_u3109_o),
    .b(_al_u3110_o),
    .o(\biu/bus_unit/mmu/n71 [33]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3112 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [96]),
    .d(satp[20]),
    .o(_al_u3112_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3113 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [96]),
    .d(\biu/bus_unit/mmu_hwdata [30]),
    .o(_al_u3113_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3114 (
    .a(_al_u3112_o),
    .b(_al_u3113_o),
    .o(\biu/bus_unit/mmu/n71 [32]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3115 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [95]),
    .d(satp[19]),
    .o(_al_u3115_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3116 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [95]),
    .d(\biu/bus_unit/mmu_hwdata [29]),
    .o(_al_u3116_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3117 (
    .a(_al_u3115_o),
    .b(_al_u3116_o),
    .o(\biu/bus_unit/mmu/n71 [31]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3118 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [94]),
    .d(satp[18]),
    .o(_al_u3118_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3119 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [94]),
    .d(\biu/bus_unit/mmu_hwdata [28]),
    .o(_al_u3119_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3120 (
    .a(_al_u3118_o),
    .b(_al_u3119_o),
    .o(\biu/bus_unit/mmu/n71 [30]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3121 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [93]),
    .d(satp[17]),
    .o(_al_u3121_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3122 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [93]),
    .d(\biu/bus_unit/mmu_hwdata [27]),
    .o(_al_u3122_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3123 (
    .a(_al_u3121_o),
    .b(_al_u3122_o),
    .o(\biu/bus_unit/mmu/n71 [29]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3124 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [92]),
    .d(satp[16]),
    .o(_al_u3124_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3125 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [92]),
    .d(\biu/bus_unit/mmu_hwdata [26]),
    .o(_al_u3125_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3126 (
    .a(_al_u3124_o),
    .b(_al_u3125_o),
    .o(\biu/bus_unit/mmu/n71 [28]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3127 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [91]),
    .d(satp[15]),
    .o(_al_u3127_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3128 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [91]),
    .d(\biu/bus_unit/mmu_hwdata [25]),
    .o(_al_u3128_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3129 (
    .a(_al_u3127_o),
    .b(_al_u3128_o),
    .o(\biu/bus_unit/mmu/n71 [27]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3130 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [90]),
    .d(satp[14]),
    .o(_al_u3130_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3131 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [90]),
    .d(\biu/bus_unit/mmu_hwdata [24]),
    .o(_al_u3131_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3132 (
    .a(_al_u3130_o),
    .b(_al_u3131_o),
    .o(\biu/bus_unit/mmu/n71 [26]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3133 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [89]),
    .d(satp[13]),
    .o(_al_u3133_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3134 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [89]),
    .d(\biu/bus_unit/mmu_hwdata [23]),
    .o(_al_u3134_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3135 (
    .a(_al_u3133_o),
    .b(_al_u3134_o),
    .o(\biu/bus_unit/mmu/n71 [25]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3136 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [88]),
    .d(satp[12]),
    .o(_al_u3136_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3137 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [88]),
    .d(\biu/bus_unit/mmu_hwdata [22]),
    .o(_al_u3137_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3138 (
    .a(_al_u3136_o),
    .b(_al_u3137_o),
    .o(\biu/bus_unit/mmu/n71 [24]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3139 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [87]),
    .d(satp[11]),
    .o(_al_u3139_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3140 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [87]),
    .d(\biu/bus_unit/mmu_hwdata [21]),
    .o(_al_u3140_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3141 (
    .a(_al_u3139_o),
    .b(_al_u3140_o),
    .o(\biu/bus_unit/mmu/n71 [23]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3142 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [86]),
    .d(satp[10]),
    .o(_al_u3142_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3143 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [86]),
    .d(\biu/bus_unit/mmu_hwdata [20]),
    .o(_al_u3143_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3144 (
    .a(_al_u3142_o),
    .b(_al_u3143_o),
    .o(\biu/bus_unit/mmu/n71 [22]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3145 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [85]),
    .d(satp[9]),
    .o(_al_u3145_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3146 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [85]),
    .d(\biu/bus_unit/mmu_hwdata [19]),
    .o(_al_u3146_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3147 (
    .a(_al_u3145_o),
    .b(_al_u3146_o),
    .o(\biu/bus_unit/mmu/n71 [21]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3148 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [84]),
    .d(satp[8]),
    .o(_al_u3148_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3149 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [84]),
    .d(\biu/bus_unit/mmu_hwdata [18]),
    .o(_al_u3149_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3150 (
    .a(_al_u3148_o),
    .b(_al_u3149_o),
    .o(\biu/bus_unit/mmu/n71 [20]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3151 (
    .a(_al_u3034_o),
    .b(\biu/paddress [66]),
    .o(\biu/bus_unit/mmu/n71 [2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3152 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [83]),
    .d(satp[7]),
    .o(_al_u3152_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3153 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [83]),
    .d(\biu/bus_unit/mmu_hwdata [17]),
    .o(_al_u3153_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3154 (
    .a(_al_u3152_o),
    .b(_al_u3153_o),
    .o(\biu/bus_unit/mmu/n71 [19]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3155 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [82]),
    .d(satp[6]),
    .o(_al_u3155_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3156 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [82]),
    .d(\biu/bus_unit/mmu_hwdata [16]),
    .o(_al_u3156_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3157 (
    .a(_al_u3155_o),
    .b(_al_u3156_o),
    .o(\biu/bus_unit/mmu/n71 [18]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3158 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [81]),
    .d(satp[5]),
    .o(_al_u3158_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3159 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [81]),
    .d(\biu/bus_unit/mmu_hwdata [15]),
    .o(_al_u3159_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3160 (
    .a(_al_u3158_o),
    .b(_al_u3159_o),
    .o(\biu/bus_unit/mmu/n71 [17]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3161 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [80]),
    .d(satp[4]),
    .o(_al_u3161_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3162 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [80]),
    .d(\biu/bus_unit/mmu_hwdata [14]),
    .o(_al_u3162_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3163 (
    .a(_al_u3161_o),
    .b(_al_u3162_o),
    .o(\biu/bus_unit/mmu/n71 [16]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3164 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [79]),
    .d(satp[3]),
    .o(_al_u3164_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3165 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [79]),
    .d(\biu/bus_unit/mmu_hwdata [13]),
    .o(_al_u3165_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3166 (
    .a(_al_u3164_o),
    .b(_al_u3165_o),
    .o(\biu/bus_unit/mmu/n71 [15]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3167 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [78]),
    .d(satp[2]),
    .o(_al_u3167_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3168 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [78]),
    .d(\biu/bus_unit/mmu_hwdata [12]),
    .o(_al_u3168_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3169 (
    .a(_al_u3167_o),
    .b(_al_u3168_o),
    .o(\biu/bus_unit/mmu/n71 [14]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3170 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [77]),
    .d(satp[1]),
    .o(_al_u3170_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3171 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [77]),
    .d(\biu/bus_unit/mmu_hwdata [11]),
    .o(_al_u3171_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3172 (
    .a(_al_u3170_o),
    .b(_al_u3171_o),
    .o(\biu/bus_unit/mmu/n71 [13]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u3173 (
    .a(_al_u3033_o),
    .b(_al_u2698_o),
    .c(\biu/paddress [76]),
    .d(satp[0]),
    .o(_al_u3173_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u3174 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .c(\biu/paddress [76]),
    .d(\biu/bus_unit/mmu_hwdata [10]),
    .o(_al_u3174_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3175 (
    .a(_al_u3173_o),
    .b(_al_u3174_o),
    .o(\biu/bus_unit/mmu/n71 [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3176 (
    .a(_al_u3034_o),
    .b(\biu/paddress [65]),
    .o(\biu/bus_unit/mmu/n71 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3177 (
    .a(_al_u3034_o),
    .b(\biu/paddress [64]),
    .o(\biu/bus_unit/mmu/n71 [0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3178 (
    .a(addr_ex[0]),
    .b(addr_ex[1]),
    .o(\exu/lsu/n0_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdd50))
    _al_u3179 (
    .a(\exu/lsu/n0_lutinv ),
    .b(addr_ex[2]),
    .c(ex_size[2]),
    .d(ex_size[3]),
    .o(_al_u3179_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3180 (
    .a(addr_ex[0]),
    .b(addr_ex[1]),
    .o(\exu/lsu/n8_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u3181 (
    .a(_al_u3179_o),
    .b(\exu/lsu/n8_lutinv ),
    .c(addr_ex[2]),
    .d(ex_size[1]),
    .o(_al_u3181_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u3182 (
    .a(_al_u3181_o),
    .b(amo),
    .c(load),
    .o(\exu/load_addr_mis ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3183 (
    .a(csr_index[0]),
    .b(csr_index[3]),
    .c(csr_index[4]),
    .d(csr_index[5]),
    .o(_al_u3183_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3184 (
    .a(wb_csr_write),
    .b(wb_valid),
    .o(_al_u3184_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3185 (
    .a(_al_u3183_o),
    .b(_al_u3184_o),
    .c(csr_index[1]),
    .d(csr_index[2]),
    .o(_al_u3185_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3186 (
    .a(csr_index[10]),
    .b(csr_index[11]),
    .c(csr_index[9]),
    .o(_al_u3186_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3187 (
    .a(_al_u3186_o),
    .b(csr_index[6]),
    .c(csr_index[7]),
    .d(csr_index[8]),
    .o(_al_u3187_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3188 (
    .a(_al_u3185_o),
    .b(_al_u3187_o),
    .o(\cu_ru/csr_satp/n0 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3189 (
    .a(csr_index[10]),
    .b(csr_index[11]),
    .c(csr_index[9]),
    .o(_al_u3189_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3190 (
    .a(_al_u3189_o),
    .b(csr_index[6]),
    .c(csr_index[7]),
    .d(csr_index[8]),
    .o(_al_u3190_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3191 (
    .a(_al_u3183_o),
    .b(_al_u3184_o),
    .c(csr_index[1]),
    .d(csr_index[2]),
    .o(_al_u3191_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3192 (
    .a(_al_u3190_o),
    .b(_al_u3191_o),
    .o(\cu_ru/m_s_ip/n0 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3193 (
    .a(_al_u3185_o),
    .b(_al_u3190_o),
    .o(\cu_ru/m_s_scratch/n0 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3194 (
    .a(csr_index[6]),
    .b(csr_index[7]),
    .c(csr_index[8]),
    .o(_al_u3194_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3195 (
    .a(_al_u3189_o),
    .b(_al_u3194_o),
    .o(_al_u3195_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3196 (
    .a(_al_u3185_o),
    .b(_al_u3195_o),
    .o(\cu_ru/m_s_status/n0 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u3197 (
    .a(csr_index[0]),
    .b(csr_index[1]),
    .c(csr_index[2]),
    .d(csr_index[5]),
    .o(_al_u3197_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3198 (
    .a(_al_u3197_o),
    .b(csr_index[3]),
    .c(csr_index[4]),
    .o(_al_u3198_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3199 (
    .a(_al_u3195_o),
    .b(_al_u3198_o),
    .c(_al_u3184_o),
    .o(\cu_ru/m_cycle_event/n13 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u3200 (
    .a(csr_index[0]),
    .b(csr_index[3]),
    .c(csr_index[4]),
    .d(csr_index[5]),
    .o(_al_u3200_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3201 (
    .a(_al_u3184_o),
    .b(_al_u3200_o),
    .c(csr_index[1]),
    .d(csr_index[2]),
    .o(_al_u3201_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3202 (
    .a(_al_u3195_o),
    .b(_al_u3201_o),
    .o(\cu_ru/m_s_tvec/n0 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3203 (
    .a(_al_u3191_o),
    .b(_al_u3195_o),
    .o(\cu_ru/m_s_ie/n0 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3204 (
    .a(_al_u3200_o),
    .b(csr_index[1]),
    .c(csr_index[2]),
    .o(_al_u3204_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3205 (
    .a(_al_u3195_o),
    .b(_al_u3204_o),
    .c(_al_u3184_o),
    .o(\cu_ru/mideleg_int_ctrl/n0 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3206 (
    .a(_al_u3183_o),
    .b(csr_index[1]),
    .c(csr_index[2]),
    .o(_al_u3206_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3207 (
    .a(_al_u3195_o),
    .b(_al_u3206_o),
    .c(_al_u3184_o),
    .o(\cu_ru/medeleg_exc_ctrl/n0 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3208 (
    .a(_al_u2909_o),
    .b(\exu/main_state [2]),
    .o(\exu/c_fence_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3209 (
    .a(\biu/cache_ctrl_logic/statu [0]),
    .b(\biu/cache_ctrl_logic/statu [1]),
    .o(_al_u3209_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u3210 (
    .a(_al_u3209_o),
    .b(\biu/cache_ctrl_logic/statu [2]),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(\biu/cache_ctrl_logic/n55_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*B*A))"),
    .INIT(16'h070f))
    _al_u3211 (
    .a(\exu/c_fence_lutinv ),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(rst_pad),
    .d(cache_flush),
    .o(\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3212 (
    .a(_al_u2940_o),
    .b(_al_u2941_o),
    .c(_al_u2942_o),
    .d(_al_u2943_o),
    .o(_al_u3212_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3213 (
    .a(_al_u2933_o),
    .b(_al_u2938_o),
    .c(_al_u2939_o),
    .d(_al_u3212_o),
    .o(_al_u3213_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3214 (
    .a(_al_u2938_o),
    .b(_al_u2939_o),
    .c(_al_u2948_o),
    .d(_al_u3212_o),
    .o(_al_u3214_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u3215 (
    .a(_al_u3213_o),
    .b(_al_u3214_o),
    .o(\ins_dec/n59 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u3216 (
    .a(\ins_fetch/ins_shift [14]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [14]),
    .o(_al_u3216_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u3217 (
    .a(\ins_fetch/ins_shift [13]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [13]),
    .o(_al_u3217_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3218 (
    .a(_al_u3216_o),
    .b(_al_u3217_o),
    .o(\ins_dec/n35_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3219 (
    .a(id_system),
    .b(\ins_dec/n35_lutinv ),
    .o(\ins_dec/ins_fence ));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(~B*~(D*~C)))"),
    .INIT(16'h7577))
    _al_u3220 (
    .a(_al_u2706_o),
    .b(ex_size[0]),
    .c(ex_size[1]),
    .d(ex_size[2]),
    .o(hsize_pad[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3221 (
    .a(_al_u2838_o),
    .b(_al_u3209_o),
    .o(\biu/cache_ctrl_logic/n97_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u3222 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u2847_o),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(_al_u3222_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u3223 (
    .a(\biu/cache_ctrl_logic/statu [1]),
    .b(\biu/cache_ctrl_logic/statu [2]),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(\biu/cache_ctrl_logic/n204_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3224 (
    .a(\biu/cache_ctrl_logic/n204_lutinv ),
    .b(\biu/cache_ctrl_logic/statu [0]),
    .o(_al_u3224_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3225 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[9]),
    .o(\biu/cache_ctrl_logic/off [9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3226 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[8]),
    .o(\biu/cache_ctrl_logic/off [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3227 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[7]),
    .o(\biu/cache_ctrl_logic/off [7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3228 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[6]),
    .o(\biu/cache_ctrl_logic/off [6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3229 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[5]),
    .o(\biu/cache_ctrl_logic/off [5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3230 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[4]),
    .o(\biu/cache_ctrl_logic/off [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3231 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[3]),
    .o(\biu/cache_ctrl_logic/off [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3232 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[2]),
    .o(\biu/cache_ctrl_logic/off [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3233 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[11]),
    .o(\biu/cache_ctrl_logic/off [11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3234 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[10]),
    .o(\biu/cache_ctrl_logic/off [10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3235 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[1]),
    .o(\biu/cache_ctrl_logic/off [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u3236 (
    .a(_al_u3222_o),
    .b(_al_u3224_o),
    .c(addr_ex[0]),
    .o(\biu/cache_ctrl_logic/off [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3237 (
    .a(\cu_ru/m_sie [7]),
    .b(\cu_ru/m_sip [7]),
    .c(\cu_ru/mie ),
    .o(_al_u3237_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3238 (
    .a(\cu_ru/m_sie [3]),
    .b(\cu_ru/m_sip [3]),
    .c(\cu_ru/mie ),
    .o(_al_u3238_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3239 (
    .a(_al_u3237_o),
    .b(_al_u3238_o),
    .o(\cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*B))"),
    .INIT(16'haa2a))
    _al_u3240 (
    .a(\cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ),
    .b(\cu_ru/m_sip [5]),
    .c(\cu_ru/mie ),
    .d(\cu_ru/mideleg [5]),
    .o(_al_u3240_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(~B*~A))"),
    .INIT(16'h00e0))
    _al_u3241 (
    .a(s_ext_int_pad),
    .b(\cu_ru/m_s_ip/seip ),
    .c(\cu_ru/mie ),
    .d(\cu_ru/mideleg [9]),
    .o(\cu_ru/mideleg_int_ctrl/sei_ack_m ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u3242 (
    .a(\cu_ru/mideleg_int_ctrl/sei_ack_m ),
    .b(\cu_ru/m_sip [1]),
    .c(\cu_ru/mie ),
    .d(\cu_ru/mideleg [1]),
    .o(_al_u3242_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3243 (
    .a(_al_u3240_o),
    .b(_al_u3242_o),
    .o(\cu_ru/mideleg_int_ctrl/n28_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*B*~(~C*~A))"),
    .INIT(16'hc800))
    _al_u3244 (
    .a(s_ext_int_pad),
    .b(\cu_ru/m_sie [9]),
    .c(\cu_ru/m_s_ip/seip ),
    .d(\cu_ru/mideleg [9]),
    .o(_al_u3244_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u3245 (
    .a(_al_u3244_o),
    .b(\cu_ru/m_sie [1]),
    .c(\cu_ru/m_sip [1]),
    .d(\cu_ru/mideleg [1]),
    .o(_al_u3245_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3246 (
    .a(priv[0]),
    .b(priv[1]),
    .o(\cu_ru/m_s_status/n5 [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3247 (
    .a(_al_u3245_o),
    .b(\cu_ru/m_s_status/n5 [1]),
    .c(\cu_ru/mstatus [1]),
    .o(\cu_ru/mideleg_int_ctrl/n29_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3248 (
    .a(\cu_ru/m_sie [5]),
    .b(\cu_ru/m_sip [5]),
    .c(\cu_ru/mideleg [5]),
    .o(_al_u3248_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u3249 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(_al_u3248_o),
    .c(\cu_ru/mstatus [1]),
    .o(\cu_ru/mideleg_int_ctrl/sti_ack_s ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3250 (
    .a(\cu_ru/mideleg_int_ctrl/n29_lutinv ),
    .b(\cu_ru/mideleg_int_ctrl/sti_ack_s ),
    .o(_al_u3250_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u3251 (
    .a(\cu_ru/mideleg_int_ctrl/n28_lutinv ),
    .b(_al_u3250_o),
    .o(int_req));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3252 (
    .a(_al_u3194_o),
    .b(csr_index[10]),
    .c(csr_index[11]),
    .d(csr_index[9]),
    .o(_al_u3252_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3253 (
    .a(_al_u3185_o),
    .b(_al_u3252_o),
    .o(_al_u3253_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3254 (
    .a(\cu_ru/m_cycle_event/n2 [9]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [9]),
    .o(_al_u3254_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3255 (
    .a(_al_u3253_o),
    .b(_al_u3254_o),
    .c(data_csr[9]),
    .o(\cu_ru/m_cycle_event/n9 [9]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3256 (
    .a(\cu_ru/m_cycle_event/n2 [8]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [8]),
    .o(_al_u3256_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3257 (
    .a(_al_u3253_o),
    .b(_al_u3256_o),
    .c(data_csr[8]),
    .o(\cu_ru/m_cycle_event/n9 [8]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3258 (
    .a(\cu_ru/m_cycle_event/n2 [7]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [7]),
    .o(_al_u3258_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3259 (
    .a(_al_u3253_o),
    .b(_al_u3258_o),
    .c(data_csr[7]),
    .o(\cu_ru/m_cycle_event/n9 [7]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3260 (
    .a(\cu_ru/m_cycle_event/n2 [63]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [63]),
    .o(_al_u3260_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3261 (
    .a(_al_u3253_o),
    .b(_al_u3260_o),
    .c(data_csr[63]),
    .o(\cu_ru/m_cycle_event/n9 [63]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3262 (
    .a(\cu_ru/m_cycle_event/n2 [62]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [62]),
    .o(_al_u3262_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3263 (
    .a(_al_u3253_o),
    .b(_al_u3262_o),
    .c(data_csr[62]),
    .o(\cu_ru/m_cycle_event/n9 [62]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3264 (
    .a(\cu_ru/m_cycle_event/n2 [61]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [61]),
    .o(_al_u3264_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3265 (
    .a(_al_u3253_o),
    .b(_al_u3264_o),
    .c(data_csr[61]),
    .o(\cu_ru/m_cycle_event/n9 [61]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3266 (
    .a(\cu_ru/m_cycle_event/n2 [60]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [60]),
    .o(_al_u3266_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3267 (
    .a(_al_u3253_o),
    .b(_al_u3266_o),
    .c(data_csr[60]),
    .o(\cu_ru/m_cycle_event/n9 [60]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3268 (
    .a(\cu_ru/m_cycle_event/n2 [6]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [6]),
    .o(_al_u3268_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3269 (
    .a(_al_u3253_o),
    .b(_al_u3268_o),
    .c(data_csr[6]),
    .o(\cu_ru/m_cycle_event/n9 [6]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3270 (
    .a(\cu_ru/m_cycle_event/n2 [59]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [59]),
    .o(_al_u3270_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3271 (
    .a(_al_u3253_o),
    .b(_al_u3270_o),
    .c(data_csr[59]),
    .o(\cu_ru/m_cycle_event/n9 [59]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3272 (
    .a(\cu_ru/m_cycle_event/n2 [58]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [58]),
    .o(_al_u3272_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3273 (
    .a(_al_u3253_o),
    .b(_al_u3272_o),
    .c(data_csr[58]),
    .o(\cu_ru/m_cycle_event/n9 [58]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3274 (
    .a(\cu_ru/m_cycle_event/n2 [57]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [57]),
    .o(_al_u3274_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3275 (
    .a(_al_u3253_o),
    .b(_al_u3274_o),
    .c(data_csr[57]),
    .o(\cu_ru/m_cycle_event/n9 [57]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3276 (
    .a(\cu_ru/m_cycle_event/n2 [56]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [56]),
    .o(_al_u3276_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3277 (
    .a(_al_u3253_o),
    .b(_al_u3276_o),
    .c(data_csr[56]),
    .o(\cu_ru/m_cycle_event/n9 [56]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3278 (
    .a(\cu_ru/m_cycle_event/n2 [55]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [55]),
    .o(_al_u3278_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3279 (
    .a(_al_u3253_o),
    .b(_al_u3278_o),
    .c(data_csr[55]),
    .o(\cu_ru/m_cycle_event/n9 [55]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3280 (
    .a(\cu_ru/m_cycle_event/n2 [54]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [54]),
    .o(_al_u3280_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3281 (
    .a(_al_u3253_o),
    .b(_al_u3280_o),
    .c(data_csr[54]),
    .o(\cu_ru/m_cycle_event/n9 [54]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3282 (
    .a(\cu_ru/m_cycle_event/n2 [53]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [53]),
    .o(_al_u3282_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3283 (
    .a(_al_u3253_o),
    .b(_al_u3282_o),
    .c(data_csr[53]),
    .o(\cu_ru/m_cycle_event/n9 [53]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3284 (
    .a(\cu_ru/m_cycle_event/n2 [52]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [52]),
    .o(_al_u3284_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3285 (
    .a(_al_u3253_o),
    .b(_al_u3284_o),
    .c(data_csr[52]),
    .o(\cu_ru/m_cycle_event/n9 [52]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3286 (
    .a(\cu_ru/m_cycle_event/n2 [51]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [51]),
    .o(_al_u3286_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3287 (
    .a(_al_u3253_o),
    .b(_al_u3286_o),
    .c(data_csr[51]),
    .o(\cu_ru/m_cycle_event/n9 [51]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3288 (
    .a(\cu_ru/m_cycle_event/n2 [50]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [50]),
    .o(_al_u3288_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3289 (
    .a(_al_u3253_o),
    .b(_al_u3288_o),
    .c(data_csr[50]),
    .o(\cu_ru/m_cycle_event/n9 [50]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3290 (
    .a(\cu_ru/m_cycle_event/n2 [5]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [5]),
    .o(_al_u3290_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3291 (
    .a(_al_u3253_o),
    .b(_al_u3290_o),
    .c(data_csr[5]),
    .o(\cu_ru/m_cycle_event/n9 [5]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3292 (
    .a(\cu_ru/m_cycle_event/n2 [49]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [49]),
    .o(_al_u3292_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3293 (
    .a(_al_u3253_o),
    .b(_al_u3292_o),
    .c(data_csr[49]),
    .o(\cu_ru/m_cycle_event/n9 [49]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3294 (
    .a(\cu_ru/m_cycle_event/n2 [48]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [48]),
    .o(_al_u3294_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3295 (
    .a(_al_u3253_o),
    .b(_al_u3294_o),
    .c(data_csr[48]),
    .o(\cu_ru/m_cycle_event/n9 [48]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3296 (
    .a(\cu_ru/m_cycle_event/n2 [47]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [47]),
    .o(_al_u3296_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3297 (
    .a(_al_u3253_o),
    .b(_al_u3296_o),
    .c(data_csr[47]),
    .o(\cu_ru/m_cycle_event/n9 [47]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3298 (
    .a(\cu_ru/m_cycle_event/n2 [46]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [46]),
    .o(_al_u3298_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3299 (
    .a(_al_u3253_o),
    .b(_al_u3298_o),
    .c(data_csr[46]),
    .o(\cu_ru/m_cycle_event/n9 [46]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3300 (
    .a(\cu_ru/m_cycle_event/n2 [45]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [45]),
    .o(_al_u3300_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3301 (
    .a(_al_u3253_o),
    .b(_al_u3300_o),
    .c(data_csr[45]),
    .o(\cu_ru/m_cycle_event/n9 [45]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3302 (
    .a(\cu_ru/m_cycle_event/n2 [44]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [44]),
    .o(_al_u3302_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3303 (
    .a(_al_u3253_o),
    .b(_al_u3302_o),
    .c(data_csr[44]),
    .o(\cu_ru/m_cycle_event/n9 [44]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3304 (
    .a(\cu_ru/m_cycle_event/n2 [43]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [43]),
    .o(_al_u3304_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3305 (
    .a(_al_u3253_o),
    .b(_al_u3304_o),
    .c(data_csr[43]),
    .o(\cu_ru/m_cycle_event/n9 [43]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3306 (
    .a(\cu_ru/m_cycle_event/n2 [42]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [42]),
    .o(_al_u3306_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3307 (
    .a(_al_u3253_o),
    .b(_al_u3306_o),
    .c(data_csr[42]),
    .o(\cu_ru/m_cycle_event/n9 [42]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3308 (
    .a(\cu_ru/m_cycle_event/n2 [41]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [41]),
    .o(_al_u3308_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3309 (
    .a(_al_u3253_o),
    .b(_al_u3308_o),
    .c(data_csr[41]),
    .o(\cu_ru/m_cycle_event/n9 [41]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3310 (
    .a(\cu_ru/m_cycle_event/n2 [40]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [40]),
    .o(_al_u3310_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3311 (
    .a(_al_u3253_o),
    .b(_al_u3310_o),
    .c(data_csr[40]),
    .o(\cu_ru/m_cycle_event/n9 [40]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3312 (
    .a(\cu_ru/m_cycle_event/n2 [4]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [4]),
    .o(_al_u3312_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3313 (
    .a(_al_u3253_o),
    .b(_al_u3312_o),
    .c(data_csr[4]),
    .o(\cu_ru/m_cycle_event/n9 [4]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3314 (
    .a(\cu_ru/m_cycle_event/n2 [39]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [39]),
    .o(_al_u3314_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3315 (
    .a(_al_u3253_o),
    .b(_al_u3314_o),
    .c(data_csr[39]),
    .o(\cu_ru/m_cycle_event/n9 [39]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3316 (
    .a(\cu_ru/m_cycle_event/n2 [38]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [38]),
    .o(_al_u3316_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3317 (
    .a(_al_u3253_o),
    .b(_al_u3316_o),
    .c(data_csr[38]),
    .o(\cu_ru/m_cycle_event/n9 [38]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3318 (
    .a(\cu_ru/m_cycle_event/n2 [37]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [37]),
    .o(_al_u3318_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3319 (
    .a(_al_u3253_o),
    .b(_al_u3318_o),
    .c(data_csr[37]),
    .o(\cu_ru/m_cycle_event/n9 [37]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3320 (
    .a(\cu_ru/m_cycle_event/n2 [36]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [36]),
    .o(_al_u3320_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3321 (
    .a(_al_u3253_o),
    .b(_al_u3320_o),
    .c(data_csr[36]),
    .o(\cu_ru/m_cycle_event/n9 [36]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3322 (
    .a(\cu_ru/m_cycle_event/n2 [35]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [35]),
    .o(_al_u3322_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3323 (
    .a(_al_u3253_o),
    .b(_al_u3322_o),
    .c(data_csr[35]),
    .o(\cu_ru/m_cycle_event/n9 [35]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3324 (
    .a(\cu_ru/m_cycle_event/n2 [34]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [34]),
    .o(_al_u3324_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3325 (
    .a(_al_u3253_o),
    .b(_al_u3324_o),
    .c(data_csr[34]),
    .o(\cu_ru/m_cycle_event/n9 [34]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3326 (
    .a(\cu_ru/m_cycle_event/n2 [33]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [33]),
    .o(_al_u3326_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3327 (
    .a(_al_u3253_o),
    .b(_al_u3326_o),
    .c(data_csr[33]),
    .o(\cu_ru/m_cycle_event/n9 [33]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3328 (
    .a(\cu_ru/m_cycle_event/n2 [32]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [32]),
    .o(_al_u3328_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3329 (
    .a(_al_u3253_o),
    .b(_al_u3328_o),
    .c(data_csr[32]),
    .o(\cu_ru/m_cycle_event/n9 [32]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3330 (
    .a(\cu_ru/m_cycle_event/n2 [31]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [31]),
    .o(_al_u3330_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3331 (
    .a(_al_u3253_o),
    .b(_al_u3330_o),
    .c(data_csr[31]),
    .o(\cu_ru/m_cycle_event/n9 [31]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3332 (
    .a(\cu_ru/m_cycle_event/n2 [30]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [30]),
    .o(_al_u3332_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3333 (
    .a(_al_u3253_o),
    .b(_al_u3332_o),
    .c(data_csr[30]),
    .o(\cu_ru/m_cycle_event/n9 [30]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3334 (
    .a(\cu_ru/m_cycle_event/n2 [3]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [3]),
    .o(_al_u3334_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3335 (
    .a(_al_u3253_o),
    .b(_al_u3334_o),
    .c(data_csr[3]),
    .o(\cu_ru/m_cycle_event/n9 [3]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3336 (
    .a(\cu_ru/m_cycle_event/n2 [29]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [29]),
    .o(_al_u3336_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3337 (
    .a(_al_u3253_o),
    .b(_al_u3336_o),
    .c(data_csr[29]),
    .o(\cu_ru/m_cycle_event/n9 [29]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3338 (
    .a(\cu_ru/m_cycle_event/n2 [28]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [28]),
    .o(_al_u3338_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3339 (
    .a(_al_u3253_o),
    .b(_al_u3338_o),
    .c(data_csr[28]),
    .o(\cu_ru/m_cycle_event/n9 [28]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3340 (
    .a(\cu_ru/m_cycle_event/n2 [27]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [27]),
    .o(_al_u3340_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3341 (
    .a(_al_u3253_o),
    .b(_al_u3340_o),
    .c(data_csr[27]),
    .o(\cu_ru/m_cycle_event/n9 [27]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3342 (
    .a(\cu_ru/m_cycle_event/n2 [26]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [26]),
    .o(_al_u3342_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3343 (
    .a(_al_u3253_o),
    .b(_al_u3342_o),
    .c(data_csr[26]),
    .o(\cu_ru/m_cycle_event/n9 [26]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3344 (
    .a(\cu_ru/m_cycle_event/n2 [25]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [25]),
    .o(_al_u3344_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3345 (
    .a(_al_u3253_o),
    .b(_al_u3344_o),
    .c(data_csr[25]),
    .o(\cu_ru/m_cycle_event/n9 [25]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3346 (
    .a(\cu_ru/m_cycle_event/n2 [24]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [24]),
    .o(_al_u3346_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3347 (
    .a(_al_u3253_o),
    .b(_al_u3346_o),
    .c(data_csr[24]),
    .o(\cu_ru/m_cycle_event/n9 [24]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3348 (
    .a(\cu_ru/m_cycle_event/n2 [23]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [23]),
    .o(_al_u3348_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3349 (
    .a(_al_u3253_o),
    .b(_al_u3348_o),
    .c(data_csr[23]),
    .o(\cu_ru/m_cycle_event/n9 [23]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3350 (
    .a(\cu_ru/m_cycle_event/n2 [22]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [22]),
    .o(_al_u3350_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3351 (
    .a(_al_u3253_o),
    .b(_al_u3350_o),
    .c(data_csr[22]),
    .o(\cu_ru/m_cycle_event/n9 [22]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3352 (
    .a(\cu_ru/m_cycle_event/n2 [21]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [21]),
    .o(_al_u3352_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3353 (
    .a(_al_u3253_o),
    .b(_al_u3352_o),
    .c(data_csr[21]),
    .o(\cu_ru/m_cycle_event/n9 [21]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3354 (
    .a(\cu_ru/m_cycle_event/n2 [20]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [20]),
    .o(_al_u3354_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3355 (
    .a(_al_u3253_o),
    .b(_al_u3354_o),
    .c(data_csr[20]),
    .o(\cu_ru/m_cycle_event/n9 [20]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3356 (
    .a(\cu_ru/m_cycle_event/n2 [2]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [2]),
    .o(_al_u3356_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3357 (
    .a(_al_u3253_o),
    .b(_al_u3356_o),
    .c(data_csr[2]),
    .o(\cu_ru/m_cycle_event/n9 [2]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3358 (
    .a(\cu_ru/m_cycle_event/n2 [19]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [19]),
    .o(_al_u3358_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3359 (
    .a(_al_u3253_o),
    .b(_al_u3358_o),
    .c(data_csr[19]),
    .o(\cu_ru/m_cycle_event/n9 [19]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3360 (
    .a(\cu_ru/m_cycle_event/n2 [18]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [18]),
    .o(_al_u3360_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3361 (
    .a(_al_u3253_o),
    .b(_al_u3360_o),
    .c(data_csr[18]),
    .o(\cu_ru/m_cycle_event/n9 [18]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3362 (
    .a(\cu_ru/m_cycle_event/n2 [17]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [17]),
    .o(_al_u3362_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3363 (
    .a(_al_u3253_o),
    .b(_al_u3362_o),
    .c(data_csr[17]),
    .o(\cu_ru/m_cycle_event/n9 [17]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3364 (
    .a(\cu_ru/m_cycle_event/n2 [16]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [16]),
    .o(_al_u3364_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3365 (
    .a(_al_u3253_o),
    .b(_al_u3364_o),
    .c(data_csr[16]),
    .o(\cu_ru/m_cycle_event/n9 [16]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3366 (
    .a(\cu_ru/m_cycle_event/n2 [15]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [15]),
    .o(_al_u3366_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3367 (
    .a(_al_u3253_o),
    .b(_al_u3366_o),
    .c(data_csr[15]),
    .o(\cu_ru/m_cycle_event/n9 [15]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3368 (
    .a(\cu_ru/m_cycle_event/n2 [14]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [14]),
    .o(_al_u3368_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3369 (
    .a(_al_u3253_o),
    .b(_al_u3368_o),
    .c(data_csr[14]),
    .o(\cu_ru/m_cycle_event/n9 [14]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3370 (
    .a(\cu_ru/m_cycle_event/n2 [13]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [13]),
    .o(_al_u3370_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3371 (
    .a(_al_u3253_o),
    .b(_al_u3370_o),
    .c(data_csr[13]),
    .o(\cu_ru/m_cycle_event/n9 [13]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3372 (
    .a(\cu_ru/m_cycle_event/n2 [12]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [12]),
    .o(_al_u3372_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3373 (
    .a(_al_u3253_o),
    .b(_al_u3372_o),
    .c(data_csr[12]),
    .o(\cu_ru/m_cycle_event/n9 [12]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3374 (
    .a(\cu_ru/m_cycle_event/n2 [11]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [11]),
    .o(_al_u3374_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3375 (
    .a(_al_u3253_o),
    .b(_al_u3374_o),
    .c(data_csr[11]),
    .o(\cu_ru/m_cycle_event/n9 [11]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3376 (
    .a(\cu_ru/m_cycle_event/n2 [10]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [10]),
    .o(_al_u3376_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3377 (
    .a(_al_u3253_o),
    .b(_al_u3376_o),
    .c(data_csr[10]),
    .o(\cu_ru/m_cycle_event/n9 [10]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3378 (
    .a(\cu_ru/m_cycle_event/n2 [1]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [1]),
    .o(_al_u3378_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3379 (
    .a(_al_u3253_o),
    .b(_al_u3378_o),
    .c(data_csr[1]),
    .o(\cu_ru/m_cycle_event/n9 [1]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u3380 (
    .a(\cu_ru/m_cycle_event/n2 [0]),
    .b(\cu_ru/mcountinhibit ),
    .c(\cu_ru/mcycle [0]),
    .o(_al_u3380_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u3381 (
    .a(_al_u3253_o),
    .b(_al_u3380_o),
    .c(data_csr[0]),
    .o(\cu_ru/m_cycle_event/n9 [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3382 (
    .a(_al_u2933_o),
    .b(_al_u2938_o),
    .c(_al_u3212_o),
    .o(_al_u3382_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u3383 (
    .a(_al_u3214_o),
    .b(_al_u3382_o),
    .o(\ins_dec/n302 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u3384 (
    .a(\ins_fetch/ins_shift [12]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [12]),
    .o(_al_u3384_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3385 (
    .a(id_system),
    .b(_al_u3217_o),
    .c(_al_u3384_o),
    .o(\ins_dec/n71 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3386 (
    .a(id_ins[29]),
    .b(id_ins[28]),
    .o(\ins_dec/n80_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(~B*~A))"),
    .INIT(16'heee0))
    _al_u3387 (
    .a(_al_u2667_o),
    .b(_al_u2668_o),
    .c(_al_u2670_o),
    .d(_al_u2671_o),
    .o(_al_u3387_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(~B*~A))"),
    .INIT(16'heee0))
    _al_u3388 (
    .a(_al_u2659_o),
    .b(_al_u2660_o),
    .c(_al_u2662_o),
    .d(_al_u2663_o),
    .o(_al_u3388_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3389 (
    .a(\ins_dec/n80_lutinv ),
    .b(_al_u3387_o),
    .c(_al_u3388_o),
    .o(\ins_dec/funct6_0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3390 (
    .a(\ins_dec/n35_lutinv ),
    .b(_al_u3384_o),
    .o(\ins_dec/funct3_0_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3391 (
    .a(\ins_dec/funct6_0_lutinv ),
    .b(\ins_dec/funct3_0_lutinv ),
    .c(id_system),
    .o(_al_u3391_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(~B*~A))"),
    .INIT(16'heee0))
    _al_u3392 (
    .a(_al_u2674_o),
    .b(_al_u2675_o),
    .c(_al_u2677_o),
    .d(_al_u2678_o),
    .o(_al_u3392_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3393 (
    .a(id_ins[25]),
    .b(_al_u3392_o),
    .o(_al_u3393_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(~B*~A))"),
    .INIT(16'heee0))
    _al_u3394 (
    .a(_al_u2680_o),
    .b(_al_u2681_o),
    .c(_al_u2683_o),
    .d(_al_u2684_o),
    .o(_al_u3394_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3395 (
    .a(_al_u3393_o),
    .b(id_ins[20]),
    .c(_al_u3394_o),
    .o(_al_u3395_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3396 (
    .a(_al_u3391_o),
    .b(_al_u3395_o),
    .o(\ins_dec/ins_ebreak ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u3397 (
    .a(id_ins[25]),
    .b(id_ins[20]),
    .c(_al_u3394_o),
    .d(_al_u3392_o),
    .o(_al_u3397_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3398 (
    .a(_al_u3391_o),
    .b(_al_u3397_o),
    .o(\ins_dec/ins_ecall ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3399 (
    .a(id_ins[29]),
    .b(_al_u3388_o),
    .o(_al_u3399_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3400 (
    .a(id_ins[28]),
    .b(_al_u3387_o),
    .o(_al_u3400_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3401 (
    .a(id_system),
    .b(_al_u3399_o),
    .c(_al_u3400_o),
    .d(id_ins[25]),
    .o(\ins_dec/ins_sfencevma ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u3402 (
    .a(\ins_dec/ins_fence ),
    .b(\ins_dec/ins_sfencevma ),
    .o(\ins_dec/n225 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3403 (
    .a(_al_u2703_o),
    .b(\biu/bus_unit/statu [0]),
    .c(\biu/bus_unit/statu [1]),
    .d(\biu/bus_unit/statu [3]),
    .o(_al_u3403_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3404 (
    .a(_al_u2955_o),
    .b(\biu/bus_unit/statu [0]),
    .c(\biu/bus_unit/statu [1]),
    .o(_al_u3404_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3405 (
    .a(_al_u3403_o),
    .b(_al_u3404_o),
    .o(\biu/bus_unit/mux10_b3_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u3406 (
    .a(\biu/bus_unit/mux10_b3_sel_is_0_o ),
    .b(_al_u2703_o),
    .c(\biu/bus_unit/statu [1]),
    .d(\biu/bus_unit/statu [3]),
    .o(\biu/bus_unit/mux11_b4_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3407 (
    .a(_al_u2889_o),
    .b(\biu/bus_unit/statu [2]),
    .c(\biu/bus_unit/statu [4]),
    .o(_al_u3407_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    .INIT(16'h7250))
    _al_u3408 (
    .a(\biu/bus_unit/mux11_b4_sel_is_2_o ),
    .b(_al_u3407_o),
    .c(hresp_pad),
    .d(\biu/bus_unit/statu [4]),
    .o(\biu/bus_unit/n30 [4]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u3409 (
    .a(_al_u2703_o),
    .b(\biu/bus_unit/statu [0]),
    .c(\biu/bus_unit/statu [1]),
    .d(\biu/bus_unit/statu [3]),
    .o(\biu/bus_unit/n45_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3410 (
    .a(\biu/bus_unit/mux10_b3_sel_is_0_o ),
    .b(_al_u2890_o),
    .c(\biu/bus_unit/n45_lutinv ),
    .o(_al_u3410_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u3411 (
    .a(\biu/bus_unit/mmu/statu [0]),
    .b(\biu/bus_unit/mmu/statu [1]),
    .c(\biu/bus_unit/mmu/statu [2]),
    .d(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u3411_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(C)*~(B)+(D*~A)*C*~(B)+~((D*~A))*C*B+(D*~A)*C*B)"),
    .INIT(16'h2e3f))
    _al_u3412 (
    .a(_al_u3410_o),
    .b(_al_u2705_o),
    .c(_al_u3411_o),
    .d(hready_pad),
    .o(\biu/cache_ctrl_logic/n100 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3413 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ),
    .o(\biu/cache_ctrl_logic/n149 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3414 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u2886_o),
    .o(\biu/cache_ctrl_logic/n135 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3415 (
    .a(ex_size[0]),
    .b(ex_size[1]),
    .o(_al_u3415_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u3416 (
    .a(_al_u2706_o),
    .b(_al_u3415_o),
    .o(hsize_pad[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3417 (
    .a(\biu/bus_unit/n37 ),
    .b(\biu/bus_unit/mux15_b4_sel_is_2_o ),
    .o(\biu/bus_unit/mux17_b4_sel_is_2_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3418 (
    .a(_al_u3181_o),
    .b(store),
    .o(\exu/store_addr_mis ));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u3419 (
    .a(\exu/load_addr_mis ),
    .b(\exu/store_addr_mis ),
    .c(_al_u2910_o),
    .o(\exu/n88 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3420 (
    .a(_al_u3186_o),
    .b(csr_index[6]),
    .c(csr_index[7]),
    .d(csr_index[8]),
    .o(_al_u3420_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3421 (
    .a(_al_u3191_o),
    .b(_al_u3420_o),
    .o(\cu_ru/m_s_ip/u12_sel_is_2_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3422 (
    .a(\cu_ru/m_s_ip/n0 ),
    .b(\cu_ru/m_s_ip/u12_sel_is_2_o ),
    .o(\cu_ru/m_s_ip/u11_sel_is_0_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3423 (
    .a(_al_u3185_o),
    .b(_al_u3420_o),
    .o(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3424 (
    .a(_al_u3253_o),
    .b(\cu_ru/m_cycle_event/mcountinhibit[2] ),
    .c(wb_valid),
    .o(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3425 (
    .a(_al_u3201_o),
    .b(_al_u3186_o),
    .c(_al_u3194_o),
    .o(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*A)"),
    .INIT(16'hfff7))
    _al_u3426 (
    .a(_al_u3191_o),
    .b(_al_u3194_o),
    .c(csr_index[10]),
    .d(csr_index[11]),
    .o(\cu_ru/m_s_ie/u11_sel_is_0_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3427 (
    .a(_al_u3185_o),
    .b(_al_u3186_o),
    .c(_al_u3194_o),
    .o(_al_u3427_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3428 (
    .a(\cu_ru/m_s_status/n0 ),
    .b(_al_u3427_o),
    .o(\cu_ru/m_s_status/u34_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C))"),
    .INIT(16'h00b2))
    _al_u3429 (
    .a(\exu/alu_au/n12 ),
    .b(ds1[63]),
    .c(ds2[63]),
    .d(unsign),
    .o(\exu/alu_au/n15 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u3430 (
    .a(\exu/alu_au/n15 ),
    .b(\exu/alu_au/n5 ),
    .c(unsign),
    .o(_al_u3430_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3431 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[9]),
    .d(ds2[9]),
    .o(\exu/alu_au/n53 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3432 (
    .a(\exu/alu_au/add_64 [9]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[9]),
    .o(_al_u3432_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3433 (
    .a(_al_u3432_o),
    .b(mem_csr_data_or),
    .c(ds1[9]),
    .d(ds2[9]),
    .o(_al_u3433_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3434 (
    .a(_al_u3433_o),
    .b(mem_csr_data_xor),
    .c(ds1[9]),
    .d(ds2[9]),
    .o(_al_u3434_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haa8e))
    _al_u3435 (
    .a(\exu/alu_au/n5 ),
    .b(ds1[63]),
    .c(ds2[63]),
    .d(unsign),
    .o(\exu/alu_au/ds1_light_than_ds2_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3436 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[9]),
    .d(ds2[9]),
    .o(\exu/alu_au/n55 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    _al_u3437 (
    .a(and_clr),
    .b(ds1[9]),
    .c(ds2[9]),
    .o(\exu/alu_au/alu_and [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3438 (
    .a(\exu/alu_au/alu_and [9]),
    .b(mem_csr_data_and),
    .o(\exu/alu_au/n47 [9]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3439 (
    .a(\exu/alu_au/n53 [9]),
    .b(_al_u3434_o),
    .c(\exu/alu_au/n55 [9]),
    .d(\exu/alu_au/n47 [9]),
    .o(\exu/alu_data_mem_csr [9]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3440 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[8]),
    .d(ds2[8]),
    .o(\exu/alu_au/n53 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3441 (
    .a(\exu/alu_au/add_64 [8]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[8]),
    .o(_al_u3441_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3442 (
    .a(_al_u3441_o),
    .b(mem_csr_data_or),
    .c(ds1[8]),
    .d(ds2[8]),
    .o(_al_u3442_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3443 (
    .a(_al_u3442_o),
    .b(mem_csr_data_xor),
    .c(ds1[8]),
    .d(ds2[8]),
    .o(_al_u3443_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3444 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[8]),
    .d(ds2[8]),
    .o(\exu/alu_au/n55 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    _al_u3445 (
    .a(and_clr),
    .b(ds1[8]),
    .c(ds2[8]),
    .o(\exu/alu_au/alu_and [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3446 (
    .a(\exu/alu_au/alu_and [8]),
    .b(mem_csr_data_and),
    .o(\exu/alu_au/n47 [8]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3447 (
    .a(\exu/alu_au/n53 [8]),
    .b(_al_u3443_o),
    .c(\exu/alu_au/n55 [8]),
    .d(\exu/alu_au/n47 [8]),
    .o(\exu/alu_data_mem_csr [8]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3448 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[7]),
    .d(ds2[7]),
    .o(\exu/alu_au/n53 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3449 (
    .a(\exu/alu_au/add_64 [7]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[7]),
    .o(_al_u3449_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3450 (
    .a(_al_u3449_o),
    .b(mem_csr_data_or),
    .c(ds1[7]),
    .d(ds2[7]),
    .o(_al_u3450_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3451 (
    .a(_al_u3450_o),
    .b(mem_csr_data_xor),
    .c(ds1[7]),
    .d(ds2[7]),
    .o(_al_u3451_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3452 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[7]),
    .d(ds2[7]),
    .o(\exu/alu_au/n55 [7]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3453 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[7]),
    .d(ds2[7]),
    .o(\exu/alu_au/n47 [7]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3454 (
    .a(\exu/alu_au/n53 [7]),
    .b(_al_u3451_o),
    .c(\exu/alu_au/n55 [7]),
    .d(\exu/alu_au/n47 [7]),
    .o(\exu/alu_data_mem_csr [7]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3455 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[63]),
    .d(ds2[63]),
    .o(\exu/alu_au/n53 [63]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h113f))
    _al_u3456 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds1[63]),
    .d(ds2[63]),
    .o(_al_u3456_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3457 (
    .a(_al_u3456_o),
    .b(mem_csr_data_xor),
    .c(ds1[63]),
    .d(ds2[63]),
    .o(_al_u3457_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3458 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[63]),
    .d(ds2[63]),
    .o(\exu/alu_au/n47 [63]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3459 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [63]),
    .c(ex_size[2]),
    .o(_al_u3459_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*~C))"),
    .INIT(16'h2022))
    _al_u3460 (
    .a(_al_u3457_o),
    .b(\exu/alu_au/n47 [63]),
    .c(_al_u3459_o),
    .d(mem_csr_data_add),
    .o(_al_u3460_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3461 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[63]),
    .d(ds2[63]),
    .o(\exu/alu_au/n55 [63]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3462 (
    .a(\exu/alu_au/n53 [63]),
    .b(_al_u3460_o),
    .c(\exu/alu_au/n55 [63]),
    .o(\exu/alu_data_mem_csr [63]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3463 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[62]),
    .d(ds2[62]),
    .o(\exu/alu_au/n53 [62]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3464 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[62]),
    .o(_al_u3464_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3465 (
    .a(_al_u3464_o),
    .b(mem_csr_data_xor),
    .c(ds1[62]),
    .d(ds2[62]),
    .o(_al_u3465_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3466 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[62]),
    .d(ds2[62]),
    .o(\exu/alu_au/n47 [62]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3467 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [62]),
    .c(ex_size[2]),
    .o(_al_u3467_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3468 (
    .a(_al_u3465_o),
    .b(\exu/alu_au/n47 [62]),
    .c(_al_u3467_o),
    .d(mem_csr_data_add),
    .o(_al_u3468_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3469 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[62]),
    .d(ds2[62]),
    .o(\exu/alu_au/n55 [62]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3470 (
    .a(\exu/alu_au/n53 [62]),
    .b(_al_u3468_o),
    .c(\exu/alu_au/n55 [62]),
    .o(\exu/alu_data_mem_csr [62]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3471 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[61]),
    .d(ds2[61]),
    .o(\exu/alu_au/n53 [61]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3472 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[61]),
    .o(_al_u3472_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3473 (
    .a(_al_u3472_o),
    .b(mem_csr_data_xor),
    .c(ds1[61]),
    .d(ds2[61]),
    .o(_al_u3473_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3474 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[61]),
    .d(ds2[61]),
    .o(\exu/alu_au/n47 [61]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3475 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [61]),
    .c(ex_size[2]),
    .o(_al_u3475_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3476 (
    .a(_al_u3473_o),
    .b(\exu/alu_au/n47 [61]),
    .c(_al_u3475_o),
    .d(mem_csr_data_add),
    .o(_al_u3476_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3477 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[61]),
    .d(ds2[61]),
    .o(\exu/alu_au/n55 [61]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3478 (
    .a(\exu/alu_au/n53 [61]),
    .b(_al_u3476_o),
    .c(\exu/alu_au/n55 [61]),
    .o(\exu/alu_data_mem_csr [61]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3479 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[60]),
    .d(ds2[60]),
    .o(\exu/alu_au/n53 [60]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3480 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[60]),
    .o(_al_u3480_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3481 (
    .a(_al_u3480_o),
    .b(mem_csr_data_xor),
    .c(ds1[60]),
    .d(ds2[60]),
    .o(_al_u3481_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3482 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[60]),
    .d(ds2[60]),
    .o(\exu/alu_au/n47 [60]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3483 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [60]),
    .c(ex_size[2]),
    .o(_al_u3483_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3484 (
    .a(_al_u3481_o),
    .b(\exu/alu_au/n47 [60]),
    .c(_al_u3483_o),
    .d(mem_csr_data_add),
    .o(_al_u3484_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3485 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[60]),
    .d(ds2[60]),
    .o(\exu/alu_au/n55 [60]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3486 (
    .a(\exu/alu_au/n53 [60]),
    .b(_al_u3484_o),
    .c(\exu/alu_au/n55 [60]),
    .o(\exu/alu_data_mem_csr [60]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3487 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[6]),
    .d(ds2[6]),
    .o(\exu/alu_au/n53 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3488 (
    .a(\exu/alu_au/add_64 [6]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[6]),
    .o(_al_u3488_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3489 (
    .a(_al_u3488_o),
    .b(mem_csr_data_or),
    .c(ds1[6]),
    .d(ds2[6]),
    .o(_al_u3489_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3490 (
    .a(_al_u3489_o),
    .b(mem_csr_data_xor),
    .c(ds1[6]),
    .d(ds2[6]),
    .o(_al_u3490_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3491 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[6]),
    .d(ds2[6]),
    .o(\exu/alu_au/n55 [6]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3492 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[6]),
    .d(ds2[6]),
    .o(\exu/alu_au/n47 [6]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3493 (
    .a(\exu/alu_au/n53 [6]),
    .b(_al_u3490_o),
    .c(\exu/alu_au/n55 [6]),
    .d(\exu/alu_au/n47 [6]),
    .o(\exu/alu_data_mem_csr [6]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3494 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[59]),
    .d(ds2[59]),
    .o(\exu/alu_au/n53 [59]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3495 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[59]),
    .o(_al_u3495_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3496 (
    .a(_al_u3495_o),
    .b(mem_csr_data_xor),
    .c(ds1[59]),
    .d(ds2[59]),
    .o(_al_u3496_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3497 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[59]),
    .d(ds2[59]),
    .o(\exu/alu_au/n47 [59]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3498 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [59]),
    .c(ex_size[2]),
    .o(_al_u3498_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3499 (
    .a(_al_u3496_o),
    .b(\exu/alu_au/n47 [59]),
    .c(_al_u3498_o),
    .d(mem_csr_data_add),
    .o(_al_u3499_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3500 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[59]),
    .d(ds2[59]),
    .o(\exu/alu_au/n55 [59]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3501 (
    .a(\exu/alu_au/n53 [59]),
    .b(_al_u3499_o),
    .c(\exu/alu_au/n55 [59]),
    .o(\exu/alu_data_mem_csr [59]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3502 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[58]),
    .d(ds2[58]),
    .o(\exu/alu_au/n53 [58]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3503 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[58]),
    .o(_al_u3503_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3504 (
    .a(_al_u3503_o),
    .b(mem_csr_data_xor),
    .c(ds1[58]),
    .d(ds2[58]),
    .o(_al_u3504_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3505 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[58]),
    .d(ds2[58]),
    .o(\exu/alu_au/n47 [58]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3506 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [58]),
    .c(ex_size[2]),
    .o(_al_u3506_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3507 (
    .a(_al_u3504_o),
    .b(\exu/alu_au/n47 [58]),
    .c(_al_u3506_o),
    .d(mem_csr_data_add),
    .o(_al_u3507_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3508 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[58]),
    .d(ds2[58]),
    .o(\exu/alu_au/n55 [58]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3509 (
    .a(\exu/alu_au/n53 [58]),
    .b(_al_u3507_o),
    .c(\exu/alu_au/n55 [58]),
    .o(\exu/alu_data_mem_csr [58]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3510 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[57]),
    .d(ds2[57]),
    .o(\exu/alu_au/n53 [57]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3511 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[57]),
    .o(_al_u3511_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3512 (
    .a(_al_u3511_o),
    .b(mem_csr_data_xor),
    .c(ds1[57]),
    .d(ds2[57]),
    .o(_al_u3512_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3513 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[57]),
    .d(ds2[57]),
    .o(\exu/alu_au/n47 [57]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3514 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [57]),
    .c(ex_size[2]),
    .o(_al_u3514_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3515 (
    .a(_al_u3512_o),
    .b(\exu/alu_au/n47 [57]),
    .c(_al_u3514_o),
    .d(mem_csr_data_add),
    .o(_al_u3515_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3516 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[57]),
    .d(ds2[57]),
    .o(\exu/alu_au/n55 [57]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3517 (
    .a(\exu/alu_au/n53 [57]),
    .b(_al_u3515_o),
    .c(\exu/alu_au/n55 [57]),
    .o(\exu/alu_data_mem_csr [57]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3518 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[56]),
    .d(ds2[56]),
    .o(\exu/alu_au/n53 [56]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3519 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[56]),
    .o(_al_u3519_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3520 (
    .a(_al_u3519_o),
    .b(mem_csr_data_xor),
    .c(ds1[56]),
    .d(ds2[56]),
    .o(_al_u3520_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3521 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[56]),
    .d(ds2[56]),
    .o(\exu/alu_au/n47 [56]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3522 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [56]),
    .c(ex_size[2]),
    .o(_al_u3522_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3523 (
    .a(_al_u3520_o),
    .b(\exu/alu_au/n47 [56]),
    .c(_al_u3522_o),
    .d(mem_csr_data_add),
    .o(_al_u3523_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3524 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[56]),
    .d(ds2[56]),
    .o(\exu/alu_au/n55 [56]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3525 (
    .a(\exu/alu_au/n53 [56]),
    .b(_al_u3523_o),
    .c(\exu/alu_au/n55 [56]),
    .o(\exu/alu_data_mem_csr [56]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3526 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[55]),
    .d(ds2[55]),
    .o(\exu/alu_au/n53 [55]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3527 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[55]),
    .o(_al_u3527_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3528 (
    .a(_al_u3527_o),
    .b(mem_csr_data_xor),
    .c(ds1[55]),
    .d(ds2[55]),
    .o(_al_u3528_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3529 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[55]),
    .d(ds2[55]),
    .o(\exu/alu_au/n47 [55]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3530 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [55]),
    .c(ex_size[2]),
    .o(_al_u3530_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3531 (
    .a(_al_u3528_o),
    .b(\exu/alu_au/n47 [55]),
    .c(_al_u3530_o),
    .d(mem_csr_data_add),
    .o(_al_u3531_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3532 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[55]),
    .d(ds2[55]),
    .o(\exu/alu_au/n55 [55]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3533 (
    .a(\exu/alu_au/n53 [55]),
    .b(_al_u3531_o),
    .c(\exu/alu_au/n55 [55]),
    .o(\exu/alu_data_mem_csr [55]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3534 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[54]),
    .d(ds2[54]),
    .o(\exu/alu_au/n53 [54]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3535 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[54]),
    .o(_al_u3535_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3536 (
    .a(_al_u3535_o),
    .b(mem_csr_data_xor),
    .c(ds1[54]),
    .d(ds2[54]),
    .o(_al_u3536_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3537 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[54]),
    .d(ds2[54]),
    .o(\exu/alu_au/n47 [54]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3538 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [54]),
    .c(ex_size[2]),
    .o(_al_u3538_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3539 (
    .a(_al_u3536_o),
    .b(\exu/alu_au/n47 [54]),
    .c(_al_u3538_o),
    .d(mem_csr_data_add),
    .o(_al_u3539_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3540 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[54]),
    .d(ds2[54]),
    .o(\exu/alu_au/n55 [54]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3541 (
    .a(\exu/alu_au/n53 [54]),
    .b(_al_u3539_o),
    .c(\exu/alu_au/n55 [54]),
    .o(\exu/alu_data_mem_csr [54]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3542 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[53]),
    .d(ds2[53]),
    .o(\exu/alu_au/n53 [53]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3543 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[53]),
    .o(_al_u3543_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3544 (
    .a(_al_u3543_o),
    .b(mem_csr_data_xor),
    .c(ds1[53]),
    .d(ds2[53]),
    .o(_al_u3544_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3545 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[53]),
    .d(ds2[53]),
    .o(\exu/alu_au/n47 [53]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3546 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [53]),
    .c(ex_size[2]),
    .o(_al_u3546_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3547 (
    .a(_al_u3544_o),
    .b(\exu/alu_au/n47 [53]),
    .c(_al_u3546_o),
    .d(mem_csr_data_add),
    .o(_al_u3547_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3548 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[53]),
    .d(ds2[53]),
    .o(\exu/alu_au/n55 [53]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3549 (
    .a(\exu/alu_au/n53 [53]),
    .b(_al_u3547_o),
    .c(\exu/alu_au/n55 [53]),
    .o(\exu/alu_data_mem_csr [53]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3550 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[52]),
    .d(ds2[52]),
    .o(\exu/alu_au/n53 [52]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3551 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[52]),
    .o(_al_u3551_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3552 (
    .a(_al_u3551_o),
    .b(mem_csr_data_xor),
    .c(ds1[52]),
    .d(ds2[52]),
    .o(_al_u3552_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3553 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[52]),
    .d(ds2[52]),
    .o(\exu/alu_au/n47 [52]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3554 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [52]),
    .c(ex_size[2]),
    .o(_al_u3554_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3555 (
    .a(_al_u3552_o),
    .b(\exu/alu_au/n47 [52]),
    .c(_al_u3554_o),
    .d(mem_csr_data_add),
    .o(_al_u3555_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3556 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[52]),
    .d(ds2[52]),
    .o(\exu/alu_au/n55 [52]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3557 (
    .a(\exu/alu_au/n53 [52]),
    .b(_al_u3555_o),
    .c(\exu/alu_au/n55 [52]),
    .o(\exu/alu_data_mem_csr [52]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3558 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[51]),
    .d(ds2[51]),
    .o(\exu/alu_au/n53 [51]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3559 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[51]),
    .o(_al_u3559_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3560 (
    .a(_al_u3559_o),
    .b(mem_csr_data_xor),
    .c(ds1[51]),
    .d(ds2[51]),
    .o(_al_u3560_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3561 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[51]),
    .d(ds2[51]),
    .o(\exu/alu_au/n47 [51]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3562 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [51]),
    .c(ex_size[2]),
    .o(_al_u3562_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3563 (
    .a(_al_u3560_o),
    .b(\exu/alu_au/n47 [51]),
    .c(_al_u3562_o),
    .d(mem_csr_data_add),
    .o(_al_u3563_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3564 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[51]),
    .d(ds2[51]),
    .o(\exu/alu_au/n55 [51]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3565 (
    .a(\exu/alu_au/n53 [51]),
    .b(_al_u3563_o),
    .c(\exu/alu_au/n55 [51]),
    .o(\exu/alu_data_mem_csr [51]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3566 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[50]),
    .d(ds2[50]),
    .o(\exu/alu_au/n53 [50]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3567 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[50]),
    .o(_al_u3567_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3568 (
    .a(_al_u3567_o),
    .b(mem_csr_data_xor),
    .c(ds1[50]),
    .d(ds2[50]),
    .o(_al_u3568_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3569 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[50]),
    .d(ds2[50]),
    .o(\exu/alu_au/n47 [50]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3570 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [50]),
    .c(ex_size[2]),
    .o(_al_u3570_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3571 (
    .a(_al_u3568_o),
    .b(\exu/alu_au/n47 [50]),
    .c(_al_u3570_o),
    .d(mem_csr_data_add),
    .o(_al_u3571_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3572 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[50]),
    .d(ds2[50]),
    .o(\exu/alu_au/n55 [50]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3573 (
    .a(\exu/alu_au/n53 [50]),
    .b(_al_u3571_o),
    .c(\exu/alu_au/n55 [50]),
    .o(\exu/alu_data_mem_csr [50]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3574 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[5]),
    .d(ds2[5]),
    .o(\exu/alu_au/n53 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3575 (
    .a(\exu/alu_au/add_64 [5]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[5]),
    .o(_al_u3575_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3576 (
    .a(_al_u3575_o),
    .b(mem_csr_data_or),
    .c(ds1[5]),
    .d(ds2[5]),
    .o(_al_u3576_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3577 (
    .a(_al_u3576_o),
    .b(mem_csr_data_xor),
    .c(ds1[5]),
    .d(ds2[5]),
    .o(_al_u3577_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3578 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[5]),
    .d(ds2[5]),
    .o(\exu/alu_au/n55 [5]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3579 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[5]),
    .d(ds2[5]),
    .o(\exu/alu_au/n47 [5]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3580 (
    .a(\exu/alu_au/n53 [5]),
    .b(_al_u3577_o),
    .c(\exu/alu_au/n55 [5]),
    .d(\exu/alu_au/n47 [5]),
    .o(\exu/alu_data_mem_csr [5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3581 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[49]),
    .d(ds2[49]),
    .o(\exu/alu_au/n53 [49]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3582 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[49]),
    .o(_al_u3582_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3583 (
    .a(_al_u3582_o),
    .b(mem_csr_data_xor),
    .c(ds1[49]),
    .d(ds2[49]),
    .o(_al_u3583_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3584 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[49]),
    .d(ds2[49]),
    .o(\exu/alu_au/n47 [49]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3585 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [49]),
    .c(ex_size[2]),
    .o(_al_u3585_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3586 (
    .a(_al_u3583_o),
    .b(\exu/alu_au/n47 [49]),
    .c(_al_u3585_o),
    .d(mem_csr_data_add),
    .o(_al_u3586_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3587 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[49]),
    .d(ds2[49]),
    .o(\exu/alu_au/n55 [49]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3588 (
    .a(\exu/alu_au/n53 [49]),
    .b(_al_u3586_o),
    .c(\exu/alu_au/n55 [49]),
    .o(\exu/alu_data_mem_csr [49]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3589 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[48]),
    .d(ds2[48]),
    .o(\exu/alu_au/n53 [48]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3590 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[48]),
    .o(_al_u3590_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3591 (
    .a(_al_u3590_o),
    .b(mem_csr_data_xor),
    .c(ds1[48]),
    .d(ds2[48]),
    .o(_al_u3591_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3592 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[48]),
    .d(ds2[48]),
    .o(\exu/alu_au/n47 [48]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3593 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [48]),
    .c(ex_size[2]),
    .o(_al_u3593_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3594 (
    .a(_al_u3591_o),
    .b(\exu/alu_au/n47 [48]),
    .c(_al_u3593_o),
    .d(mem_csr_data_add),
    .o(_al_u3594_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3595 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[48]),
    .d(ds2[48]),
    .o(\exu/alu_au/n55 [48]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3596 (
    .a(\exu/alu_au/n53 [48]),
    .b(_al_u3594_o),
    .c(\exu/alu_au/n55 [48]),
    .o(\exu/alu_data_mem_csr [48]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3597 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[47]),
    .d(ds2[47]),
    .o(\exu/alu_au/n53 [47]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3598 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[47]),
    .o(_al_u3598_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3599 (
    .a(_al_u3598_o),
    .b(mem_csr_data_xor),
    .c(ds1[47]),
    .d(ds2[47]),
    .o(_al_u3599_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3600 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[47]),
    .d(ds2[47]),
    .o(\exu/alu_au/n47 [47]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3601 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [47]),
    .c(ex_size[2]),
    .o(_al_u3601_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3602 (
    .a(_al_u3599_o),
    .b(\exu/alu_au/n47 [47]),
    .c(_al_u3601_o),
    .d(mem_csr_data_add),
    .o(_al_u3602_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3603 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[47]),
    .d(ds2[47]),
    .o(\exu/alu_au/n55 [47]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3604 (
    .a(\exu/alu_au/n53 [47]),
    .b(_al_u3602_o),
    .c(\exu/alu_au/n55 [47]),
    .o(\exu/alu_data_mem_csr [47]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3605 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[46]),
    .d(ds2[46]),
    .o(\exu/alu_au/n53 [46]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3606 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[46]),
    .o(_al_u3606_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3607 (
    .a(_al_u3606_o),
    .b(mem_csr_data_xor),
    .c(ds1[46]),
    .d(ds2[46]),
    .o(_al_u3607_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3608 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[46]),
    .d(ds2[46]),
    .o(\exu/alu_au/n47 [46]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3609 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [46]),
    .c(ex_size[2]),
    .o(_al_u3609_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3610 (
    .a(_al_u3607_o),
    .b(\exu/alu_au/n47 [46]),
    .c(_al_u3609_o),
    .d(mem_csr_data_add),
    .o(_al_u3610_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3611 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[46]),
    .d(ds2[46]),
    .o(\exu/alu_au/n55 [46]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3612 (
    .a(\exu/alu_au/n53 [46]),
    .b(_al_u3610_o),
    .c(\exu/alu_au/n55 [46]),
    .o(\exu/alu_data_mem_csr [46]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3613 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[45]),
    .d(ds2[45]),
    .o(\exu/alu_au/n53 [45]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3614 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[45]),
    .o(_al_u3614_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3615 (
    .a(_al_u3614_o),
    .b(mem_csr_data_xor),
    .c(ds1[45]),
    .d(ds2[45]),
    .o(_al_u3615_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3616 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[45]),
    .d(ds2[45]),
    .o(\exu/alu_au/n47 [45]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3617 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [45]),
    .c(ex_size[2]),
    .o(_al_u3617_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3618 (
    .a(_al_u3615_o),
    .b(\exu/alu_au/n47 [45]),
    .c(_al_u3617_o),
    .d(mem_csr_data_add),
    .o(_al_u3618_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3619 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[45]),
    .d(ds2[45]),
    .o(\exu/alu_au/n55 [45]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3620 (
    .a(\exu/alu_au/n53 [45]),
    .b(_al_u3618_o),
    .c(\exu/alu_au/n55 [45]),
    .o(\exu/alu_data_mem_csr [45]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3621 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[44]),
    .d(ds2[44]),
    .o(\exu/alu_au/n53 [44]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3622 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[44]),
    .o(_al_u3622_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3623 (
    .a(_al_u3622_o),
    .b(mem_csr_data_xor),
    .c(ds1[44]),
    .d(ds2[44]),
    .o(_al_u3623_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3624 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[44]),
    .d(ds2[44]),
    .o(\exu/alu_au/n47 [44]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3625 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [44]),
    .c(ex_size[2]),
    .o(_al_u3625_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3626 (
    .a(_al_u3623_o),
    .b(\exu/alu_au/n47 [44]),
    .c(_al_u3625_o),
    .d(mem_csr_data_add),
    .o(_al_u3626_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3627 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[44]),
    .d(ds2[44]),
    .o(\exu/alu_au/n55 [44]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3628 (
    .a(\exu/alu_au/n53 [44]),
    .b(_al_u3626_o),
    .c(\exu/alu_au/n55 [44]),
    .o(\exu/alu_data_mem_csr [44]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3629 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[43]),
    .d(ds2[43]),
    .o(\exu/alu_au/n53 [43]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3630 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[43]),
    .o(_al_u3630_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3631 (
    .a(_al_u3630_o),
    .b(mem_csr_data_xor),
    .c(ds1[43]),
    .d(ds2[43]),
    .o(_al_u3631_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3632 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[43]),
    .d(ds2[43]),
    .o(\exu/alu_au/n47 [43]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3633 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [43]),
    .c(ex_size[2]),
    .o(_al_u3633_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3634 (
    .a(_al_u3631_o),
    .b(\exu/alu_au/n47 [43]),
    .c(_al_u3633_o),
    .d(mem_csr_data_add),
    .o(_al_u3634_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3635 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[43]),
    .d(ds2[43]),
    .o(\exu/alu_au/n55 [43]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3636 (
    .a(\exu/alu_au/n53 [43]),
    .b(_al_u3634_o),
    .c(\exu/alu_au/n55 [43]),
    .o(\exu/alu_data_mem_csr [43]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3637 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[42]),
    .d(ds2[42]),
    .o(\exu/alu_au/n53 [42]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3638 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[42]),
    .o(_al_u3638_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3639 (
    .a(_al_u3638_o),
    .b(mem_csr_data_xor),
    .c(ds1[42]),
    .d(ds2[42]),
    .o(_al_u3639_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3640 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[42]),
    .d(ds2[42]),
    .o(\exu/alu_au/n47 [42]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3641 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [42]),
    .c(ex_size[2]),
    .o(_al_u3641_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3642 (
    .a(_al_u3639_o),
    .b(\exu/alu_au/n47 [42]),
    .c(_al_u3641_o),
    .d(mem_csr_data_add),
    .o(_al_u3642_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3643 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[42]),
    .d(ds2[42]),
    .o(\exu/alu_au/n55 [42]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3644 (
    .a(\exu/alu_au/n53 [42]),
    .b(_al_u3642_o),
    .c(\exu/alu_au/n55 [42]),
    .o(\exu/alu_data_mem_csr [42]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3645 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[41]),
    .d(ds2[41]),
    .o(\exu/alu_au/n53 [41]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3646 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[41]),
    .o(_al_u3646_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3647 (
    .a(_al_u3646_o),
    .b(mem_csr_data_xor),
    .c(ds1[41]),
    .d(ds2[41]),
    .o(_al_u3647_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3648 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[41]),
    .d(ds2[41]),
    .o(\exu/alu_au/n47 [41]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3649 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [41]),
    .c(ex_size[2]),
    .o(_al_u3649_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3650 (
    .a(_al_u3647_o),
    .b(\exu/alu_au/n47 [41]),
    .c(_al_u3649_o),
    .d(mem_csr_data_add),
    .o(_al_u3650_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3651 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[41]),
    .d(ds2[41]),
    .o(\exu/alu_au/n55 [41]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3652 (
    .a(\exu/alu_au/n53 [41]),
    .b(_al_u3650_o),
    .c(\exu/alu_au/n55 [41]),
    .o(\exu/alu_data_mem_csr [41]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3653 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[40]),
    .d(ds2[40]),
    .o(\exu/alu_au/n53 [40]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3654 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[40]),
    .o(_al_u3654_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3655 (
    .a(_al_u3654_o),
    .b(mem_csr_data_xor),
    .c(ds1[40]),
    .d(ds2[40]),
    .o(_al_u3655_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3656 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[40]),
    .d(ds2[40]),
    .o(\exu/alu_au/n47 [40]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3657 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [40]),
    .c(ex_size[2]),
    .o(_al_u3657_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3658 (
    .a(_al_u3655_o),
    .b(\exu/alu_au/n47 [40]),
    .c(_al_u3657_o),
    .d(mem_csr_data_add),
    .o(_al_u3658_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3659 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[40]),
    .d(ds2[40]),
    .o(\exu/alu_au/n55 [40]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3660 (
    .a(\exu/alu_au/n53 [40]),
    .b(_al_u3658_o),
    .c(\exu/alu_au/n55 [40]),
    .o(\exu/alu_data_mem_csr [40]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3661 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[4]),
    .d(ds2[4]),
    .o(\exu/alu_au/n53 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3662 (
    .a(\exu/alu_au/add_64 [4]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[4]),
    .o(_al_u3662_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3663 (
    .a(_al_u3662_o),
    .b(mem_csr_data_or),
    .c(ds1[4]),
    .d(ds2[4]),
    .o(_al_u3663_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3664 (
    .a(_al_u3663_o),
    .b(mem_csr_data_xor),
    .c(ds1[4]),
    .d(ds2[4]),
    .o(_al_u3664_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3665 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[4]),
    .d(ds2[4]),
    .o(\exu/alu_au/n55 [4]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3666 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[4]),
    .d(ds2[4]),
    .o(\exu/alu_au/n47 [4]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3667 (
    .a(\exu/alu_au/n53 [4]),
    .b(_al_u3664_o),
    .c(\exu/alu_au/n55 [4]),
    .d(\exu/alu_au/n47 [4]),
    .o(\exu/alu_data_mem_csr [4]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3668 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[39]),
    .d(ds2[39]),
    .o(\exu/alu_au/n53 [39]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3669 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[39]),
    .o(_al_u3669_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3670 (
    .a(_al_u3669_o),
    .b(mem_csr_data_xor),
    .c(ds1[39]),
    .d(ds2[39]),
    .o(_al_u3670_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3671 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[39]),
    .d(ds2[39]),
    .o(\exu/alu_au/n47 [39]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3672 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [39]),
    .c(ex_size[2]),
    .o(_al_u3672_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3673 (
    .a(_al_u3670_o),
    .b(\exu/alu_au/n47 [39]),
    .c(_al_u3672_o),
    .d(mem_csr_data_add),
    .o(_al_u3673_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3674 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[39]),
    .d(ds2[39]),
    .o(\exu/alu_au/n55 [39]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3675 (
    .a(\exu/alu_au/n53 [39]),
    .b(_al_u3673_o),
    .c(\exu/alu_au/n55 [39]),
    .o(\exu/alu_data_mem_csr [39]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3676 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[38]),
    .d(ds2[38]),
    .o(\exu/alu_au/n53 [38]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3677 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[38]),
    .o(_al_u3677_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3678 (
    .a(_al_u3677_o),
    .b(mem_csr_data_xor),
    .c(ds1[38]),
    .d(ds2[38]),
    .o(_al_u3678_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3679 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[38]),
    .d(ds2[38]),
    .o(\exu/alu_au/n47 [38]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3680 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [38]),
    .c(ex_size[2]),
    .o(_al_u3680_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3681 (
    .a(_al_u3678_o),
    .b(\exu/alu_au/n47 [38]),
    .c(_al_u3680_o),
    .d(mem_csr_data_add),
    .o(_al_u3681_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3682 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[38]),
    .d(ds2[38]),
    .o(\exu/alu_au/n55 [38]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3683 (
    .a(\exu/alu_au/n53 [38]),
    .b(_al_u3681_o),
    .c(\exu/alu_au/n55 [38]),
    .o(\exu/alu_data_mem_csr [38]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3684 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[37]),
    .d(ds2[37]),
    .o(\exu/alu_au/n53 [37]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3685 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[37]),
    .o(_al_u3685_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3686 (
    .a(_al_u3685_o),
    .b(mem_csr_data_xor),
    .c(ds1[37]),
    .d(ds2[37]),
    .o(_al_u3686_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3687 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[37]),
    .d(ds2[37]),
    .o(\exu/alu_au/n47 [37]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3688 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [37]),
    .c(ex_size[2]),
    .o(_al_u3688_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3689 (
    .a(_al_u3686_o),
    .b(\exu/alu_au/n47 [37]),
    .c(_al_u3688_o),
    .d(mem_csr_data_add),
    .o(_al_u3689_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3690 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[37]),
    .d(ds2[37]),
    .o(\exu/alu_au/n55 [37]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3691 (
    .a(\exu/alu_au/n53 [37]),
    .b(_al_u3689_o),
    .c(\exu/alu_au/n55 [37]),
    .o(\exu/alu_data_mem_csr [37]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3692 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[36]),
    .d(ds2[36]),
    .o(\exu/alu_au/n53 [36]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3693 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[36]),
    .o(_al_u3693_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3694 (
    .a(_al_u3693_o),
    .b(mem_csr_data_xor),
    .c(ds1[36]),
    .d(ds2[36]),
    .o(_al_u3694_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3695 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[36]),
    .d(ds2[36]),
    .o(\exu/alu_au/n47 [36]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3696 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [36]),
    .c(ex_size[2]),
    .o(_al_u3696_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3697 (
    .a(_al_u3694_o),
    .b(\exu/alu_au/n47 [36]),
    .c(_al_u3696_o),
    .d(mem_csr_data_add),
    .o(_al_u3697_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3698 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[36]),
    .d(ds2[36]),
    .o(\exu/alu_au/n55 [36]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3699 (
    .a(\exu/alu_au/n53 [36]),
    .b(_al_u3697_o),
    .c(\exu/alu_au/n55 [36]),
    .o(\exu/alu_data_mem_csr [36]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3700 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[35]),
    .d(ds2[35]),
    .o(\exu/alu_au/n53 [35]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3701 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[35]),
    .o(_al_u3701_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3702 (
    .a(_al_u3701_o),
    .b(mem_csr_data_xor),
    .c(ds1[35]),
    .d(ds2[35]),
    .o(_al_u3702_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3703 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[35]),
    .d(ds2[35]),
    .o(\exu/alu_au/n47 [35]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3704 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [35]),
    .c(ex_size[2]),
    .o(_al_u3704_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3705 (
    .a(_al_u3702_o),
    .b(\exu/alu_au/n47 [35]),
    .c(_al_u3704_o),
    .d(mem_csr_data_add),
    .o(_al_u3705_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3706 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[35]),
    .d(ds2[35]),
    .o(\exu/alu_au/n55 [35]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3707 (
    .a(\exu/alu_au/n53 [35]),
    .b(_al_u3705_o),
    .c(\exu/alu_au/n55 [35]),
    .o(\exu/alu_data_mem_csr [35]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3708 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[34]),
    .d(ds2[34]),
    .o(\exu/alu_au/n53 [34]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3709 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[34]),
    .o(_al_u3709_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3710 (
    .a(_al_u3709_o),
    .b(mem_csr_data_xor),
    .c(ds1[34]),
    .d(ds2[34]),
    .o(_al_u3710_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3711 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[34]),
    .d(ds2[34]),
    .o(\exu/alu_au/n47 [34]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3712 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [34]),
    .c(ex_size[2]),
    .o(_al_u3712_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3713 (
    .a(_al_u3710_o),
    .b(\exu/alu_au/n47 [34]),
    .c(_al_u3712_o),
    .d(mem_csr_data_add),
    .o(_al_u3713_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3714 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[34]),
    .d(ds2[34]),
    .o(\exu/alu_au/n55 [34]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3715 (
    .a(\exu/alu_au/n53 [34]),
    .b(_al_u3713_o),
    .c(\exu/alu_au/n55 [34]),
    .o(\exu/alu_data_mem_csr [34]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3716 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[33]),
    .d(ds2[33]),
    .o(\exu/alu_au/n53 [33]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3717 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[33]),
    .o(_al_u3717_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3718 (
    .a(_al_u3717_o),
    .b(mem_csr_data_xor),
    .c(ds1[33]),
    .d(ds2[33]),
    .o(_al_u3718_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3719 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[33]),
    .d(ds2[33]),
    .o(\exu/alu_au/n47 [33]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3720 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [33]),
    .c(ex_size[2]),
    .o(_al_u3720_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3721 (
    .a(_al_u3718_o),
    .b(\exu/alu_au/n47 [33]),
    .c(_al_u3720_o),
    .d(mem_csr_data_add),
    .o(_al_u3721_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3722 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[33]),
    .d(ds2[33]),
    .o(\exu/alu_au/n55 [33]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3723 (
    .a(\exu/alu_au/n53 [33]),
    .b(_al_u3721_o),
    .c(\exu/alu_au/n55 [33]),
    .o(\exu/alu_data_mem_csr [33]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3724 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[32]),
    .d(ds2[32]),
    .o(\exu/alu_au/n53 [32]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u3725 (
    .a(mem_csr_data_ds2),
    .b(mem_csr_data_or),
    .c(ds2[32]),
    .o(_al_u3725_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u3726 (
    .a(_al_u3725_o),
    .b(mem_csr_data_xor),
    .c(ds1[32]),
    .d(ds2[32]),
    .o(_al_u3726_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3727 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[32]),
    .d(ds2[32]),
    .o(\exu/alu_au/n47 [32]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u3728 (
    .a(\exu/alu_au/add_64 [31]),
    .b(\exu/alu_au/add_64 [32]),
    .c(ex_size[2]),
    .o(_al_u3728_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*~C))"),
    .INIT(16'h1011))
    _al_u3729 (
    .a(_al_u3726_o),
    .b(\exu/alu_au/n47 [32]),
    .c(_al_u3728_o),
    .d(mem_csr_data_add),
    .o(_al_u3729_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3730 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[32]),
    .d(ds2[32]),
    .o(\exu/alu_au/n55 [32]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u3731 (
    .a(\exu/alu_au/n53 [32]),
    .b(_al_u3729_o),
    .c(\exu/alu_au/n55 [32]),
    .o(\exu/alu_data_mem_csr [32]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3732 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[31]),
    .d(ds2[31]),
    .o(\exu/alu_au/n53 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3733 (
    .a(\exu/alu_au/add_64 [31]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[31]),
    .o(_al_u3733_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3734 (
    .a(_al_u3733_o),
    .b(mem_csr_data_or),
    .c(ds1[31]),
    .d(ds2[31]),
    .o(_al_u3734_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3735 (
    .a(_al_u3734_o),
    .b(mem_csr_data_xor),
    .c(ds1[31]),
    .d(ds2[31]),
    .o(_al_u3735_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3736 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[31]),
    .d(ds2[31]),
    .o(\exu/alu_au/n55 [31]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3737 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[31]),
    .d(ds2[31]),
    .o(\exu/alu_au/n47 [31]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3738 (
    .a(\exu/alu_au/n53 [31]),
    .b(_al_u3735_o),
    .c(\exu/alu_au/n55 [31]),
    .d(\exu/alu_au/n47 [31]),
    .o(\exu/alu_data_mem_csr [31]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3739 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[30]),
    .d(ds2[30]),
    .o(\exu/alu_au/n53 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3740 (
    .a(\exu/alu_au/add_64 [30]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[30]),
    .o(_al_u3740_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3741 (
    .a(_al_u3740_o),
    .b(mem_csr_data_or),
    .c(ds1[30]),
    .d(ds2[30]),
    .o(_al_u3741_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3742 (
    .a(_al_u3741_o),
    .b(mem_csr_data_xor),
    .c(ds1[30]),
    .d(ds2[30]),
    .o(_al_u3742_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3743 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[30]),
    .d(ds2[30]),
    .o(\exu/alu_au/n55 [30]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3744 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[30]),
    .d(ds2[30]),
    .o(\exu/alu_au/n47 [30]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3745 (
    .a(\exu/alu_au/n53 [30]),
    .b(_al_u3742_o),
    .c(\exu/alu_au/n55 [30]),
    .d(\exu/alu_au/n47 [30]),
    .o(\exu/alu_data_mem_csr [30]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3746 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[3]),
    .d(ds2[3]),
    .o(\exu/alu_au/n53 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3747 (
    .a(\exu/alu_au/add_64 [3]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[3]),
    .o(_al_u3747_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3748 (
    .a(_al_u3747_o),
    .b(mem_csr_data_or),
    .c(ds1[3]),
    .d(ds2[3]),
    .o(_al_u3748_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3749 (
    .a(_al_u3748_o),
    .b(mem_csr_data_xor),
    .c(ds1[3]),
    .d(ds2[3]),
    .o(_al_u3749_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3750 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[3]),
    .d(ds2[3]),
    .o(\exu/alu_au/n55 [3]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3751 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[3]),
    .d(ds2[3]),
    .o(\exu/alu_au/n47 [3]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3752 (
    .a(\exu/alu_au/n53 [3]),
    .b(_al_u3749_o),
    .c(\exu/alu_au/n55 [3]),
    .d(\exu/alu_au/n47 [3]),
    .o(\exu/alu_data_mem_csr [3]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3753 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[29]),
    .d(ds2[29]),
    .o(\exu/alu_au/n53 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3754 (
    .a(\exu/alu_au/add_64 [29]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[29]),
    .o(_al_u3754_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3755 (
    .a(_al_u3754_o),
    .b(mem_csr_data_or),
    .c(ds1[29]),
    .d(ds2[29]),
    .o(_al_u3755_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3756 (
    .a(_al_u3755_o),
    .b(mem_csr_data_xor),
    .c(ds1[29]),
    .d(ds2[29]),
    .o(_al_u3756_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3757 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[29]),
    .d(ds2[29]),
    .o(\exu/alu_au/n55 [29]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3758 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[29]),
    .d(ds2[29]),
    .o(\exu/alu_au/n47 [29]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3759 (
    .a(\exu/alu_au/n53 [29]),
    .b(_al_u3756_o),
    .c(\exu/alu_au/n55 [29]),
    .d(\exu/alu_au/n47 [29]),
    .o(\exu/alu_data_mem_csr [29]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3760 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[28]),
    .d(ds2[28]),
    .o(\exu/alu_au/n53 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3761 (
    .a(\exu/alu_au/add_64 [28]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[28]),
    .o(_al_u3761_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3762 (
    .a(_al_u3761_o),
    .b(mem_csr_data_or),
    .c(ds1[28]),
    .d(ds2[28]),
    .o(_al_u3762_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3763 (
    .a(_al_u3762_o),
    .b(mem_csr_data_xor),
    .c(ds1[28]),
    .d(ds2[28]),
    .o(_al_u3763_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3764 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[28]),
    .d(ds2[28]),
    .o(\exu/alu_au/n55 [28]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3765 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[28]),
    .d(ds2[28]),
    .o(\exu/alu_au/n47 [28]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3766 (
    .a(\exu/alu_au/n53 [28]),
    .b(_al_u3763_o),
    .c(\exu/alu_au/n55 [28]),
    .d(\exu/alu_au/n47 [28]),
    .o(\exu/alu_data_mem_csr [28]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3767 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[27]),
    .d(ds2[27]),
    .o(\exu/alu_au/n53 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3768 (
    .a(\exu/alu_au/add_64 [27]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[27]),
    .o(_al_u3768_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3769 (
    .a(_al_u3768_o),
    .b(mem_csr_data_or),
    .c(ds1[27]),
    .d(ds2[27]),
    .o(_al_u3769_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3770 (
    .a(_al_u3769_o),
    .b(mem_csr_data_xor),
    .c(ds1[27]),
    .d(ds2[27]),
    .o(_al_u3770_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3771 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[27]),
    .d(ds2[27]),
    .o(\exu/alu_au/n55 [27]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3772 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[27]),
    .d(ds2[27]),
    .o(\exu/alu_au/n47 [27]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3773 (
    .a(\exu/alu_au/n53 [27]),
    .b(_al_u3770_o),
    .c(\exu/alu_au/n55 [27]),
    .d(\exu/alu_au/n47 [27]),
    .o(\exu/alu_data_mem_csr [27]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3774 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[26]),
    .d(ds2[26]),
    .o(\exu/alu_au/n53 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3775 (
    .a(\exu/alu_au/add_64 [26]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[26]),
    .o(_al_u3775_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3776 (
    .a(_al_u3775_o),
    .b(mem_csr_data_or),
    .c(ds1[26]),
    .d(ds2[26]),
    .o(_al_u3776_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3777 (
    .a(_al_u3776_o),
    .b(mem_csr_data_xor),
    .c(ds1[26]),
    .d(ds2[26]),
    .o(_al_u3777_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3778 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[26]),
    .d(ds2[26]),
    .o(\exu/alu_au/n55 [26]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3779 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[26]),
    .d(ds2[26]),
    .o(\exu/alu_au/n47 [26]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3780 (
    .a(\exu/alu_au/n53 [26]),
    .b(_al_u3777_o),
    .c(\exu/alu_au/n55 [26]),
    .d(\exu/alu_au/n47 [26]),
    .o(\exu/alu_data_mem_csr [26]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3781 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[25]),
    .d(ds2[25]),
    .o(\exu/alu_au/n53 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3782 (
    .a(\exu/alu_au/add_64 [25]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[25]),
    .o(_al_u3782_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3783 (
    .a(_al_u3782_o),
    .b(mem_csr_data_or),
    .c(ds1[25]),
    .d(ds2[25]),
    .o(_al_u3783_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3784 (
    .a(_al_u3783_o),
    .b(mem_csr_data_xor),
    .c(ds1[25]),
    .d(ds2[25]),
    .o(_al_u3784_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3785 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[25]),
    .d(ds2[25]),
    .o(\exu/alu_au/n55 [25]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3786 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[25]),
    .d(ds2[25]),
    .o(\exu/alu_au/n47 [25]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3787 (
    .a(\exu/alu_au/n53 [25]),
    .b(_al_u3784_o),
    .c(\exu/alu_au/n55 [25]),
    .d(\exu/alu_au/n47 [25]),
    .o(\exu/alu_data_mem_csr [25]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3788 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[24]),
    .d(ds2[24]),
    .o(\exu/alu_au/n53 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3789 (
    .a(\exu/alu_au/add_64 [24]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[24]),
    .o(_al_u3789_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3790 (
    .a(_al_u3789_o),
    .b(mem_csr_data_or),
    .c(ds1[24]),
    .d(ds2[24]),
    .o(_al_u3790_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3791 (
    .a(_al_u3790_o),
    .b(mem_csr_data_xor),
    .c(ds1[24]),
    .d(ds2[24]),
    .o(_al_u3791_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3792 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[24]),
    .d(ds2[24]),
    .o(\exu/alu_au/n55 [24]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3793 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[24]),
    .d(ds2[24]),
    .o(\exu/alu_au/n47 [24]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3794 (
    .a(\exu/alu_au/n53 [24]),
    .b(_al_u3791_o),
    .c(\exu/alu_au/n55 [24]),
    .d(\exu/alu_au/n47 [24]),
    .o(\exu/alu_data_mem_csr [24]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3795 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[23]),
    .d(ds2[23]),
    .o(\exu/alu_au/n53 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3796 (
    .a(\exu/alu_au/add_64 [23]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[23]),
    .o(_al_u3796_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3797 (
    .a(_al_u3796_o),
    .b(mem_csr_data_or),
    .c(ds1[23]),
    .d(ds2[23]),
    .o(_al_u3797_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3798 (
    .a(_al_u3797_o),
    .b(mem_csr_data_xor),
    .c(ds1[23]),
    .d(ds2[23]),
    .o(_al_u3798_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3799 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[23]),
    .d(ds2[23]),
    .o(\exu/alu_au/n55 [23]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3800 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[23]),
    .d(ds2[23]),
    .o(\exu/alu_au/n47 [23]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3801 (
    .a(\exu/alu_au/n53 [23]),
    .b(_al_u3798_o),
    .c(\exu/alu_au/n55 [23]),
    .d(\exu/alu_au/n47 [23]),
    .o(\exu/alu_data_mem_csr [23]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3802 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[22]),
    .d(ds2[22]),
    .o(\exu/alu_au/n53 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3803 (
    .a(\exu/alu_au/add_64 [22]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[22]),
    .o(_al_u3803_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3804 (
    .a(_al_u3803_o),
    .b(mem_csr_data_or),
    .c(ds1[22]),
    .d(ds2[22]),
    .o(_al_u3804_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3805 (
    .a(_al_u3804_o),
    .b(mem_csr_data_xor),
    .c(ds1[22]),
    .d(ds2[22]),
    .o(_al_u3805_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3806 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[22]),
    .d(ds2[22]),
    .o(\exu/alu_au/n55 [22]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3807 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[22]),
    .d(ds2[22]),
    .o(\exu/alu_au/n47 [22]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3808 (
    .a(\exu/alu_au/n53 [22]),
    .b(_al_u3805_o),
    .c(\exu/alu_au/n55 [22]),
    .d(\exu/alu_au/n47 [22]),
    .o(\exu/alu_data_mem_csr [22]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3809 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[21]),
    .d(ds2[21]),
    .o(\exu/alu_au/n53 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3810 (
    .a(\exu/alu_au/add_64 [21]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[21]),
    .o(_al_u3810_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3811 (
    .a(_al_u3810_o),
    .b(mem_csr_data_or),
    .c(ds1[21]),
    .d(ds2[21]),
    .o(_al_u3811_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3812 (
    .a(_al_u3811_o),
    .b(mem_csr_data_xor),
    .c(ds1[21]),
    .d(ds2[21]),
    .o(_al_u3812_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3813 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[21]),
    .d(ds2[21]),
    .o(\exu/alu_au/n55 [21]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3814 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[21]),
    .d(ds2[21]),
    .o(\exu/alu_au/n47 [21]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3815 (
    .a(\exu/alu_au/n53 [21]),
    .b(_al_u3812_o),
    .c(\exu/alu_au/n55 [21]),
    .d(\exu/alu_au/n47 [21]),
    .o(\exu/alu_data_mem_csr [21]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3816 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[20]),
    .d(ds2[20]),
    .o(\exu/alu_au/n53 [20]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3817 (
    .a(\exu/alu_au/add_64 [20]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[20]),
    .o(_al_u3817_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3818 (
    .a(_al_u3817_o),
    .b(mem_csr_data_or),
    .c(ds1[20]),
    .d(ds2[20]),
    .o(_al_u3818_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3819 (
    .a(_al_u3818_o),
    .b(mem_csr_data_xor),
    .c(ds1[20]),
    .d(ds2[20]),
    .o(_al_u3819_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3820 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[20]),
    .d(ds2[20]),
    .o(\exu/alu_au/n55 [20]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3821 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[20]),
    .d(ds2[20]),
    .o(\exu/alu_au/n47 [20]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3822 (
    .a(\exu/alu_au/n53 [20]),
    .b(_al_u3819_o),
    .c(\exu/alu_au/n55 [20]),
    .d(\exu/alu_au/n47 [20]),
    .o(\exu/alu_data_mem_csr [20]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3823 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[2]),
    .d(ds2[2]),
    .o(\exu/alu_au/n53 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3824 (
    .a(\exu/alu_au/add_64 [2]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[2]),
    .o(_al_u3824_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3825 (
    .a(_al_u3824_o),
    .b(mem_csr_data_or),
    .c(ds1[2]),
    .d(ds2[2]),
    .o(_al_u3825_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3826 (
    .a(_al_u3825_o),
    .b(mem_csr_data_xor),
    .c(ds1[2]),
    .d(ds2[2]),
    .o(_al_u3826_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3827 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[2]),
    .d(ds2[2]),
    .o(\exu/alu_au/n55 [2]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3828 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[2]),
    .d(ds2[2]),
    .o(\exu/alu_au/n47 [2]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3829 (
    .a(\exu/alu_au/n53 [2]),
    .b(_al_u3826_o),
    .c(\exu/alu_au/n55 [2]),
    .d(\exu/alu_au/n47 [2]),
    .o(\exu/alu_data_mem_csr [2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3830 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[19]),
    .d(ds2[19]),
    .o(\exu/alu_au/n53 [19]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3831 (
    .a(\exu/alu_au/add_64 [19]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[19]),
    .o(_al_u3831_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3832 (
    .a(_al_u3831_o),
    .b(mem_csr_data_or),
    .c(ds1[19]),
    .d(ds2[19]),
    .o(_al_u3832_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3833 (
    .a(_al_u3832_o),
    .b(mem_csr_data_xor),
    .c(ds1[19]),
    .d(ds2[19]),
    .o(_al_u3833_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3834 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[19]),
    .d(ds2[19]),
    .o(\exu/alu_au/n55 [19]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3835 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[19]),
    .d(ds2[19]),
    .o(\exu/alu_au/n47 [19]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3836 (
    .a(\exu/alu_au/n53 [19]),
    .b(_al_u3833_o),
    .c(\exu/alu_au/n55 [19]),
    .d(\exu/alu_au/n47 [19]),
    .o(\exu/alu_data_mem_csr [19]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3837 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[18]),
    .d(ds2[18]),
    .o(\exu/alu_au/n53 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3838 (
    .a(\exu/alu_au/add_64 [18]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[18]),
    .o(_al_u3838_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3839 (
    .a(_al_u3838_o),
    .b(mem_csr_data_or),
    .c(ds1[18]),
    .d(ds2[18]),
    .o(_al_u3839_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3840 (
    .a(_al_u3839_o),
    .b(mem_csr_data_xor),
    .c(ds1[18]),
    .d(ds2[18]),
    .o(_al_u3840_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3841 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[18]),
    .d(ds2[18]),
    .o(\exu/alu_au/n55 [18]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3842 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[18]),
    .d(ds2[18]),
    .o(\exu/alu_au/n47 [18]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3843 (
    .a(\exu/alu_au/n53 [18]),
    .b(_al_u3840_o),
    .c(\exu/alu_au/n55 [18]),
    .d(\exu/alu_au/n47 [18]),
    .o(\exu/alu_data_mem_csr [18]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3844 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[17]),
    .d(ds2[17]),
    .o(\exu/alu_au/n53 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3845 (
    .a(\exu/alu_au/add_64 [17]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[17]),
    .o(_al_u3845_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3846 (
    .a(_al_u3845_o),
    .b(mem_csr_data_or),
    .c(ds1[17]),
    .d(ds2[17]),
    .o(_al_u3846_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3847 (
    .a(_al_u3846_o),
    .b(mem_csr_data_xor),
    .c(ds1[17]),
    .d(ds2[17]),
    .o(_al_u3847_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3848 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[17]),
    .d(ds2[17]),
    .o(\exu/alu_au/n55 [17]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3849 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[17]),
    .d(ds2[17]),
    .o(\exu/alu_au/n47 [17]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3850 (
    .a(\exu/alu_au/n53 [17]),
    .b(_al_u3847_o),
    .c(\exu/alu_au/n55 [17]),
    .d(\exu/alu_au/n47 [17]),
    .o(\exu/alu_data_mem_csr [17]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3851 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[16]),
    .d(ds2[16]),
    .o(\exu/alu_au/n53 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3852 (
    .a(\exu/alu_au/add_64 [16]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[16]),
    .o(_al_u3852_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3853 (
    .a(_al_u3852_o),
    .b(mem_csr_data_or),
    .c(ds1[16]),
    .d(ds2[16]),
    .o(_al_u3853_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3854 (
    .a(_al_u3853_o),
    .b(mem_csr_data_xor),
    .c(ds1[16]),
    .d(ds2[16]),
    .o(_al_u3854_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3855 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[16]),
    .d(ds2[16]),
    .o(\exu/alu_au/n55 [16]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3856 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[16]),
    .d(ds2[16]),
    .o(\exu/alu_au/n47 [16]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3857 (
    .a(\exu/alu_au/n53 [16]),
    .b(_al_u3854_o),
    .c(\exu/alu_au/n55 [16]),
    .d(\exu/alu_au/n47 [16]),
    .o(\exu/alu_data_mem_csr [16]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3858 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[15]),
    .d(ds2[15]),
    .o(\exu/alu_au/n53 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3859 (
    .a(\exu/alu_au/add_64 [15]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[15]),
    .o(_al_u3859_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3860 (
    .a(_al_u3859_o),
    .b(mem_csr_data_or),
    .c(ds1[15]),
    .d(ds2[15]),
    .o(_al_u3860_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3861 (
    .a(_al_u3860_o),
    .b(mem_csr_data_xor),
    .c(ds1[15]),
    .d(ds2[15]),
    .o(_al_u3861_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3862 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[15]),
    .d(ds2[15]),
    .o(\exu/alu_au/n55 [15]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3863 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[15]),
    .d(ds2[15]),
    .o(\exu/alu_au/n47 [15]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3864 (
    .a(\exu/alu_au/n53 [15]),
    .b(_al_u3861_o),
    .c(\exu/alu_au/n55 [15]),
    .d(\exu/alu_au/n47 [15]),
    .o(\exu/alu_data_mem_csr [15]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3865 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[14]),
    .d(ds2[14]),
    .o(\exu/alu_au/n53 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3866 (
    .a(\exu/alu_au/add_64 [14]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[14]),
    .o(_al_u3866_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3867 (
    .a(_al_u3866_o),
    .b(mem_csr_data_or),
    .c(ds1[14]),
    .d(ds2[14]),
    .o(_al_u3867_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3868 (
    .a(_al_u3867_o),
    .b(mem_csr_data_xor),
    .c(ds1[14]),
    .d(ds2[14]),
    .o(_al_u3868_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3869 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[14]),
    .d(ds2[14]),
    .o(\exu/alu_au/n55 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    _al_u3870 (
    .a(and_clr),
    .b(ds1[14]),
    .c(ds2[14]),
    .o(\exu/alu_au/alu_and [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3871 (
    .a(\exu/alu_au/alu_and [14]),
    .b(mem_csr_data_and),
    .o(\exu/alu_au/n47 [14]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3872 (
    .a(\exu/alu_au/n53 [14]),
    .b(_al_u3868_o),
    .c(\exu/alu_au/n55 [14]),
    .d(\exu/alu_au/n47 [14]),
    .o(\exu/alu_data_mem_csr [14]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3873 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[13]),
    .d(ds2[13]),
    .o(\exu/alu_au/n53 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3874 (
    .a(\exu/alu_au/add_64 [13]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[13]),
    .o(_al_u3874_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3875 (
    .a(_al_u3874_o),
    .b(mem_csr_data_or),
    .c(ds1[13]),
    .d(ds2[13]),
    .o(_al_u3875_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3876 (
    .a(_al_u3875_o),
    .b(mem_csr_data_xor),
    .c(ds1[13]),
    .d(ds2[13]),
    .o(_al_u3876_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3877 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[13]),
    .d(ds2[13]),
    .o(\exu/alu_au/n55 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    _al_u3878 (
    .a(and_clr),
    .b(ds1[13]),
    .c(ds2[13]),
    .o(\exu/alu_au/alu_and [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3879 (
    .a(\exu/alu_au/alu_and [13]),
    .b(mem_csr_data_and),
    .o(\exu/alu_au/n47 [13]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3880 (
    .a(\exu/alu_au/n53 [13]),
    .b(_al_u3876_o),
    .c(\exu/alu_au/n55 [13]),
    .d(\exu/alu_au/n47 [13]),
    .o(\exu/alu_data_mem_csr [13]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3881 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[12]),
    .d(ds2[12]),
    .o(\exu/alu_au/n53 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3882 (
    .a(\exu/alu_au/add_64 [12]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[12]),
    .o(_al_u3882_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3883 (
    .a(_al_u3882_o),
    .b(mem_csr_data_or),
    .c(ds1[12]),
    .d(ds2[12]),
    .o(_al_u3883_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3884 (
    .a(_al_u3883_o),
    .b(mem_csr_data_xor),
    .c(ds1[12]),
    .d(ds2[12]),
    .o(_al_u3884_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3885 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[12]),
    .d(ds2[12]),
    .o(\exu/alu_au/n55 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    _al_u3886 (
    .a(and_clr),
    .b(ds1[12]),
    .c(ds2[12]),
    .o(\exu/alu_au/alu_and [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3887 (
    .a(\exu/alu_au/alu_and [12]),
    .b(mem_csr_data_and),
    .o(\exu/alu_au/n47 [12]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3888 (
    .a(\exu/alu_au/n53 [12]),
    .b(_al_u3884_o),
    .c(\exu/alu_au/n55 [12]),
    .d(\exu/alu_au/n47 [12]),
    .o(\exu/alu_data_mem_csr [12]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3889 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[11]),
    .d(ds2[11]),
    .o(\exu/alu_au/n53 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3890 (
    .a(\exu/alu_au/add_64 [11]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[11]),
    .o(_al_u3890_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3891 (
    .a(_al_u3890_o),
    .b(mem_csr_data_or),
    .c(ds1[11]),
    .d(ds2[11]),
    .o(_al_u3891_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3892 (
    .a(_al_u3891_o),
    .b(mem_csr_data_xor),
    .c(ds1[11]),
    .d(ds2[11]),
    .o(_al_u3892_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3893 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[11]),
    .d(ds2[11]),
    .o(\exu/alu_au/n55 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    _al_u3894 (
    .a(and_clr),
    .b(ds1[11]),
    .c(ds2[11]),
    .o(\exu/alu_au/alu_and [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3895 (
    .a(\exu/alu_au/alu_and [11]),
    .b(mem_csr_data_and),
    .o(\exu/alu_au/n47 [11]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3896 (
    .a(\exu/alu_au/n53 [11]),
    .b(_al_u3892_o),
    .c(\exu/alu_au/n55 [11]),
    .d(\exu/alu_au/n47 [11]),
    .o(\exu/alu_data_mem_csr [11]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3897 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[10]),
    .d(ds2[10]),
    .o(\exu/alu_au/n53 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3898 (
    .a(\exu/alu_au/add_64 [10]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[10]),
    .o(_al_u3898_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3899 (
    .a(_al_u3898_o),
    .b(mem_csr_data_or),
    .c(ds1[10]),
    .d(ds2[10]),
    .o(_al_u3899_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3900 (
    .a(_al_u3899_o),
    .b(mem_csr_data_xor),
    .c(ds1[10]),
    .d(ds2[10]),
    .o(_al_u3900_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3901 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[10]),
    .d(ds2[10]),
    .o(\exu/alu_au/n55 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    _al_u3902 (
    .a(and_clr),
    .b(ds1[10]),
    .c(ds2[10]),
    .o(\exu/alu_au/alu_and [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3903 (
    .a(\exu/alu_au/alu_and [10]),
    .b(mem_csr_data_and),
    .o(\exu/alu_au/n47 [10]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3904 (
    .a(\exu/alu_au/n53 [10]),
    .b(_al_u3900_o),
    .c(\exu/alu_au/n55 [10]),
    .d(\exu/alu_au/n47 [10]),
    .o(\exu/alu_data_mem_csr [10]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3905 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[1]),
    .d(ds2[1]),
    .o(\exu/alu_au/n53 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3906 (
    .a(\exu/alu_au/add_64 [1]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[1]),
    .o(_al_u3906_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3907 (
    .a(_al_u3906_o),
    .b(mem_csr_data_or),
    .c(ds1[1]),
    .d(ds2[1]),
    .o(_al_u3907_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3908 (
    .a(_al_u3907_o),
    .b(mem_csr_data_xor),
    .c(ds1[1]),
    .d(ds2[1]),
    .o(_al_u3908_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3909 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[1]),
    .d(ds2[1]),
    .o(\exu/alu_au/n55 [1]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3910 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[1]),
    .d(ds2[1]),
    .o(\exu/alu_au/n47 [1]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3911 (
    .a(\exu/alu_au/n53 [1]),
    .b(_al_u3908_o),
    .c(\exu/alu_au/n55 [1]),
    .d(\exu/alu_au/n47 [1]),
    .o(\exu/alu_data_mem_csr [1]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u3912 (
    .a(_al_u3430_o),
    .b(mem_csr_data_max),
    .c(ds1[0]),
    .d(ds2[0]),
    .o(\exu/alu_au/n53 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u3913 (
    .a(\exu/alu_au/add_64 [0]),
    .b(mem_csr_data_add),
    .c(mem_csr_data_ds2),
    .d(ds2[0]),
    .o(_al_u3913_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u3914 (
    .a(_al_u3913_o),
    .b(mem_csr_data_or),
    .c(ds1[0]),
    .d(ds2[0]),
    .o(_al_u3914_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u3915 (
    .a(_al_u3914_o),
    .b(mem_csr_data_xor),
    .c(ds1[0]),
    .d(ds2[0]),
    .o(_al_u3915_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u3916 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(mem_csr_data_min),
    .c(ds1[0]),
    .d(ds2[0]),
    .o(\exu/alu_au/n55 [0]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u3917 (
    .a(and_clr),
    .b(mem_csr_data_and),
    .c(ds1[0]),
    .d(ds2[0]),
    .o(\exu/alu_au/n47 [0]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*~A)"),
    .INIT(16'hfffb))
    _al_u3918 (
    .a(\exu/alu_au/n53 [0]),
    .b(_al_u3915_o),
    .c(\exu/alu_au/n55 [0]),
    .d(\exu/alu_au/n47 [0]),
    .o(\exu/alu_data_mem_csr [0]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u3919 (
    .a(\ins_dec/op_store ),
    .b(\ins_dec/op_load ),
    .c(_al_u3216_o),
    .o(_al_u3919_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3920 (
    .a(_al_u3919_o),
    .b(_al_u3217_o),
    .c(_al_u3384_o),
    .o(\ins_dec/dbyte ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3921 (
    .a(_al_u3919_o),
    .b(_al_u3217_o),
    .c(_al_u3384_o),
    .o(\ins_dec/sbyte ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u3922 (
    .a(\ins_dec/funct6_0_lutinv ),
    .b(id_ins[25]),
    .o(\ins_dec/funct7_0_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*~C))"),
    .INIT(16'h1110))
    _al_u3923 (
    .a(_al_u2929_o),
    .b(_al_u2930_o),
    .c(_al_u2931_o),
    .d(_al_u2932_o),
    .o(_al_u3923_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3924 (
    .a(_al_u2929_o),
    .b(_al_u2930_o),
    .o(_al_u3924_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3925 (
    .a(_al_u3924_o),
    .b(_al_u2938_o),
    .c(_al_u2939_o),
    .d(_al_u2944_o),
    .o(_al_u3925_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3926 (
    .a(\ins_dec/funct7_0_lutinv ),
    .b(_al_u3923_o),
    .c(_al_u3925_o),
    .o(_al_u3926_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u3927 (
    .a(_al_u3924_o),
    .b(_al_u2938_o),
    .c(_al_u2939_o),
    .d(_al_u2946_o),
    .o(_al_u3927_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3928 (
    .a(_al_u2931_o),
    .b(_al_u2932_o),
    .o(_al_u3928_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u3929 (
    .a(_al_u3926_o),
    .b(_al_u3927_o),
    .c(_al_u3928_o),
    .o(_al_u3929_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u3930 (
    .a(_al_u3929_o),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .d(_al_u3384_o),
    .o(\ins_dec/n135 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u3931 (
    .a(_al_u3929_o),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .d(_al_u3384_o),
    .o(\ins_dec/n136 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u3932 (
    .a(id_ins[31]),
    .b(id_ins[30]),
    .c(id_ins[28]),
    .d(id_ins[26]),
    .o(_al_u3932_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3933 (
    .a(_al_u3932_o),
    .b(id_ins[29]),
    .c(id_ins[27]),
    .d(id_ins[25]),
    .o(\ins_dec/funct7_32_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3934 (
    .a(\ins_dec/funct3_0_lutinv ),
    .b(\ins_dec/funct7_32_lutinv ),
    .c(_al_u3925_o),
    .o(\ins_dec/n133 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u3935 (
    .a(_al_u3929_o),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .d(_al_u3384_o),
    .o(\ins_dec/n134 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3936 (
    .a(_al_u3925_o),
    .b(_al_u3928_o),
    .o(\ins_dec/op_32_reg_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3937 (
    .a(\ins_dec/funct7_0_lutinv ),
    .b(\ins_dec/funct3_0_lutinv ),
    .c(\ins_dec/op_32_reg_lutinv ),
    .o(\ins_dec/ins_addw ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3938 (
    .a(\ins_dec/op_amo ),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .o(_al_u3938_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3939 (
    .a(_al_u3938_o),
    .b(id_ins[28]),
    .c(id_ins[27]),
    .o(_al_u3939_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*C*B))"),
    .INIT(16'heaaa))
    _al_u3940 (
    .a(\ins_dec/ins_addw ),
    .b(_al_u3939_o),
    .c(_al_u3399_o),
    .d(_al_u3384_o),
    .o(\ins_dec/n146 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3941 (
    .a(_al_u3939_o),
    .b(id_ins[29]),
    .c(_al_u3388_o),
    .o(\ins_dec/n152 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3942 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u2914_o),
    .o(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3943 (
    .a(_al_u2705_o),
    .b(hrdata_pad[7]),
    .o(uncache_data[7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3944 (
    .a(\biu/cache_ctrl_logic/statu [2]),
    .b(\biu/cache_ctrl_logic/statu [3]),
    .c(\biu/cache_ctrl_logic/statu [4]),
    .o(_al_u3944_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3945 (
    .a(_al_u3209_o),
    .b(_al_u3944_o),
    .o(_al_u3945_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A)"),
    .INIT(16'hddd8))
    _al_u3946 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(uncache_data[7]),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [7]),
    .o(\biu/cache_ctrl_logic/n165 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3947 (
    .a(_al_u2837_o),
    .b(_al_u3944_o),
    .o(_al_u3947_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(D)*~(A)+~(~C*~B)*D*~(A)+~(~(~C*~B))*D*A+~(~C*~B)*D*A)"),
    .INIT(16'hfe54))
    _al_u3948 (
    .a(\biu/cache_ctrl_logic/n149 ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [7]),
    .d(\biu/cache_ctrl_logic/pte_temp [7]),
    .o(\biu/cache_ctrl_logic/n158 [7]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u3949 (
    .a(\biu/cache_ctrl_logic/n149 ),
    .b(\biu/cache_ctrl_logic/l1d_value ),
    .o(\biu/cache_ctrl_logic/l1d_value_d ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3950 (
    .a(_al_u3944_o),
    .b(\biu/cache_ctrl_logic/statu [0]),
    .c(\biu/cache_ctrl_logic/statu [1]),
    .o(_al_u3950_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(D)*~(A)+~(~C*~B)*D*~(A)+~(~(~C*~B))*D*A+~(~C*~B)*D*A)"),
    .INIT(16'hfe54))
    _al_u3951 (
    .a(\biu/cache_ctrl_logic/n135 ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [7]),
    .d(\biu/cache_ctrl_logic/pte_temp [7]),
    .o(\biu/cache_ctrl_logic/n147 [7]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u3952 (
    .a(\biu/cache_ctrl_logic/n135 ),
    .b(\biu/cache_ctrl_logic/l1i_value ),
    .o(\biu/cache_ctrl_logic/l1i_value_d ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3953 (
    .a(_al_u3929_o),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .o(\ins_dec/n139 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3954 (
    .a(_al_u2938_o),
    .b(_al_u2939_o),
    .c(_al_u2944_o),
    .d(_al_u3923_o),
    .o(\ins_dec/op_lui_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u3955 (
    .a(_al_u2938_o),
    .b(_al_u2939_o),
    .c(_al_u2946_o),
    .d(_al_u3923_o),
    .o(_al_u3955_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u3956 (
    .a(_al_u3213_o),
    .b(_al_u3214_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(_al_u3955_o),
    .o(_al_u3956_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u3957 (
    .a(\ins_fetch/ins_shift [19]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [19]),
    .o(id_ins[19]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3958 (
    .a(_al_u3956_o),
    .b(id_ins[19]),
    .o(id_rs1_index[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u3959 (
    .a(\ins_fetch/ins_shift [18]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [18]),
    .o(id_ins[18]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3960 (
    .a(_al_u3956_o),
    .b(id_ins[18]),
    .o(id_rs1_index[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u3961 (
    .a(\ins_fetch/ins_shift [17]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [17]),
    .o(id_ins[17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3962 (
    .a(_al_u3956_o),
    .b(id_ins[17]),
    .o(id_rs1_index[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u3963 (
    .a(\ins_fetch/ins_shift [16]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [16]),
    .o(id_ins[16]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3964 (
    .a(_al_u3956_o),
    .b(id_ins[16]),
    .o(id_rs1_index[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u3965 (
    .a(\ins_fetch/ins_shift [15]),
    .b(\ins_fetch/hold ),
    .c(\ins_fetch/ins_hold [15]),
    .o(id_ins[15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3966 (
    .a(_al_u3956_o),
    .b(id_ins[15]),
    .o(id_rs1_index[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3967 (
    .a(\ins_dec/op_store ),
    .b(\ins_dec/op_load ),
    .o(\ins_dec/mux24_b10_sel_is_0_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u3968 (
    .a(\ins_dec/n302 ),
    .b(\ins_dec/mux24_b10_sel_is_0_o ),
    .c(id_ins[31]),
    .o(\ins_dec/n291 [20]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u3969 (
    .a(_al_u3939_o),
    .b(id_ins[31]),
    .c(id_ins[30]),
    .d(id_ins[29]),
    .o(_al_u3969_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u3970 (
    .a(_al_u3969_o),
    .b(\ins_dec/n71 ),
    .o(\ins_dec/n148 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u3971 (
    .a(id_system),
    .b(_al_u3217_o),
    .c(_al_u3384_o),
    .o(\ins_dec/n149_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u3972 (
    .a(id_ins[31]),
    .b(id_ins[30]),
    .c(id_ins[29]),
    .o(_al_u3972_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u3973 (
    .a(_al_u3972_o),
    .b(id_ins[28]),
    .c(id_ins[27]),
    .o(\ins_dec/funct5_8_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u3974 (
    .a(_al_u3938_o),
    .b(\ins_dec/n149_lutinv ),
    .c(\ins_dec/funct5_8_lutinv ),
    .o(\ins_dec/n151 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3975 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [9]),
    .c(\biu/cache_ctrl_logic/pa_temp [9]),
    .o(\biu/cache_ctrl_logic/n166 [9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3976 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [8]),
    .c(\biu/cache_ctrl_logic/pa_temp [8]),
    .o(\biu/cache_ctrl_logic/n166 [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3977 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [7]),
    .c(\biu/cache_ctrl_logic/pa_temp [7]),
    .o(\biu/cache_ctrl_logic/n166 [7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3978 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [63]),
    .c(\biu/cache_ctrl_logic/pa_temp [63]),
    .o(\biu/cache_ctrl_logic/n166 [63]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3979 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [62]),
    .c(\biu/cache_ctrl_logic/pa_temp [62]),
    .o(\biu/cache_ctrl_logic/n166 [62]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3980 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [61]),
    .c(\biu/cache_ctrl_logic/pa_temp [61]),
    .o(\biu/cache_ctrl_logic/n166 [61]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3981 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [60]),
    .c(\biu/cache_ctrl_logic/pa_temp [60]),
    .o(\biu/cache_ctrl_logic/n166 [60]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3982 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [6]),
    .c(\biu/cache_ctrl_logic/pa_temp [6]),
    .o(\biu/cache_ctrl_logic/n166 [6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3983 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [59]),
    .c(\biu/cache_ctrl_logic/pa_temp [59]),
    .o(\biu/cache_ctrl_logic/n166 [59]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3984 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [58]),
    .c(\biu/cache_ctrl_logic/pa_temp [58]),
    .o(\biu/cache_ctrl_logic/n166 [58]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3985 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [57]),
    .c(\biu/cache_ctrl_logic/pa_temp [57]),
    .o(\biu/cache_ctrl_logic/n166 [57]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3986 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [56]),
    .c(\biu/cache_ctrl_logic/pa_temp [56]),
    .o(\biu/cache_ctrl_logic/n166 [56]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3987 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [55]),
    .c(\biu/cache_ctrl_logic/pa_temp [55]),
    .o(\biu/cache_ctrl_logic/n166 [55]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3988 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [54]),
    .c(\biu/cache_ctrl_logic/pa_temp [54]),
    .o(\biu/cache_ctrl_logic/n166 [54]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3989 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [53]),
    .c(\biu/cache_ctrl_logic/pa_temp [53]),
    .o(\biu/cache_ctrl_logic/n166 [53]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3990 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [52]),
    .c(\biu/cache_ctrl_logic/pa_temp [52]),
    .o(\biu/cache_ctrl_logic/n166 [52]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3991 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [51]),
    .c(\biu/cache_ctrl_logic/pa_temp [51]),
    .o(\biu/cache_ctrl_logic/n166 [51]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3992 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [50]),
    .c(\biu/cache_ctrl_logic/pa_temp [50]),
    .o(\biu/cache_ctrl_logic/n166 [50]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3993 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [5]),
    .c(\biu/cache_ctrl_logic/pa_temp [5]),
    .o(\biu/cache_ctrl_logic/n166 [5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3994 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [49]),
    .c(\biu/cache_ctrl_logic/pa_temp [49]),
    .o(\biu/cache_ctrl_logic/n166 [49]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3995 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [48]),
    .c(\biu/cache_ctrl_logic/pa_temp [48]),
    .o(\biu/cache_ctrl_logic/n166 [48]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3996 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [47]),
    .c(\biu/cache_ctrl_logic/pa_temp [47]),
    .o(\biu/cache_ctrl_logic/n166 [47]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3997 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [46]),
    .c(\biu/cache_ctrl_logic/pa_temp [46]),
    .o(\biu/cache_ctrl_logic/n166 [46]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3998 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [45]),
    .c(\biu/cache_ctrl_logic/pa_temp [45]),
    .o(\biu/cache_ctrl_logic/n166 [45]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u3999 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [44]),
    .c(\biu/cache_ctrl_logic/pa_temp [44]),
    .o(\biu/cache_ctrl_logic/n166 [44]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4000 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [43]),
    .c(\biu/cache_ctrl_logic/pa_temp [43]),
    .o(\biu/cache_ctrl_logic/n166 [43]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4001 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [42]),
    .c(\biu/cache_ctrl_logic/pa_temp [42]),
    .o(\biu/cache_ctrl_logic/n166 [42]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4002 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [41]),
    .c(\biu/cache_ctrl_logic/pa_temp [41]),
    .o(\biu/cache_ctrl_logic/n166 [41]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4003 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [40]),
    .c(\biu/cache_ctrl_logic/pa_temp [40]),
    .o(\biu/cache_ctrl_logic/n166 [40]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4004 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [4]),
    .c(\biu/cache_ctrl_logic/pa_temp [4]),
    .o(\biu/cache_ctrl_logic/n166 [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4005 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [39]),
    .c(\biu/cache_ctrl_logic/pa_temp [39]),
    .o(\biu/cache_ctrl_logic/n166 [39]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4006 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [38]),
    .c(\biu/cache_ctrl_logic/pa_temp [38]),
    .o(\biu/cache_ctrl_logic/n166 [38]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4007 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [37]),
    .c(\biu/cache_ctrl_logic/pa_temp [37]),
    .o(\biu/cache_ctrl_logic/n166 [37]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4008 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [36]),
    .c(\biu/cache_ctrl_logic/pa_temp [36]),
    .o(\biu/cache_ctrl_logic/n166 [36]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4009 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [35]),
    .c(\biu/cache_ctrl_logic/pa_temp [35]),
    .o(\biu/cache_ctrl_logic/n166 [35]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4010 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [34]),
    .c(\biu/cache_ctrl_logic/pa_temp [34]),
    .o(\biu/cache_ctrl_logic/n166 [34]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4011 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [33]),
    .c(\biu/cache_ctrl_logic/pa_temp [33]),
    .o(\biu/cache_ctrl_logic/n166 [33]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4012 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [32]),
    .c(\biu/cache_ctrl_logic/pa_temp [32]),
    .o(\biu/cache_ctrl_logic/n166 [32]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4013 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [31]),
    .c(\biu/cache_ctrl_logic/pa_temp [31]),
    .o(\biu/cache_ctrl_logic/n166 [31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4014 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [30]),
    .c(\biu/cache_ctrl_logic/pa_temp [30]),
    .o(\biu/cache_ctrl_logic/n166 [30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4015 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [3]),
    .c(\biu/cache_ctrl_logic/pa_temp [3]),
    .o(\biu/cache_ctrl_logic/n166 [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4016 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [29]),
    .c(\biu/cache_ctrl_logic/pa_temp [29]),
    .o(\biu/cache_ctrl_logic/n166 [29]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4017 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [28]),
    .c(\biu/cache_ctrl_logic/pa_temp [28]),
    .o(\biu/cache_ctrl_logic/n166 [28]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4018 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [27]),
    .c(\biu/cache_ctrl_logic/pa_temp [27]),
    .o(\biu/cache_ctrl_logic/n166 [27]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4019 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [26]),
    .c(\biu/cache_ctrl_logic/pa_temp [26]),
    .o(\biu/cache_ctrl_logic/n166 [26]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4020 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [25]),
    .c(\biu/cache_ctrl_logic/pa_temp [25]),
    .o(\biu/cache_ctrl_logic/n166 [25]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4021 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [24]),
    .c(\biu/cache_ctrl_logic/pa_temp [24]),
    .o(\biu/cache_ctrl_logic/n166 [24]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4022 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [23]),
    .c(\biu/cache_ctrl_logic/pa_temp [23]),
    .o(\biu/cache_ctrl_logic/n166 [23]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4023 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [22]),
    .c(\biu/cache_ctrl_logic/pa_temp [22]),
    .o(\biu/cache_ctrl_logic/n166 [22]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4024 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [21]),
    .c(\biu/cache_ctrl_logic/pa_temp [21]),
    .o(\biu/cache_ctrl_logic/n166 [21]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4025 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [20]),
    .c(\biu/cache_ctrl_logic/pa_temp [20]),
    .o(\biu/cache_ctrl_logic/n166 [20]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4026 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [2]),
    .c(\biu/cache_ctrl_logic/pa_temp [2]),
    .o(\biu/cache_ctrl_logic/n166 [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4027 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [19]),
    .c(\biu/cache_ctrl_logic/pa_temp [19]),
    .o(\biu/cache_ctrl_logic/n166 [19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4028 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [18]),
    .c(\biu/cache_ctrl_logic/pa_temp [18]),
    .o(\biu/cache_ctrl_logic/n166 [18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4029 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [17]),
    .c(\biu/cache_ctrl_logic/pa_temp [17]),
    .o(\biu/cache_ctrl_logic/n166 [17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4030 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [16]),
    .c(\biu/cache_ctrl_logic/pa_temp [16]),
    .o(\biu/cache_ctrl_logic/n166 [16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4031 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [15]),
    .c(\biu/cache_ctrl_logic/pa_temp [15]),
    .o(\biu/cache_ctrl_logic/n166 [15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4032 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [14]),
    .c(\biu/cache_ctrl_logic/pa_temp [14]),
    .o(\biu/cache_ctrl_logic/n166 [14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4033 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [13]),
    .c(\biu/cache_ctrl_logic/pa_temp [13]),
    .o(\biu/cache_ctrl_logic/n166 [13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4034 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [12]),
    .c(\biu/cache_ctrl_logic/pa_temp [12]),
    .o(\biu/cache_ctrl_logic/n166 [12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4035 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [11]),
    .c(\biu/cache_ctrl_logic/pa_temp [11]),
    .o(\biu/cache_ctrl_logic/n166 [11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4036 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [10]),
    .c(\biu/cache_ctrl_logic/pa_temp [10]),
    .o(\biu/cache_ctrl_logic/n166 [10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4037 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [1]),
    .c(\biu/cache_ctrl_logic/pa_temp [1]),
    .o(\biu/cache_ctrl_logic/n166 [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u4038 (
    .a(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .b(\biu/paddress [0]),
    .c(\biu/cache_ctrl_logic/pa_temp [0]),
    .o(\biu/cache_ctrl_logic/n166 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4039 (
    .a(\exu/alu_data_mem_csr [7]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n1 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4040 (
    .a(\exu/lsu/n1 [7]),
    .b(uncache_data[7]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4041 (
    .a(\exu/alu_data_mem_csr [6]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n1 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4042 (
    .a(\exu/lsu/n1 [6]),
    .b(uncache_data[6]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4043 (
    .a(\exu/alu_data_mem_csr [5]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n1 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4044 (
    .a(\exu/lsu/n1 [5]),
    .b(uncache_data[5]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4045 (
    .a(\exu/alu_data_mem_csr [4]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n1 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4046 (
    .a(\exu/lsu/n1 [4]),
    .b(uncache_data[4]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4047 (
    .a(\exu/alu_data_mem_csr [3]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n1 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4048 (
    .a(\exu/lsu/n1 [3]),
    .b(uncache_data[3]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4049 (
    .a(\exu/alu_data_mem_csr [2]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n1 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4050 (
    .a(\exu/lsu/n1 [2]),
    .b(uncache_data[2]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4051 (
    .a(\exu/alu_data_mem_csr [1]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n1 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4052 (
    .a(\exu/lsu/n1 [1]),
    .b(uncache_data[1]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4053 (
    .a(\exu/alu_data_mem_csr [0]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n1 [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4054 (
    .a(\exu/lsu/n1 [0]),
    .b(uncache_data[0]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u4055 (
    .a(\ins_dec/mux24_b10_sel_is_0_o ),
    .b(_al_u3382_o),
    .c(id_ins[31]),
    .o(_al_u4055_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4056 (
    .a(_al_u4055_o),
    .b(_al_u3214_o),
    .c(id_ins[30]),
    .o(\ins_dec/n291 [19]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4057 (
    .a(_al_u4055_o),
    .b(_al_u3214_o),
    .c(id_ins[29]),
    .o(\ins_dec/n291 [18]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4058 (
    .a(_al_u4055_o),
    .b(_al_u3214_o),
    .c(id_ins[28]),
    .o(\ins_dec/n291 [17]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4059 (
    .a(_al_u4055_o),
    .b(_al_u3214_o),
    .c(id_ins[27]),
    .o(\ins_dec/n291 [16]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4060 (
    .a(_al_u4055_o),
    .b(_al_u3214_o),
    .c(id_ins[26]),
    .o(\ins_dec/n291 [15]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4061 (
    .a(_al_u4055_o),
    .b(_al_u3214_o),
    .c(id_ins[25]),
    .o(\ins_dec/n291 [14]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4062 (
    .a(_al_u4055_o),
    .b(_al_u3214_o),
    .c(id_ins[24]),
    .o(\ins_dec/n291 [13]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u4063 (
    .a(_al_u4055_o),
    .b(_al_u3214_o),
    .c(id_ins[23]),
    .o(\ins_dec/n291 [12]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u4064 (
    .a(_al_u2933_o),
    .b(_al_u2938_o),
    .c(_al_u2939_o),
    .d(_al_u3212_o),
    .o(_al_u4064_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4065 (
    .a(_al_u3213_o),
    .b(_al_u4064_o),
    .o(\ins_dec/mux27_b12_sel_is_0_o ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4066 (
    .a(\ins_dec/mux27_b12_sel_is_0_o ),
    .b(_al_u3214_o),
    .c(id_ins[15]),
    .o(_al_u4066_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(~D*C)))"),
    .INIT(16'h88c8))
    _al_u4067 (
    .a(\ins_dec/mux24_b10_sel_is_0_o ),
    .b(_al_u4066_o),
    .c(\ins_dec/op_store ),
    .d(id_ins[11]),
    .o(_al_u4067_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4068 (
    .a(\ins_dec/op_store ),
    .b(_al_u3214_o),
    .c(_al_u4064_o),
    .o(\ins_dec/mux27_b56_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u4069 (
    .a(\ins_dec/mux27_b56_sel_is_0_o ),
    .b(_al_u4064_o),
    .c(id_ins[24]),
    .d(id_ins[10]),
    .o(_al_u4069_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4070 (
    .a(_al_u4067_o),
    .b(_al_u4069_o),
    .o(\ins_dec/n291 [4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4071 (
    .a(\ins_dec/mux27_b12_sel_is_0_o ),
    .b(_al_u3214_o),
    .c(_al_u3216_o),
    .o(_al_u4071_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(~D*C)))"),
    .INIT(16'h88c8))
    _al_u4072 (
    .a(\ins_dec/mux24_b10_sel_is_0_o ),
    .b(_al_u4071_o),
    .c(\ins_dec/op_store ),
    .d(id_ins[10]),
    .o(_al_u4072_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4073 (
    .a(\ins_dec/mux27_b56_sel_is_0_o ),
    .b(_al_u4064_o),
    .c(id_ins[9]),
    .d(id_ins[23]),
    .o(_al_u4073_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4074 (
    .a(_al_u4072_o),
    .b(_al_u4073_o),
    .o(\ins_dec/n291 [3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4075 (
    .a(\ins_dec/mux27_b12_sel_is_0_o ),
    .b(_al_u3214_o),
    .c(_al_u3217_o),
    .o(_al_u4075_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(~D*C)))"),
    .INIT(16'h88c8))
    _al_u4076 (
    .a(\ins_dec/mux24_b10_sel_is_0_o ),
    .b(_al_u4075_o),
    .c(\ins_dec/op_store ),
    .d(id_ins[9]),
    .o(_al_u4076_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4077 (
    .a(\ins_dec/mux27_b56_sel_is_0_o ),
    .b(_al_u4064_o),
    .c(id_ins[8]),
    .d(id_ins[22]),
    .o(_al_u4077_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4078 (
    .a(_al_u4076_o),
    .b(_al_u4077_o),
    .o(\ins_dec/n291 [2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4079 (
    .a(\ins_dec/mux27_b12_sel_is_0_o ),
    .b(_al_u3214_o),
    .c(_al_u3384_o),
    .o(_al_u4079_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(~D*C)))"),
    .INIT(16'h88c8))
    _al_u4080 (
    .a(\ins_dec/mux24_b10_sel_is_0_o ),
    .b(_al_u4079_o),
    .c(\ins_dec/op_store ),
    .d(id_ins[8]),
    .o(_al_u4080_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u4081 (
    .a(\ins_dec/mux27_b56_sel_is_0_o ),
    .b(_al_u4064_o),
    .c(id_ins[7]),
    .d(id_ins[21]),
    .o(_al_u4081_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4082 (
    .a(_al_u4080_o),
    .b(_al_u4081_o),
    .o(\ins_dec/n291 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4083 (
    .a(\ins_dec/op_store ),
    .b(id_ins[7]),
    .o(_al_u4083_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4084 (
    .a(\ins_dec/op_load ),
    .b(_al_u3213_o),
    .o(_al_u4084_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    _al_u4085 (
    .a(_al_u4083_o),
    .b(_al_u4084_o),
    .c(id_ins[20]),
    .o(\ins_dec/n291 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u4086 (
    .a(\ins_dec/op_store ),
    .b(\ins_dec/op_amo ),
    .c(_al_u3925_o),
    .d(_al_u4064_o),
    .o(_al_u4086_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4087 (
    .a(_al_u4086_o),
    .b(id_ins[24]),
    .o(id_rs2_index[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4088 (
    .a(_al_u4086_o),
    .b(id_ins[23]),
    .o(id_rs2_index[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4089 (
    .a(_al_u4086_o),
    .b(id_ins[22]),
    .o(id_rs2_index[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4090 (
    .a(_al_u4086_o),
    .b(id_ins[21]),
    .o(id_rs2_index[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4091 (
    .a(_al_u4086_o),
    .b(id_ins[20]),
    .o(id_rs2_index[0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4092 (
    .a(\ins_dec/funct6_0_lutinv ),
    .b(_al_u3927_o),
    .c(_al_u3928_o),
    .o(_al_u4092_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4093 (
    .a(_al_u4092_o),
    .b(\ins_dec/n35_lutinv ),
    .c(_al_u3384_o),
    .o(\ins_dec/ins_slli ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4094 (
    .a(\ins_dec/funct7_0_lutinv ),
    .b(\ins_dec/n35_lutinv ),
    .c(_al_u3384_o),
    .o(_al_u4094_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4095 (
    .a(_al_u3927_o),
    .b(_al_u3928_o),
    .o(\ins_dec/op_32_imm_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(B*~(~D*~C)))"),
    .INIT(16'heeea))
    _al_u4096 (
    .a(\ins_dec/ins_slli ),
    .b(_al_u4094_o),
    .c(\ins_dec/op_32_imm_lutinv ),
    .d(_al_u3925_o),
    .o(\ins_dec/n235 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4097 (
    .a(_al_u3939_o),
    .b(id_ins[31]),
    .c(id_ins[29]),
    .o(\ins_dec/n155 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4098 (
    .a(_al_u3939_o),
    .b(id_ins[31]),
    .c(id_ins[29]),
    .o(\ins_dec/n158 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4099 (
    .a(hready_pad),
    .b(hresp_pad),
    .o(_al_u4099_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C)*~(A)+~(D*~B)*C*~(A)+~(~(D*~B))*C*A+~(D*~B)*C*A)"),
    .INIT(16'he4f5))
    _al_u4100 (
    .a(_al_u2890_o),
    .b(_al_u3407_o),
    .c(_al_u4099_o),
    .d(\biu/bus_unit/statu [3]),
    .o(_al_u4100_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B)*~(A)+~C*B*~(A)+~(~C)*B*A+~C*B*A)"),
    .INIT(8'h8d))
    _al_u4101 (
    .a(\biu/bus_unit/mux10_b3_sel_is_0_o ),
    .b(_al_u4100_o),
    .c(hresp_pad),
    .o(_al_u4101_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u4102 (
    .a(_al_u2833_o),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(_al_u4101_o),
    .o(\biu/bus_unit/n35 [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u4103 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(\cu_ru/medeleg [15]),
    .c(wb_st_page_fault),
    .o(\cu_ru/medeleg_exc_ctrl/spf_target_s ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u4104 (
    .a(priv[3]),
    .b(\cu_ru/medeleg [15]),
    .c(wb_st_page_fault),
    .o(\cu_ru/medeleg_exc_ctrl/spf_target_m_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4105 (
    .a(\cu_ru/medeleg_exc_ctrl/spf_target_s ),
    .b(\cu_ru/medeleg_exc_ctrl/spf_target_m_lutinv ),
    .o(\cu_ru/medeleg_exc_ctrl/n85_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u4106 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(priv[3]),
    .c(\cu_ru/medeleg [13]),
    .d(wb_ld_page_fault),
    .o(_al_u4106_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4107 (
    .a(\cu_ru/medeleg_exc_ctrl/n85_neg_lutinv ),
    .b(_al_u4106_o),
    .o(_al_u4107_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4108 (
    .a(\cu_ru/medeleg [7]),
    .b(wb_st_acc_fault),
    .o(_al_u4108_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u4109 (
    .a(priv[3]),
    .b(\cu_ru/medeleg [7]),
    .c(wb_st_acc_fault),
    .o(\cu_ru/medeleg_exc_ctrl/saf_target_m_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u4110 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(_al_u4108_o),
    .c(\cu_ru/medeleg_exc_ctrl/saf_target_m_lutinv ),
    .o(\cu_ru/medeleg_exc_ctrl/n87_neg_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u4111 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(\cu_ru/medeleg [5]),
    .c(wb_ld_acc_fault),
    .o(\cu_ru/medeleg_exc_ctrl/laf_target_s ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u4112 (
    .a(priv[3]),
    .b(\cu_ru/medeleg [5]),
    .c(wb_ld_acc_fault),
    .o(\cu_ru/medeleg_exc_ctrl/laf_target_m_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u4113 (
    .a(_al_u4107_o),
    .b(\cu_ru/medeleg_exc_ctrl/n87_neg_lutinv ),
    .c(\cu_ru/medeleg_exc_ctrl/laf_target_s ),
    .d(\cu_ru/medeleg_exc_ctrl/laf_target_m_lutinv ),
    .o(_al_u4113_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u4114 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(\cu_ru/medeleg [0]),
    .c(wb_ins_addr_mis),
    .o(\cu_ru/medeleg_exc_ctrl/iam_target_s ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u4115 (
    .a(priv[3]),
    .b(\cu_ru/medeleg [0]),
    .c(wb_ins_addr_mis),
    .o(\cu_ru/medeleg_exc_ctrl/iam_target_m_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4116 (
    .a(\cu_ru/medeleg_exc_ctrl/iam_target_s ),
    .b(\cu_ru/medeleg_exc_ctrl/iam_target_m_lutinv ),
    .o(\cu_ru/medeleg_exc_ctrl/n80_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u4117 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(priv[3]),
    .c(\cu_ru/medeleg [2]),
    .d(wb_ill_ins),
    .o(_al_u4117_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4118 (
    .a(\cu_ru/medeleg_exc_ctrl/n80_neg_lutinv ),
    .b(_al_u4117_o),
    .o(\cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4119 (
    .a(\cu_ru/medeleg [1]),
    .b(wb_ins_acc_fault),
    .o(_al_u4119_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u4120 (
    .a(priv[3]),
    .b(\cu_ru/medeleg [1]),
    .c(wb_ins_acc_fault),
    .o(\cu_ru/medeleg_exc_ctrl/iaf_target_m_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u4121 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(_al_u4119_o),
    .c(\cu_ru/medeleg_exc_ctrl/iaf_target_m_lutinv ),
    .o(_al_u4121_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4122 (
    .a(\cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o ),
    .b(_al_u4121_o),
    .o(_al_u4122_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4123 (
    .a(\cu_ru/medeleg [4]),
    .b(wb_ld_addr_mis),
    .o(_al_u4123_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u4124 (
    .a(priv[3]),
    .b(\cu_ru/medeleg [4]),
    .c(wb_ld_addr_mis),
    .o(\cu_ru/medeleg_exc_ctrl/lam_target_m_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u4125 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(_al_u4123_o),
    .c(\cu_ru/medeleg_exc_ctrl/lam_target_m_lutinv ),
    .o(\cu_ru/medeleg_exc_ctrl/n84_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u4126 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(priv[3]),
    .c(\cu_ru/medeleg [6]),
    .d(wb_st_addr_mis),
    .o(_al_u4126_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4127 (
    .a(\cu_ru/medeleg_exc_ctrl/n84_neg_lutinv ),
    .b(_al_u4126_o),
    .o(_al_u4127_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u4128 (
    .a(priv[0]),
    .b(priv[1]),
    .c(wb_ecall),
    .o(_al_u4128_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(C*A))"),
    .INIT(16'h004c))
    _al_u4129 (
    .a(_al_u4113_o),
    .b(_al_u4122_o),
    .c(_al_u4127_o),
    .d(_al_u4128_o),
    .o(\cu_ru/medeleg_exc_ctrl/n98 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4130 (
    .a(\cu_ru/mideleg_int_ctrl/n29_lutinv ),
    .b(_al_u3242_o),
    .o(\cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u4131 (
    .a(\cu_ru/mideleg_int_ctrl/sti_ack_s ),
    .b(\cu_ru/m_sip [5]),
    .c(\cu_ru/mie ),
    .d(\cu_ru/mideleg [5]),
    .o(_al_u4131_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u4132 (
    .a(\cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o ),
    .b(_al_u4131_o),
    .c(_al_u3237_o),
    .o(_al_u4132_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4133 (
    .a(wb_ins_acc_fault),
    .b(wb_ins_addr_mis),
    .c(wb_ins_page_fault),
    .o(_al_u4133_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u4134 (
    .a(_al_u4133_o),
    .b(wb_st_acc_fault),
    .c(wb_st_addr_mis),
    .d(wb_st_page_fault),
    .o(_al_u4134_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u4135 (
    .a(wb_ill_ins),
    .b(wb_ld_acc_fault),
    .c(wb_ld_addr_mis),
    .d(wb_ld_page_fault),
    .o(_al_u4135_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u4136 (
    .a(_al_u4135_o),
    .b(wb_ebreak),
    .c(wb_ecall),
    .o(_al_u4136_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4137 (
    .a(_al_u4134_o),
    .b(_al_u4136_o),
    .o(_al_u4137_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4138 (
    .a(_al_u4137_o),
    .b(wb_valid),
    .o(_al_u4138_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4139 (
    .a(\cu_ru/m_sie [11]),
    .b(\cu_ru/m_sip [11]),
    .c(\cu_ru/mie ),
    .o(_al_u4139_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u4140 (
    .a(_al_u4132_o),
    .b(_al_u4138_o),
    .c(_al_u3238_o),
    .d(_al_u4139_o),
    .o(_al_u4140_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u4141 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(priv[3]),
    .c(\cu_ru/medeleg [3]),
    .d(wb_ebreak),
    .o(_al_u4141_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4142 (
    .a(_al_u4138_o),
    .b(_al_u4141_o),
    .o(_al_u4142_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u4143 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(priv[3]),
    .c(\cu_ru/medeleg [12]),
    .d(wb_ins_page_fault),
    .o(_al_u4143_o));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(C*~(~D*~A)))"),
    .INIT(16'hfcec))
    _al_u4144 (
    .a(\cu_ru/medeleg_exc_ctrl/n98 [2]),
    .b(_al_u4140_o),
    .c(_al_u4142_o),
    .d(_al_u4143_o),
    .o(\cu_ru/trap_cause [2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u4145 (
    .a(\exu/alu_data_mem_csr [7]),
    .b(\exu/alu_data_mem_csr [15]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(\exu/lsu/n4 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4146 (
    .a(\exu/lsu/n4 [15]),
    .b(uncache_data[15]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [15]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u4147 (
    .a(\exu/alu_data_mem_csr [6]),
    .b(\exu/alu_data_mem_csr [14]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(\exu/lsu/n4 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4148 (
    .a(\exu/lsu/n4 [14]),
    .b(uncache_data[14]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [14]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u4149 (
    .a(\exu/alu_data_mem_csr [5]),
    .b(\exu/alu_data_mem_csr [13]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(\exu/lsu/n4 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4150 (
    .a(\exu/lsu/n4 [13]),
    .b(uncache_data[13]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [13]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u4151 (
    .a(\exu/alu_data_mem_csr [4]),
    .b(\exu/alu_data_mem_csr [12]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(\exu/lsu/n4 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4152 (
    .a(\exu/lsu/n4 [12]),
    .b(uncache_data[12]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [12]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u4153 (
    .a(\exu/alu_data_mem_csr [3]),
    .b(\exu/alu_data_mem_csr [11]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(\exu/lsu/n4 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4154 (
    .a(\exu/lsu/n4 [11]),
    .b(uncache_data[11]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [11]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u4155 (
    .a(\exu/alu_data_mem_csr [2]),
    .b(\exu/alu_data_mem_csr [10]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(\exu/lsu/n4 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4156 (
    .a(\exu/lsu/n4 [10]),
    .b(uncache_data[10]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [10]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u4157 (
    .a(\exu/alu_data_mem_csr [9]),
    .b(\exu/alu_data_mem_csr [1]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(\exu/lsu/n4 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4158 (
    .a(\exu/lsu/n4 [9]),
    .b(uncache_data[9]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [9]));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u4159 (
    .a(\exu/alu_data_mem_csr [8]),
    .b(\exu/alu_data_mem_csr [0]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(\exu/lsu/n4 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u4160 (
    .a(\exu/lsu/n4 [8]),
    .b(uncache_data[8]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [8]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4161 (
    .a(\ins_dec/op_store ),
    .b(\ins_dec/op_amo ),
    .o(_al_u4161_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u4162 (
    .a(_al_u4161_o),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .d(_al_u3384_o),
    .o(_al_u4162_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4163 (
    .a(\ins_dec/op_load ),
    .b(_al_u3217_o),
    .c(_al_u3384_o),
    .o(\ins_dec/n48_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*~B*~A)"),
    .INIT(16'hfffe))
    _al_u4164 (
    .a(_al_u4162_o),
    .b(\ins_dec/op_32_reg_lutinv ),
    .c(\ins_dec/op_32_imm_lutinv ),
    .d(\ins_dec/n48_lutinv ),
    .o(\ins_dec/qbyte ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4165 (
    .a(\ins_dec/mux24_b10_sel_is_0_o ),
    .b(_al_u3213_o),
    .o(_al_u4165_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4166 (
    .a(_al_u4165_o),
    .b(id_ins[29]),
    .o(_al_u4166_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4167 (
    .a(_al_u3214_o),
    .b(id_ins[20]),
    .o(_al_u4167_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u4168 (
    .a(_al_u4166_o),
    .b(_al_u4167_o),
    .c(_al_u4064_o),
    .d(id_ins[28]),
    .o(\ins_dec/n291 [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4169 (
    .a(_al_u4165_o),
    .b(id_ins[28]),
    .o(_al_u4169_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4170 (
    .a(_al_u3214_o),
    .b(id_ins[19]),
    .o(_al_u4170_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u4171 (
    .a(_al_u4169_o),
    .b(_al_u4170_o),
    .c(_al_u4064_o),
    .d(id_ins[27]),
    .o(\ins_dec/n291 [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4172 (
    .a(_al_u4165_o),
    .b(id_ins[27]),
    .o(_al_u4172_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4173 (
    .a(_al_u3214_o),
    .b(id_ins[18]),
    .o(_al_u4173_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u4174 (
    .a(_al_u4172_o),
    .b(_al_u4173_o),
    .c(_al_u4064_o),
    .d(id_ins[26]),
    .o(\ins_dec/n291 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4175 (
    .a(_al_u3214_o),
    .b(_al_u4064_o),
    .c(id_ins[25]),
    .d(id_ins[17]),
    .o(_al_u4175_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u4176 (
    .a(_al_u4165_o),
    .b(_al_u4175_o),
    .c(id_ins[26]),
    .o(\ins_dec/n291 [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4177 (
    .a(_al_u4165_o),
    .b(id_ins[25]),
    .o(_al_u4177_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4178 (
    .a(_al_u3214_o),
    .b(id_ins[16]),
    .o(_al_u4178_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u4179 (
    .a(_al_u4177_o),
    .b(_al_u4178_o),
    .c(_al_u4064_o),
    .d(id_ins[11]),
    .o(\ins_dec/n291 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4180 (
    .a(_al_u3214_o),
    .b(id_ins[22]),
    .o(_al_u4180_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'hfbea))
    _al_u4181 (
    .a(_al_u4180_o),
    .b(_al_u4064_o),
    .c(id_ins[30]),
    .d(_al_u4055_o),
    .o(\ins_dec/n291 [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4182 (
    .a(_al_u4165_o),
    .b(id_ins[30]),
    .o(_al_u4182_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4183 (
    .a(_al_u3214_o),
    .b(id_ins[21]),
    .o(_al_u4183_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u4184 (
    .a(_al_u4182_o),
    .b(_al_u4183_o),
    .c(_al_u4064_o),
    .d(id_ins[29]),
    .o(\ins_dec/n291 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u4185 (
    .a(_al_u3926_o),
    .b(\ins_dec/funct3_0_lutinv ),
    .c(_al_u3927_o),
    .o(_al_u4185_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*~B*~A)"),
    .INIT(16'hfffe))
    _al_u4186 (
    .a(_al_u4185_o),
    .b(\ins_dec/ins_addw ),
    .c(\ins_dec/n59 ),
    .d(_al_u3955_o),
    .o(\ins_dec/n132 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u4187 (
    .a(id_system),
    .b(_al_u3217_o),
    .c(_al_u3384_o),
    .o(\ins_dec/n239 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u4188 (
    .a(id_system),
    .b(_al_u3217_o),
    .c(_al_u3384_o),
    .o(\ins_dec/n141_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D*C*A))"),
    .INIT(16'heccc))
    _al_u4189 (
    .a(_al_u3938_o),
    .b(\ins_dec/n141_lutinv ),
    .c(_al_u3399_o),
    .d(id_ins[27]),
    .o(\ins_dec/n145 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4190 (
    .a(_al_u3407_o),
    .b(\biu/bus_unit/statu [0]),
    .o(\biu/bus_unit/n26 [0]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(B)*~((~C*A))+~D*B*~((~C*A))+~(~D)*B*(~C*A)+~D*B*(~C*A))"),
    .INIT(16'hf702))
    _al_u4191 (
    .a(\biu/bus_unit/mux10_b3_sel_is_0_o ),
    .b(\biu/bus_unit/n26 [0]),
    .c(_al_u2890_o),
    .d(_al_u4099_o),
    .o(_al_u4191_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'hcc80))
    _al_u4192 (
    .a(\biu/bus_unit/n15_lutinv ),
    .b(htrans_pad[0]),
    .c(hready_pad),
    .d(hresp_pad),
    .o(_al_u4192_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u4193 (
    .a(_al_u4191_o),
    .b(_al_u2957_o),
    .c(_al_u4192_o),
    .o(_al_u4193_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u4194 (
    .a(_al_u2833_o),
    .b(\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ),
    .c(\biu/cache_ctrl_logic/n75_lutinv ),
    .d(_al_u2885_o),
    .o(_al_u4194_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u4195 (
    .a(\biu/bus_unit/mmu/statu [1]),
    .b(\biu/bus_unit/mmu/statu [2]),
    .c(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u4195_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4196 (
    .a(_al_u3411_o),
    .b(_al_u4195_o),
    .o(\biu/bus_unit/mmu/mux10_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4197 (
    .a(_al_u2704_o),
    .b(\biu/bus_unit/mmu/mux10_b0_sel_is_2_o ),
    .c(\biu/bus_unit/statu [0]),
    .o(_al_u4197_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~C*~(~D*~A)))"),
    .INIT(16'h3031))
    _al_u4198 (
    .a(_al_u4193_o),
    .b(_al_u4194_o),
    .c(_al_u4197_o),
    .d(_al_u2958_o),
    .o(\biu/bus_unit/n35 [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4199 (
    .a(_al_u2903_o),
    .b(_al_u2905_o),
    .c(_al_u2907_o),
    .o(_al_u4199_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4200 (
    .a(_al_u2891_o),
    .b(_al_u2893_o),
    .o(_al_u4200_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4201 (
    .a(_al_u2895_o),
    .b(_al_u2897_o),
    .c(_al_u2899_o),
    .d(_al_u2901_o),
    .o(_al_u4201_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u4202 (
    .a(\biu/cache_ctrl_logic/n149 ),
    .b(_al_u4199_o),
    .c(_al_u4200_o),
    .d(_al_u4201_o),
    .o(\biu/cache_ctrl_logic/n140 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4203 (
    .a(\exu/alu_data_mem_csr [17]),
    .b(\exu/alu_data_mem_csr [1]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4203_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4204 (
    .a(addr_ex[0]),
    .b(addr_ex[1]),
    .o(\exu/lsu/n2_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u4205 (
    .a(_al_u4203_o),
    .b(\exu/alu_data_mem_csr [9]),
    .c(\exu/lsu/n2_lutinv ),
    .o(_al_u4205_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4206 (
    .a(_al_u4205_o),
    .b(uncache_data[17]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [17]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4207 (
    .a(\exu/alu_data_mem_csr [16]),
    .b(\exu/alu_data_mem_csr [0]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4207_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u4208 (
    .a(_al_u4207_o),
    .b(\exu/alu_data_mem_csr [8]),
    .c(\exu/lsu/n2_lutinv ),
    .o(_al_u4208_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4209 (
    .a(_al_u4208_o),
    .b(uncache_data[16]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [16]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u4210 (
    .a(\exu/alu_data_mem_csr [7]),
    .b(\exu/alu_data_mem_csr [15]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4210_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4211 (
    .a(_al_u4210_o),
    .b(\exu/alu_data_mem_csr [23]),
    .c(\exu/lsu/n0_lutinv ),
    .o(_al_u4211_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4212 (
    .a(_al_u4211_o),
    .b(uncache_data[23]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u4213 (
    .a(\exu/alu_data_mem_csr [6]),
    .b(\exu/alu_data_mem_csr [14]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4213_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4214 (
    .a(_al_u4213_o),
    .b(\exu/alu_data_mem_csr [22]),
    .c(\exu/lsu/n0_lutinv ),
    .o(_al_u4214_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4215 (
    .a(_al_u4214_o),
    .b(uncache_data[22]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [22]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u4216 (
    .a(\exu/alu_data_mem_csr [5]),
    .b(\exu/alu_data_mem_csr [13]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4216_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4217 (
    .a(_al_u4216_o),
    .b(\exu/alu_data_mem_csr [21]),
    .c(\exu/lsu/n0_lutinv ),
    .o(_al_u4217_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4218 (
    .a(_al_u4217_o),
    .b(uncache_data[21]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u4219 (
    .a(\exu/alu_data_mem_csr [4]),
    .b(\exu/alu_data_mem_csr [12]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4219_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4220 (
    .a(_al_u4219_o),
    .b(\exu/alu_data_mem_csr [20]),
    .c(\exu/lsu/n0_lutinv ),
    .o(_al_u4220_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4221 (
    .a(_al_u4220_o),
    .b(uncache_data[20]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [20]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u4222 (
    .a(\exu/alu_data_mem_csr [3]),
    .b(\exu/alu_data_mem_csr [11]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4222_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4223 (
    .a(_al_u4222_o),
    .b(\exu/alu_data_mem_csr [19]),
    .c(\exu/lsu/n0_lutinv ),
    .o(_al_u4223_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4224 (
    .a(_al_u4223_o),
    .b(uncache_data[19]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [19]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u4225 (
    .a(\exu/alu_data_mem_csr [2]),
    .b(\exu/alu_data_mem_csr [10]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4225_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4226 (
    .a(_al_u4225_o),
    .b(\exu/alu_data_mem_csr [18]),
    .c(\exu/lsu/n0_lutinv ),
    .o(_al_u4226_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4227 (
    .a(_al_u4226_o),
    .b(uncache_data[18]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [18]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u4228 (
    .a(\ins_dec/mux27_b56_sel_is_0_o ),
    .b(id_ins[31]),
    .o(\ins_dec/n291 [56]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4229 (
    .a(priv[1]),
    .b(wb_ecall),
    .o(_al_u4229_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*B*~A))"),
    .INIT(16'h0f0b))
    _al_u4230 (
    .a(_al_u4113_o),
    .b(_al_u4127_o),
    .c(_al_u4229_o),
    .d(_al_u4128_o),
    .o(_al_u4230_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u4231 (
    .a(_al_u4230_o),
    .b(\cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o ),
    .c(_al_u4143_o),
    .d(_al_u4121_o),
    .o(\cu_ru/medeleg_exc_ctrl/n99 [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u4232 (
    .a(\cu_ru/medeleg_exc_ctrl/n99 [0]),
    .b(_al_u4138_o),
    .c(_al_u4141_o),
    .o(_al_u4232_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4233 (
    .a(\cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ),
    .b(_al_u4139_o),
    .o(_al_u4233_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u4234 (
    .a(_al_u4138_o),
    .b(\cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o ),
    .c(_al_u4131_o),
    .d(_al_u4233_o),
    .o(_al_u4234_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u4235 (
    .a(_al_u4232_o),
    .b(_al_u4234_o),
    .o(\cu_ru/trap_cause [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4236 (
    .a(\exu/alu_data_mem_csr [55]),
    .b(\exu/alu_data_mem_csr [47]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4236_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4237 (
    .a(\exu/alu_data_mem_csr [63]),
    .b(\exu/alu_data_mem_csr [39]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4237_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4238 (
    .a(_al_u4236_o),
    .b(_al_u4237_o),
    .o(_al_u4238_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4239 (
    .a(_al_u4238_o),
    .b(uncache_data[63]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [63]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4240 (
    .a(\exu/alu_data_mem_csr [62]),
    .b(\exu/alu_data_mem_csr [46]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4240_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4241 (
    .a(\exu/alu_data_mem_csr [54]),
    .b(\exu/alu_data_mem_csr [38]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4241_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4242 (
    .a(_al_u4240_o),
    .b(_al_u4241_o),
    .o(_al_u4242_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4243 (
    .a(_al_u4242_o),
    .b(uncache_data[62]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [62]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4244 (
    .a(\exu/alu_data_mem_csr [53]),
    .b(\exu/alu_data_mem_csr [45]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4244_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4245 (
    .a(\exu/alu_data_mem_csr [61]),
    .b(\exu/alu_data_mem_csr [37]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4245_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4246 (
    .a(_al_u4244_o),
    .b(_al_u4245_o),
    .o(_al_u4246_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4247 (
    .a(_al_u4246_o),
    .b(uncache_data[61]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [61]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4248 (
    .a(\exu/alu_data_mem_csr [52]),
    .b(\exu/alu_data_mem_csr [44]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4248_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4249 (
    .a(\exu/alu_data_mem_csr [60]),
    .b(\exu/alu_data_mem_csr [36]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4249_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4250 (
    .a(_al_u4248_o),
    .b(_al_u4249_o),
    .o(_al_u4250_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4251 (
    .a(_al_u4250_o),
    .b(uncache_data[60]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [60]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4252 (
    .a(\exu/alu_data_mem_csr [59]),
    .b(\exu/alu_data_mem_csr [43]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4252_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4253 (
    .a(\exu/alu_data_mem_csr [51]),
    .b(\exu/alu_data_mem_csr [35]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4253_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4254 (
    .a(_al_u4252_o),
    .b(_al_u4253_o),
    .o(_al_u4254_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4255 (
    .a(_al_u4254_o),
    .b(uncache_data[59]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [59]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4256 (
    .a(\exu/alu_data_mem_csr [58]),
    .b(\exu/alu_data_mem_csr [42]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4256_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4257 (
    .a(\exu/alu_data_mem_csr [50]),
    .b(\exu/alu_data_mem_csr [34]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4257_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4258 (
    .a(_al_u4256_o),
    .b(_al_u4257_o),
    .o(_al_u4258_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4259 (
    .a(_al_u4258_o),
    .b(uncache_data[58]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [58]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4260 (
    .a(\exu/alu_data_mem_csr [49]),
    .b(\exu/alu_data_mem_csr [41]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4260_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4261 (
    .a(\exu/alu_data_mem_csr [57]),
    .b(\exu/alu_data_mem_csr [33]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4261_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4262 (
    .a(_al_u4260_o),
    .b(_al_u4261_o),
    .o(_al_u4262_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4263 (
    .a(_al_u4262_o),
    .b(uncache_data[57]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [57]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4264 (
    .a(\exu/alu_data_mem_csr [56]),
    .b(\exu/alu_data_mem_csr [40]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4264_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4265 (
    .a(\exu/alu_data_mem_csr [48]),
    .b(\exu/alu_data_mem_csr [32]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4265_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4266 (
    .a(_al_u4264_o),
    .b(_al_u4265_o),
    .o(_al_u4266_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4267 (
    .a(_al_u4266_o),
    .b(uncache_data[56]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [56]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4268 (
    .a(\exu/alu_data_mem_csr [47]),
    .b(\exu/alu_data_mem_csr [39]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4268_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4269 (
    .a(\exu/alu_data_mem_csr [55]),
    .b(\exu/alu_data_mem_csr [31]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4269_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4270 (
    .a(_al_u4268_o),
    .b(_al_u4269_o),
    .o(_al_u4270_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4271 (
    .a(_al_u4270_o),
    .b(uncache_data[55]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [55]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4272 (
    .a(\exu/alu_data_mem_csr [54]),
    .b(\exu/alu_data_mem_csr [38]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4272_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4273 (
    .a(\exu/alu_data_mem_csr [46]),
    .b(\exu/alu_data_mem_csr [30]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4273_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4274 (
    .a(_al_u4272_o),
    .b(_al_u4273_o),
    .o(_al_u4274_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4275 (
    .a(_al_u4274_o),
    .b(uncache_data[54]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [54]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4276 (
    .a(\exu/alu_data_mem_csr [53]),
    .b(\exu/alu_data_mem_csr [37]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4276_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4277 (
    .a(\exu/alu_data_mem_csr [45]),
    .b(\exu/alu_data_mem_csr [29]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4277_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4278 (
    .a(_al_u4276_o),
    .b(_al_u4277_o),
    .o(_al_u4278_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4279 (
    .a(_al_u4278_o),
    .b(uncache_data[53]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [53]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4280 (
    .a(\exu/alu_data_mem_csr [52]),
    .b(\exu/alu_data_mem_csr [36]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4280_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4281 (
    .a(\exu/alu_data_mem_csr [44]),
    .b(\exu/alu_data_mem_csr [28]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4281_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4282 (
    .a(_al_u4280_o),
    .b(_al_u4281_o),
    .o(_al_u4282_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4283 (
    .a(_al_u4282_o),
    .b(uncache_data[52]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [52]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4284 (
    .a(\exu/alu_data_mem_csr [51]),
    .b(\exu/alu_data_mem_csr [35]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4284_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4285 (
    .a(\exu/alu_data_mem_csr [43]),
    .b(\exu/alu_data_mem_csr [27]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4285_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4286 (
    .a(_al_u4284_o),
    .b(_al_u4285_o),
    .o(_al_u4286_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4287 (
    .a(_al_u4286_o),
    .b(uncache_data[51]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [51]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4288 (
    .a(\exu/alu_data_mem_csr [50]),
    .b(\exu/alu_data_mem_csr [34]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4288_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4289 (
    .a(\exu/alu_data_mem_csr [42]),
    .b(\exu/alu_data_mem_csr [26]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4289_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4290 (
    .a(_al_u4288_o),
    .b(_al_u4289_o),
    .o(_al_u4290_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4291 (
    .a(_al_u4290_o),
    .b(uncache_data[50]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [50]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4292 (
    .a(\exu/alu_data_mem_csr [41]),
    .b(\exu/alu_data_mem_csr [33]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4292_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4293 (
    .a(\exu/alu_data_mem_csr [49]),
    .b(\exu/alu_data_mem_csr [25]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4293_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4294 (
    .a(_al_u4292_o),
    .b(_al_u4293_o),
    .o(_al_u4294_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4295 (
    .a(_al_u4294_o),
    .b(uncache_data[49]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [49]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4296 (
    .a(\exu/alu_data_mem_csr [40]),
    .b(\exu/alu_data_mem_csr [32]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4296_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4297 (
    .a(\exu/alu_data_mem_csr [48]),
    .b(\exu/alu_data_mem_csr [24]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4297_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4298 (
    .a(_al_u4296_o),
    .b(_al_u4297_o),
    .o(_al_u4298_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4299 (
    .a(_al_u4298_o),
    .b(uncache_data[48]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [48]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4300 (
    .a(\exu/alu_data_mem_csr [47]),
    .b(\exu/alu_data_mem_csr [31]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4300_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4301 (
    .a(\exu/alu_data_mem_csr [39]),
    .b(\exu/alu_data_mem_csr [23]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4301_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4302 (
    .a(_al_u4300_o),
    .b(_al_u4301_o),
    .o(_al_u4302_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4303 (
    .a(_al_u4302_o),
    .b(uncache_data[47]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [47]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4304 (
    .a(\exu/alu_data_mem_csr [38]),
    .b(\exu/alu_data_mem_csr [30]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4304_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4305 (
    .a(\exu/alu_data_mem_csr [46]),
    .b(\exu/alu_data_mem_csr [22]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4305_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4306 (
    .a(_al_u4304_o),
    .b(_al_u4305_o),
    .o(_al_u4306_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4307 (
    .a(_al_u4306_o),
    .b(uncache_data[46]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [46]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4308 (
    .a(\exu/alu_data_mem_csr [45]),
    .b(\exu/alu_data_mem_csr [29]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4308_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4309 (
    .a(\exu/alu_data_mem_csr [37]),
    .b(\exu/alu_data_mem_csr [21]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4309_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4310 (
    .a(_al_u4308_o),
    .b(_al_u4309_o),
    .o(_al_u4310_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4311 (
    .a(_al_u4310_o),
    .b(uncache_data[45]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [45]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4312 (
    .a(\exu/alu_data_mem_csr [44]),
    .b(\exu/alu_data_mem_csr [28]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4312_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4313 (
    .a(\exu/alu_data_mem_csr [36]),
    .b(\exu/alu_data_mem_csr [20]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4313_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4314 (
    .a(_al_u4312_o),
    .b(_al_u4313_o),
    .o(_al_u4314_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4315 (
    .a(_al_u4314_o),
    .b(uncache_data[44]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [44]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4316 (
    .a(\exu/alu_data_mem_csr [35]),
    .b(\exu/alu_data_mem_csr [27]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4316_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4317 (
    .a(\exu/alu_data_mem_csr [43]),
    .b(\exu/alu_data_mem_csr [19]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4317_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4318 (
    .a(_al_u4316_o),
    .b(_al_u4317_o),
    .o(_al_u4318_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4319 (
    .a(_al_u4318_o),
    .b(uncache_data[43]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [43]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4320 (
    .a(\exu/alu_data_mem_csr [34]),
    .b(\exu/alu_data_mem_csr [26]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4320_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4321 (
    .a(\exu/alu_data_mem_csr [42]),
    .b(\exu/alu_data_mem_csr [18]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4321_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4322 (
    .a(_al_u4320_o),
    .b(_al_u4321_o),
    .o(_al_u4322_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4323 (
    .a(_al_u4322_o),
    .b(uncache_data[42]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [42]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4324 (
    .a(\exu/alu_data_mem_csr [33]),
    .b(\exu/alu_data_mem_csr [25]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4324_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4325 (
    .a(\exu/alu_data_mem_csr [41]),
    .b(\exu/alu_data_mem_csr [17]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4325_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4326 (
    .a(_al_u4324_o),
    .b(_al_u4325_o),
    .o(_al_u4326_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4327 (
    .a(_al_u4326_o),
    .b(uncache_data[41]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [41]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4328 (
    .a(\exu/alu_data_mem_csr [40]),
    .b(\exu/alu_data_mem_csr [24]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4328_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4329 (
    .a(\exu/alu_data_mem_csr [32]),
    .b(\exu/alu_data_mem_csr [16]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4329_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4330 (
    .a(_al_u4328_o),
    .b(_al_u4329_o),
    .o(_al_u4330_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4331 (
    .a(_al_u4330_o),
    .b(uncache_data[40]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [40]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4332 (
    .a(\exu/alu_data_mem_csr [31]),
    .b(\exu/alu_data_mem_csr [23]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4332_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4333 (
    .a(\exu/alu_data_mem_csr [39]),
    .b(\exu/alu_data_mem_csr [15]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4333_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4334 (
    .a(_al_u4332_o),
    .b(_al_u4333_o),
    .o(_al_u4334_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4335 (
    .a(_al_u4334_o),
    .b(uncache_data[39]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [39]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4336 (
    .a(\exu/alu_data_mem_csr [30]),
    .b(\exu/alu_data_mem_csr [22]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4336_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4337 (
    .a(\exu/alu_data_mem_csr [38]),
    .b(\exu/alu_data_mem_csr [14]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4337_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4338 (
    .a(_al_u4336_o),
    .b(_al_u4337_o),
    .o(_al_u4338_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4339 (
    .a(_al_u4338_o),
    .b(uncache_data[38]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [38]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4340 (
    .a(\exu/alu_data_mem_csr [29]),
    .b(\exu/alu_data_mem_csr [21]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4340_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4341 (
    .a(\exu/alu_data_mem_csr [37]),
    .b(\exu/alu_data_mem_csr [13]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4341_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4342 (
    .a(_al_u4340_o),
    .b(_al_u4341_o),
    .o(_al_u4342_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4343 (
    .a(_al_u4342_o),
    .b(uncache_data[37]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [37]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4344 (
    .a(\exu/alu_data_mem_csr [28]),
    .b(\exu/alu_data_mem_csr [20]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4344_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4345 (
    .a(\exu/alu_data_mem_csr [36]),
    .b(\exu/alu_data_mem_csr [12]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4345_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4346 (
    .a(_al_u4344_o),
    .b(_al_u4345_o),
    .o(_al_u4346_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4347 (
    .a(_al_u4346_o),
    .b(uncache_data[36]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [36]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4348 (
    .a(\exu/alu_data_mem_csr [27]),
    .b(\exu/alu_data_mem_csr [19]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4348_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4349 (
    .a(\exu/alu_data_mem_csr [35]),
    .b(\exu/alu_data_mem_csr [11]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4349_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4350 (
    .a(_al_u4348_o),
    .b(_al_u4349_o),
    .o(_al_u4350_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4351 (
    .a(_al_u4350_o),
    .b(uncache_data[35]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [35]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4352 (
    .a(\exu/alu_data_mem_csr [34]),
    .b(\exu/alu_data_mem_csr [18]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4352_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4353 (
    .a(\exu/alu_data_mem_csr [26]),
    .b(\exu/alu_data_mem_csr [10]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4353_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4354 (
    .a(_al_u4352_o),
    .b(_al_u4353_o),
    .o(_al_u4354_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4355 (
    .a(_al_u4354_o),
    .b(uncache_data[34]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [34]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4356 (
    .a(\exu/alu_data_mem_csr [33]),
    .b(\exu/alu_data_mem_csr [17]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4356_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u4357 (
    .a(\exu/alu_data_mem_csr [9]),
    .b(\exu/alu_data_mem_csr [25]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4357_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4358 (
    .a(_al_u4356_o),
    .b(_al_u4357_o),
    .o(_al_u4358_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4359 (
    .a(_al_u4358_o),
    .b(uncache_data[33]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [33]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4360 (
    .a(\exu/alu_data_mem_csr [24]),
    .b(\exu/alu_data_mem_csr [16]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4360_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u4361 (
    .a(\exu/alu_data_mem_csr [8]),
    .b(\exu/alu_data_mem_csr [32]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4361_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4362 (
    .a(_al_u4360_o),
    .b(_al_u4361_o),
    .o(_al_u4362_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4363 (
    .a(_al_u4362_o),
    .b(uncache_data[32]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [32]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4364 (
    .a(\exu/alu_data_mem_csr [31]),
    .b(\exu/alu_data_mem_csr [15]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4364_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u4365 (
    .a(\exu/alu_data_mem_csr [7]),
    .b(\exu/alu_data_mem_csr [23]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4365_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4366 (
    .a(_al_u4364_o),
    .b(_al_u4365_o),
    .o(_al_u4366_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4367 (
    .a(_al_u4366_o),
    .b(uncache_data[31]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [31]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4368 (
    .a(\exu/alu_data_mem_csr [22]),
    .b(\exu/alu_data_mem_csr [14]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4368_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u4369 (
    .a(\exu/alu_data_mem_csr [6]),
    .b(\exu/alu_data_mem_csr [30]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4369_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4370 (
    .a(_al_u4368_o),
    .b(_al_u4369_o),
    .o(_al_u4370_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4371 (
    .a(_al_u4370_o),
    .b(uncache_data[30]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [30]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4372 (
    .a(\exu/alu_data_mem_csr [29]),
    .b(\exu/alu_data_mem_csr [13]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4372_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u4373 (
    .a(\exu/alu_data_mem_csr [5]),
    .b(\exu/alu_data_mem_csr [21]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4373_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4374 (
    .a(_al_u4372_o),
    .b(_al_u4373_o),
    .o(_al_u4374_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4375 (
    .a(_al_u4374_o),
    .b(uncache_data[29]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [29]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u4376 (
    .a(\exu/alu_data_mem_csr [20]),
    .b(\exu/alu_data_mem_csr [12]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4376_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u4377 (
    .a(\exu/alu_data_mem_csr [4]),
    .b(\exu/alu_data_mem_csr [28]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4377_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4378 (
    .a(_al_u4376_o),
    .b(_al_u4377_o),
    .o(_al_u4378_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4379 (
    .a(_al_u4378_o),
    .b(uncache_data[28]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [28]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4380 (
    .a(\exu/alu_data_mem_csr [27]),
    .b(\exu/alu_data_mem_csr [11]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4380_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u4381 (
    .a(\exu/alu_data_mem_csr [3]),
    .b(\exu/alu_data_mem_csr [19]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4381_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4382 (
    .a(_al_u4380_o),
    .b(_al_u4381_o),
    .o(_al_u4382_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4383 (
    .a(_al_u4382_o),
    .b(uncache_data[27]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [27]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u4384 (
    .a(\exu/alu_data_mem_csr [26]),
    .b(\exu/alu_data_mem_csr [10]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4384_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u4385 (
    .a(\exu/alu_data_mem_csr [2]),
    .b(\exu/alu_data_mem_csr [18]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4385_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4386 (
    .a(_al_u4384_o),
    .b(_al_u4385_o),
    .o(_al_u4386_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4387 (
    .a(_al_u4386_o),
    .b(uncache_data[26]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [26]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u4388 (
    .a(\exu/alu_data_mem_csr [9]),
    .b(\exu/alu_data_mem_csr [25]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4388_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u4389 (
    .a(\exu/alu_data_mem_csr [17]),
    .b(\exu/alu_data_mem_csr [1]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4389_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4390 (
    .a(_al_u4388_o),
    .b(_al_u4389_o),
    .o(_al_u4390_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4391 (
    .a(_al_u4390_o),
    .b(uncache_data[25]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [25]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u4392 (
    .a(\exu/alu_data_mem_csr [8]),
    .b(\exu/alu_data_mem_csr [16]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4392_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u4393 (
    .a(\exu/alu_data_mem_csr [24]),
    .b(\exu/alu_data_mem_csr [0]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u4393_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u4394 (
    .a(_al_u4392_o),
    .b(_al_u4393_o),
    .o(_al_u4394_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u4395 (
    .a(_al_u4394_o),
    .b(uncache_data[24]),
    .c(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .o(\biu/l1i_in [24]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u4396 (
    .a(\ins_dec/qbyte ),
    .b(_al_u3919_o),
    .c(_al_u3217_o),
    .o(\ins_dec/obyte ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4397 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [9]),
    .d(\biu/cache_ctrl_logic/l1i_pa [73]),
    .o(_al_u4397_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4398 (
    .a(_al_u4397_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[9]),
    .o(_al_u4398_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u4399 (
    .a(_al_u2847_o),
    .b(\biu/cache_ctrl_logic/statu [2]),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(_al_u4399_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4400 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [9]),
    .d(\biu/cache_ctrl_logic/l1d_pa [73]),
    .o(_al_u4400_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4401 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [73]),
    .d(addr_ex[9]),
    .o(_al_u4401_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4402 (
    .a(_al_u4398_o),
    .b(_al_u4400_o),
    .c(_al_u4401_o),
    .o(_al_u4402_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4403 (
    .a(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .b(\biu/cache_ctrl_logic/n204_lutinv ),
    .o(_al_u4403_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4404 (
    .a(_al_u4402_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [9]),
    .o(\biu/maddress [9]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4405 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [72]),
    .d(\biu/cache_ctrl_logic/pa_temp [72]),
    .o(_al_u4405_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4406 (
    .a(_al_u4405_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[8]),
    .o(_al_u4406_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4407 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [72]),
    .d(addr_ex[8]),
    .o(_al_u4407_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4408 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [8]),
    .d(\biu/cache_ctrl_logic/n212 [8]),
    .o(_al_u4408_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4409 (
    .a(_al_u4406_o),
    .b(_al_u4407_o),
    .c(_al_u4408_o),
    .o(_al_u4409_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4410 (
    .a(_al_u4409_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [8]),
    .o(\biu/maddress [8]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4411 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [71]),
    .d(addr_ex[7]),
    .o(_al_u4411_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4412 (
    .a(_al_u4411_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[7]),
    .o(_al_u4412_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4413 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [7]),
    .d(\biu/cache_ctrl_logic/n212 [7]),
    .o(_al_u4413_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4414 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [71]),
    .d(\biu/cache_ctrl_logic/pa_temp [71]),
    .o(_al_u4414_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4415 (
    .a(_al_u4412_o),
    .b(_al_u4413_o),
    .c(_al_u4414_o),
    .o(_al_u4415_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4416 (
    .a(_al_u4415_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [7]),
    .o(\biu/maddress [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4417 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [127]),
    .d(\biu/cache_ctrl_logic/pa_temp [127]),
    .o(_al_u4417_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4418 (
    .a(_al_u4417_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[63]),
    .o(_al_u4418_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4419 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [127]),
    .d(addr_ex[63]),
    .o(_al_u4419_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4420 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [63]),
    .d(\biu/cache_ctrl_logic/n212 [63]),
    .o(_al_u4420_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4421 (
    .a(_al_u4418_o),
    .b(_al_u4419_o),
    .c(_al_u4420_o),
    .o(_al_u4421_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4422 (
    .a(_al_u4421_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [63]),
    .o(\biu/maddress [63]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4423 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [62]),
    .d(addr_ex[62]),
    .o(_al_u4423_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4424 (
    .a(_al_u4423_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[62]),
    .o(_al_u4424_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4425 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [62]),
    .d(\biu/cache_ctrl_logic/l1i_pa [126]),
    .o(_al_u4425_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4426 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [126]),
    .d(\biu/cache_ctrl_logic/pa_temp [126]),
    .o(_al_u4426_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4427 (
    .a(_al_u4424_o),
    .b(_al_u4425_o),
    .c(_al_u4426_o),
    .o(_al_u4427_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4428 (
    .a(_al_u4427_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [62]),
    .o(\biu/maddress [62]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4429 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [61]),
    .d(\biu/cache_ctrl_logic/l1i_pa [125]),
    .o(_al_u4429_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4430 (
    .a(_al_u4429_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[61]),
    .o(_al_u4430_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4431 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [61]),
    .d(addr_ex[61]),
    .o(_al_u4431_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4432 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [125]),
    .d(\biu/cache_ctrl_logic/pa_temp [125]),
    .o(_al_u4432_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4433 (
    .a(_al_u4430_o),
    .b(_al_u4431_o),
    .c(_al_u4432_o),
    .o(_al_u4433_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4434 (
    .a(_al_u4433_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [61]),
    .o(\biu/maddress [61]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4435 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [60]),
    .d(\biu/cache_ctrl_logic/n212 [60]),
    .o(_al_u4435_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4436 (
    .a(_al_u4435_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[60]),
    .o(_al_u4436_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4437 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [124]),
    .d(addr_ex[60]),
    .o(_al_u4437_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4438 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [124]),
    .d(\biu/cache_ctrl_logic/pa_temp [124]),
    .o(_al_u4438_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4439 (
    .a(_al_u4436_o),
    .b(_al_u4437_o),
    .c(_al_u4438_o),
    .o(_al_u4439_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4440 (
    .a(_al_u4439_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [60]),
    .o(\biu/maddress [60]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4441 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [6]),
    .d(addr_ex[6]),
    .o(_al_u4441_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4442 (
    .a(_al_u4441_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[6]),
    .o(_al_u4442_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4443 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/n212 [6]),
    .d(\biu/cache_ctrl_logic/l1d_pa [70]),
    .o(_al_u4443_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4444 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [70]),
    .d(\biu/cache_ctrl_logic/pa_temp [70]),
    .o(_al_u4444_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4445 (
    .a(_al_u4442_o),
    .b(_al_u4443_o),
    .c(_al_u4444_o),
    .o(_al_u4445_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4446 (
    .a(_al_u4445_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [6]),
    .o(\biu/maddress [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4447 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [59]),
    .d(\biu/cache_ctrl_logic/l1i_pa [123]),
    .o(_al_u4447_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4448 (
    .a(_al_u4447_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[59]),
    .o(_al_u4448_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4449 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [59]),
    .d(addr_ex[59]),
    .o(_al_u4449_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4450 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [123]),
    .d(\biu/cache_ctrl_logic/pa_temp [123]),
    .o(_al_u4450_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4451 (
    .a(_al_u4448_o),
    .b(_al_u4449_o),
    .c(_al_u4450_o),
    .o(_al_u4451_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4452 (
    .a(_al_u4451_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [59]),
    .o(\biu/maddress [59]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4453 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [122]),
    .d(\biu/cache_ctrl_logic/pa_temp [122]),
    .o(_al_u4453_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4454 (
    .a(_al_u4453_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[58]),
    .o(_al_u4454_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4455 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [58]),
    .d(\biu/cache_ctrl_logic/l1i_pa [122]),
    .o(_al_u4455_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4456 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/n212 [58]),
    .d(addr_ex[58]),
    .o(_al_u4456_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4457 (
    .a(_al_u4454_o),
    .b(_al_u4455_o),
    .c(_al_u4456_o),
    .o(_al_u4457_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4458 (
    .a(_al_u4457_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [58]),
    .o(\biu/maddress [58]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4459 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [57]),
    .d(\biu/cache_ctrl_logic/l1i_pa [121]),
    .o(_al_u4459_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4460 (
    .a(_al_u4459_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[57]),
    .o(_al_u4460_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4461 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [57]),
    .d(addr_ex[57]),
    .o(_al_u4461_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4462 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [121]),
    .d(\biu/cache_ctrl_logic/pa_temp [121]),
    .o(_al_u4462_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4463 (
    .a(_al_u4460_o),
    .b(_al_u4461_o),
    .c(_al_u4462_o),
    .o(_al_u4463_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4464 (
    .a(_al_u4463_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [57]),
    .o(\biu/maddress [57]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4465 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [56]),
    .d(addr_ex[56]),
    .o(_al_u4465_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4466 (
    .a(_al_u4465_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[56]),
    .o(_al_u4466_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4467 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [56]),
    .d(\biu/cache_ctrl_logic/l1i_pa [120]),
    .o(_al_u4467_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4468 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [120]),
    .d(\biu/cache_ctrl_logic/pa_temp [120]),
    .o(_al_u4468_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4469 (
    .a(_al_u4466_o),
    .b(_al_u4467_o),
    .c(_al_u4468_o),
    .o(_al_u4469_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4470 (
    .a(_al_u4469_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [56]),
    .o(\biu/maddress [56]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4471 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [119]),
    .d(\biu/cache_ctrl_logic/pa_temp [119]),
    .o(_al_u4471_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4472 (
    .a(_al_u4471_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[55]),
    .o(_al_u4472_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4473 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [55]),
    .d(\biu/cache_ctrl_logic/l1i_pa [119]),
    .o(_al_u4473_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4474 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/n212 [55]),
    .d(addr_ex[55]),
    .o(_al_u4474_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4475 (
    .a(_al_u4472_o),
    .b(_al_u4473_o),
    .c(_al_u4474_o),
    .o(_al_u4475_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4476 (
    .a(_al_u4475_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [55]),
    .o(\biu/maddress [55]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4477 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [118]),
    .d(\biu/cache_ctrl_logic/pa_temp [118]),
    .o(_al_u4477_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4478 (
    .a(_al_u4477_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[54]),
    .o(_al_u4478_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4479 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [118]),
    .d(addr_ex[54]),
    .o(_al_u4479_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4480 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [54]),
    .d(\biu/cache_ctrl_logic/n212 [54]),
    .o(_al_u4480_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4481 (
    .a(_al_u4478_o),
    .b(_al_u4479_o),
    .c(_al_u4480_o),
    .o(_al_u4481_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4482 (
    .a(_al_u4481_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [54]),
    .o(\biu/maddress [54]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4483 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [53]),
    .d(\biu/cache_ctrl_logic/n212 [53]),
    .o(_al_u4483_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4484 (
    .a(_al_u4483_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[53]),
    .o(_al_u4484_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4485 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [117]),
    .d(addr_ex[53]),
    .o(_al_u4485_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4486 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [117]),
    .d(\biu/cache_ctrl_logic/pa_temp [117]),
    .o(_al_u4486_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4487 (
    .a(_al_u4484_o),
    .b(_al_u4485_o),
    .c(_al_u4486_o),
    .o(_al_u4487_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4488 (
    .a(_al_u4487_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [53]),
    .o(\biu/maddress [53]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4489 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [52]),
    .d(addr_ex[52]),
    .o(_al_u4489_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4490 (
    .a(_al_u4489_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[52]),
    .o(_al_u4490_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4491 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/n212 [52]),
    .d(\biu/cache_ctrl_logic/l1d_pa [116]),
    .o(_al_u4491_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4492 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [116]),
    .d(\biu/cache_ctrl_logic/pa_temp [116]),
    .o(_al_u4492_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4493 (
    .a(_al_u4490_o),
    .b(_al_u4491_o),
    .c(_al_u4492_o),
    .o(_al_u4493_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4494 (
    .a(_al_u4493_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [52]),
    .o(\biu/maddress [52]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4495 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [115]),
    .d(\biu/cache_ctrl_logic/pa_temp [115]),
    .o(_al_u4495_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4496 (
    .a(_al_u4495_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[51]),
    .o(_al_u4496_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4497 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [51]),
    .d(\biu/cache_ctrl_logic/l1i_pa [115]),
    .o(_al_u4497_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4498 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/n212 [51]),
    .d(addr_ex[51]),
    .o(_al_u4498_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4499 (
    .a(_al_u4496_o),
    .b(_al_u4497_o),
    .c(_al_u4498_o),
    .o(_al_u4499_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4500 (
    .a(_al_u4499_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [51]),
    .o(\biu/maddress [51]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4501 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [50]),
    .d(\biu/cache_ctrl_logic/l1i_pa [114]),
    .o(_al_u4501_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4502 (
    .a(_al_u4501_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[50]),
    .o(_al_u4502_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4503 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [50]),
    .d(\biu/cache_ctrl_logic/l1d_pa [114]),
    .o(_al_u4503_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4504 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [114]),
    .d(addr_ex[50]),
    .o(_al_u4504_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4505 (
    .a(_al_u4502_o),
    .b(_al_u4503_o),
    .c(_al_u4504_o),
    .o(_al_u4505_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4506 (
    .a(_al_u4505_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [50]),
    .o(\biu/maddress [50]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4507 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [5]),
    .d(\biu/cache_ctrl_logic/n212 [5]),
    .o(_al_u4507_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4508 (
    .a(_al_u4507_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[5]),
    .o(_al_u4508_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4509 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [69]),
    .d(addr_ex[5]),
    .o(_al_u4509_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4510 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [69]),
    .d(\biu/cache_ctrl_logic/pa_temp [69]),
    .o(_al_u4510_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4511 (
    .a(_al_u4508_o),
    .b(_al_u4509_o),
    .c(_al_u4510_o),
    .o(_al_u4511_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4512 (
    .a(_al_u4511_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [5]),
    .o(\biu/maddress [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4513 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [113]),
    .d(\biu/cache_ctrl_logic/pa_temp [113]),
    .o(_al_u4513_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4514 (
    .a(_al_u4513_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[49]),
    .o(_al_u4514_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4515 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [49]),
    .d(\biu/cache_ctrl_logic/l1i_pa [113]),
    .o(_al_u4515_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4516 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/n212 [49]),
    .d(addr_ex[49]),
    .o(_al_u4516_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4517 (
    .a(_al_u4514_o),
    .b(_al_u4515_o),
    .c(_al_u4516_o),
    .o(_al_u4517_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4518 (
    .a(_al_u4517_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [49]),
    .o(\biu/maddress [49]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4519 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [112]),
    .d(\biu/cache_ctrl_logic/pa_temp [112]),
    .o(_al_u4519_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4520 (
    .a(_al_u4519_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[48]),
    .o(_al_u4520_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4521 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [112]),
    .d(addr_ex[48]),
    .o(_al_u4521_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4522 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [48]),
    .d(\biu/cache_ctrl_logic/n212 [48]),
    .o(_al_u4522_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4523 (
    .a(_al_u4520_o),
    .b(_al_u4521_o),
    .c(_al_u4522_o),
    .o(_al_u4523_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4524 (
    .a(_al_u4523_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [48]),
    .o(\biu/maddress [48]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4525 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [111]),
    .d(\biu/cache_ctrl_logic/pa_temp [111]),
    .o(_al_u4525_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4526 (
    .a(_al_u4525_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[47]),
    .o(_al_u4526_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4527 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [47]),
    .d(\biu/cache_ctrl_logic/l1i_pa [111]),
    .o(_al_u4527_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4528 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/n212 [47]),
    .d(addr_ex[47]),
    .o(_al_u4528_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4529 (
    .a(_al_u4526_o),
    .b(_al_u4527_o),
    .c(_al_u4528_o),
    .o(_al_u4529_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4530 (
    .a(_al_u4529_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [47]),
    .o(\biu/maddress [47]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4531 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [46]),
    .d(\biu/cache_ctrl_logic/l1i_pa [110]),
    .o(_al_u4531_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4532 (
    .a(_al_u4531_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[46]),
    .o(_al_u4532_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4533 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/n212 [46]),
    .d(addr_ex[46]),
    .o(_al_u4533_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4534 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [110]),
    .d(\biu/cache_ctrl_logic/pa_temp [110]),
    .o(_al_u4534_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4535 (
    .a(_al_u4532_o),
    .b(_al_u4533_o),
    .c(_al_u4534_o),
    .o(_al_u4535_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4536 (
    .a(_al_u4535_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [46]),
    .o(\biu/maddress [46]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4537 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [45]),
    .d(\biu/cache_ctrl_logic/l1i_pa [109]),
    .o(_al_u4537_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4538 (
    .a(_al_u4537_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[45]),
    .o(_al_u4538_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4539 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [45]),
    .d(\biu/cache_ctrl_logic/l1d_pa [109]),
    .o(_al_u4539_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4540 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [109]),
    .d(addr_ex[45]),
    .o(_al_u4540_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4541 (
    .a(_al_u4538_o),
    .b(_al_u4539_o),
    .c(_al_u4540_o),
    .o(_al_u4541_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4542 (
    .a(_al_u4541_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [45]),
    .o(\biu/maddress [45]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4543 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [108]),
    .d(addr_ex[44]),
    .o(_al_u4543_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4544 (
    .a(_al_u4543_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[44]),
    .o(_al_u4544_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4545 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [44]),
    .d(\biu/cache_ctrl_logic/n212 [44]),
    .o(_al_u4545_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4546 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [108]),
    .d(\biu/cache_ctrl_logic/pa_temp [108]),
    .o(_al_u4546_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4547 (
    .a(_al_u4544_o),
    .b(_al_u4545_o),
    .c(_al_u4546_o),
    .o(_al_u4547_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4548 (
    .a(_al_u4547_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [44]),
    .o(\biu/maddress [44]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4549 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [107]),
    .d(addr_ex[43]),
    .o(_al_u4549_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4550 (
    .a(_al_u4549_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[43]),
    .o(_al_u4550_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4551 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [43]),
    .d(\biu/cache_ctrl_logic/n212 [43]),
    .o(_al_u4551_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4552 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [107]),
    .d(\biu/cache_ctrl_logic/pa_temp [107]),
    .o(_al_u4552_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4553 (
    .a(_al_u4550_o),
    .b(_al_u4551_o),
    .c(_al_u4552_o),
    .o(_al_u4553_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4554 (
    .a(_al_u4553_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [43]),
    .o(\biu/maddress [43]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4555 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [42]),
    .d(\biu/cache_ctrl_logic/n212 [42]),
    .o(_al_u4555_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4556 (
    .a(_al_u4555_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[42]),
    .o(_al_u4556_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4557 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [106]),
    .d(addr_ex[42]),
    .o(_al_u4557_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4558 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [106]),
    .d(\biu/cache_ctrl_logic/pa_temp [106]),
    .o(_al_u4558_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4559 (
    .a(_al_u4556_o),
    .b(_al_u4557_o),
    .c(_al_u4558_o),
    .o(_al_u4559_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4560 (
    .a(_al_u4559_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [42]),
    .o(\biu/maddress [42]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4561 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [41]),
    .d(\biu/cache_ctrl_logic/l1i_pa [105]),
    .o(_al_u4561_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4562 (
    .a(_al_u4561_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[41]),
    .o(_al_u4562_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4563 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [41]),
    .d(\biu/cache_ctrl_logic/l1d_pa [105]),
    .o(_al_u4563_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4564 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [105]),
    .d(addr_ex[41]),
    .o(_al_u4564_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4565 (
    .a(_al_u4562_o),
    .b(_al_u4563_o),
    .c(_al_u4564_o),
    .o(_al_u4565_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4566 (
    .a(_al_u4565_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [41]),
    .o(\biu/maddress [41]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4567 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [40]),
    .d(\biu/cache_ctrl_logic/l1i_pa [104]),
    .o(_al_u4567_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4568 (
    .a(_al_u4567_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[40]),
    .o(_al_u4568_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4569 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [40]),
    .d(\biu/cache_ctrl_logic/l1d_pa [104]),
    .o(_al_u4569_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4570 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [104]),
    .d(addr_ex[40]),
    .o(_al_u4570_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4571 (
    .a(_al_u4568_o),
    .b(_al_u4569_o),
    .c(_al_u4570_o),
    .o(_al_u4571_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4572 (
    .a(_al_u4571_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [40]),
    .o(\biu/maddress [40]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4573 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [4]),
    .d(addr_ex[4]),
    .o(_al_u4573_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4574 (
    .a(_al_u4573_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[4]),
    .o(_al_u4574_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4575 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/n212 [4]),
    .d(\biu/cache_ctrl_logic/l1d_pa [68]),
    .o(_al_u4575_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4576 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [68]),
    .d(\biu/cache_ctrl_logic/pa_temp [68]),
    .o(_al_u4576_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4577 (
    .a(_al_u4574_o),
    .b(_al_u4575_o),
    .c(_al_u4576_o),
    .o(_al_u4577_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4578 (
    .a(_al_u4577_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [4]),
    .o(\biu/maddress [4]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4579 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [103]),
    .d(\biu/cache_ctrl_logic/pa_temp [103]),
    .o(_al_u4579_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4580 (
    .a(_al_u4579_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[39]),
    .o(_al_u4580_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4581 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [39]),
    .d(\biu/cache_ctrl_logic/l1i_pa [103]),
    .o(_al_u4581_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4582 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/n212 [39]),
    .d(addr_ex[39]),
    .o(_al_u4582_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4583 (
    .a(_al_u4580_o),
    .b(_al_u4581_o),
    .c(_al_u4582_o),
    .o(_al_u4583_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4584 (
    .a(_al_u4583_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [39]),
    .o(\biu/maddress [39]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4585 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [102]),
    .d(\biu/cache_ctrl_logic/pa_temp [102]),
    .o(_al_u4585_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4586 (
    .a(_al_u4585_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[38]),
    .o(_al_u4586_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4587 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [38]),
    .d(\biu/cache_ctrl_logic/l1i_pa [102]),
    .o(_al_u4587_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4588 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [38]),
    .d(addr_ex[38]),
    .o(_al_u4588_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4589 (
    .a(_al_u4586_o),
    .b(_al_u4587_o),
    .c(_al_u4588_o),
    .o(_al_u4589_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4590 (
    .a(_al_u4589_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [38]),
    .o(\biu/maddress [38]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4591 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [37]),
    .d(\biu/cache_ctrl_logic/l1i_pa [101]),
    .o(_al_u4591_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4592 (
    .a(_al_u4591_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[37]),
    .o(_al_u4592_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4593 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [37]),
    .d(\biu/cache_ctrl_logic/l1d_pa [101]),
    .o(_al_u4593_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4594 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [101]),
    .d(addr_ex[37]),
    .o(_al_u4594_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4595 (
    .a(_al_u4592_o),
    .b(_al_u4593_o),
    .c(_al_u4594_o),
    .o(_al_u4595_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4596 (
    .a(_al_u4595_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [37]),
    .o(\biu/maddress [37]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4597 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [36]),
    .d(addr_ex[36]),
    .o(_al_u4597_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4598 (
    .a(_al_u4597_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[36]),
    .o(_al_u4598_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4599 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/n212 [36]),
    .d(\biu/cache_ctrl_logic/l1d_pa [100]),
    .o(_al_u4599_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4600 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [100]),
    .d(\biu/cache_ctrl_logic/pa_temp [100]),
    .o(_al_u4600_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4601 (
    .a(_al_u4598_o),
    .b(_al_u4599_o),
    .c(_al_u4600_o),
    .o(_al_u4601_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4602 (
    .a(_al_u4601_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [36]),
    .o(\biu/maddress [36]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4603 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [35]),
    .d(addr_ex[35]),
    .o(_al_u4603_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4604 (
    .a(_al_u4603_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[35]),
    .o(_al_u4604_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4605 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [35]),
    .d(\biu/cache_ctrl_logic/l1i_pa [99]),
    .o(_al_u4605_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4606 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [99]),
    .d(\biu/cache_ctrl_logic/pa_temp [99]),
    .o(_al_u4606_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4607 (
    .a(_al_u4604_o),
    .b(_al_u4605_o),
    .c(_al_u4606_o),
    .o(_al_u4607_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4608 (
    .a(_al_u4607_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [35]),
    .o(\biu/maddress [35]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4609 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [98]),
    .d(\biu/cache_ctrl_logic/pa_temp [98]),
    .o(_al_u4609_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4610 (
    .a(_al_u4609_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[34]),
    .o(_al_u4610_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4611 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [98]),
    .d(addr_ex[34]),
    .o(_al_u4611_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4612 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [34]),
    .d(\biu/cache_ctrl_logic/n212 [34]),
    .o(_al_u4612_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4613 (
    .a(_al_u4610_o),
    .b(_al_u4611_o),
    .c(_al_u4612_o),
    .o(_al_u4613_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4614 (
    .a(_al_u4613_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [34]),
    .o(\biu/maddress [34]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4615 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [33]),
    .d(\biu/cache_ctrl_logic/n212 [33]),
    .o(_al_u4615_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4616 (
    .a(_al_u4615_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[33]),
    .o(_al_u4616_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4617 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [97]),
    .d(addr_ex[33]),
    .o(_al_u4617_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4618 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [97]),
    .d(\biu/cache_ctrl_logic/pa_temp [97]),
    .o(_al_u4618_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4619 (
    .a(_al_u4616_o),
    .b(_al_u4617_o),
    .c(_al_u4618_o),
    .o(_al_u4619_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4620 (
    .a(_al_u4619_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [33]),
    .o(\biu/maddress [33]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4621 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [32]),
    .d(addr_ex[32]),
    .o(_al_u4621_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4622 (
    .a(_al_u4621_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[32]),
    .o(_al_u4622_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4623 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/n212 [32]),
    .d(\biu/cache_ctrl_logic/l1d_pa [96]),
    .o(_al_u4623_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4624 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [96]),
    .d(\biu/cache_ctrl_logic/pa_temp [96]),
    .o(_al_u4624_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4625 (
    .a(_al_u4622_o),
    .b(_al_u4623_o),
    .c(_al_u4624_o),
    .o(_al_u4625_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4626 (
    .a(_al_u4625_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [32]),
    .o(\biu/maddress [32]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4627 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [95]),
    .d(\biu/cache_ctrl_logic/pa_temp [95]),
    .o(_al_u4627_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4628 (
    .a(_al_u4627_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[31]),
    .o(_al_u4628_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4629 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [31]),
    .d(\biu/cache_ctrl_logic/l1i_pa [95]),
    .o(_al_u4629_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4630 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/n212 [31]),
    .d(addr_ex[31]),
    .o(_al_u4630_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4631 (
    .a(_al_u4628_o),
    .b(_al_u4629_o),
    .c(_al_u4630_o),
    .o(_al_u4631_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4632 (
    .a(_al_u4631_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [31]),
    .o(\biu/maddress [31]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4633 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [30]),
    .d(addr_ex[30]),
    .o(_al_u4633_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4634 (
    .a(_al_u4633_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[30]),
    .o(_al_u4634_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4635 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/n212 [30]),
    .d(\biu/cache_ctrl_logic/l1d_pa [94]),
    .o(_al_u4635_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4636 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [94]),
    .d(\biu/cache_ctrl_logic/pa_temp [94]),
    .o(_al_u4636_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4637 (
    .a(_al_u4634_o),
    .b(_al_u4635_o),
    .c(_al_u4636_o),
    .o(_al_u4637_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4638 (
    .a(_al_u4637_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [30]),
    .o(\biu/maddress [30]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4639 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [3]),
    .d(\biu/cache_ctrl_logic/n212 [3]),
    .o(_al_u4639_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4640 (
    .a(_al_u4639_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[3]),
    .o(_al_u4640_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4641 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [67]),
    .d(addr_ex[3]),
    .o(_al_u4641_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4642 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [67]),
    .d(\biu/cache_ctrl_logic/pa_temp [67]),
    .o(_al_u4642_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4643 (
    .a(_al_u4640_o),
    .b(_al_u4641_o),
    .c(_al_u4642_o),
    .o(_al_u4643_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4644 (
    .a(_al_u4643_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [3]),
    .o(\biu/maddress [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4645 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [29]),
    .d(\biu/cache_ctrl_logic/n212 [29]),
    .o(_al_u4645_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4646 (
    .a(_al_u4645_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[29]),
    .o(_al_u4646_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4647 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [93]),
    .d(addr_ex[29]),
    .o(_al_u4647_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4648 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [93]),
    .d(\biu/cache_ctrl_logic/pa_temp [93]),
    .o(_al_u4648_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4649 (
    .a(_al_u4646_o),
    .b(_al_u4647_o),
    .c(_al_u4648_o),
    .o(_al_u4649_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4650 (
    .a(_al_u4649_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [29]),
    .o(\biu/maddress [29]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4651 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [28]),
    .d(\biu/cache_ctrl_logic/n212 [28]),
    .o(_al_u4651_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4652 (
    .a(_al_u4651_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[28]),
    .o(_al_u4652_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4653 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [92]),
    .d(addr_ex[28]),
    .o(_al_u4653_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4654 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [92]),
    .d(\biu/cache_ctrl_logic/pa_temp [92]),
    .o(_al_u4654_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4655 (
    .a(_al_u4652_o),
    .b(_al_u4653_o),
    .c(_al_u4654_o),
    .o(_al_u4655_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4656 (
    .a(_al_u4655_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [28]),
    .o(\biu/maddress [28]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4657 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [27]),
    .d(addr_ex[27]),
    .o(_al_u4657_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4658 (
    .a(_al_u4657_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[27]),
    .o(_al_u4658_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4659 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [27]),
    .d(\biu/cache_ctrl_logic/l1i_pa [91]),
    .o(_al_u4659_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4660 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [91]),
    .d(\biu/cache_ctrl_logic/pa_temp [91]),
    .o(_al_u4660_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4661 (
    .a(_al_u4658_o),
    .b(_al_u4659_o),
    .c(_al_u4660_o),
    .o(_al_u4661_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4662 (
    .a(_al_u4661_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [27]),
    .o(\biu/maddress [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4663 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [90]),
    .d(\biu/cache_ctrl_logic/pa_temp [90]),
    .o(_al_u4663_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4664 (
    .a(_al_u4663_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[26]),
    .o(_al_u4664_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4665 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [26]),
    .d(\biu/cache_ctrl_logic/l1i_pa [90]),
    .o(_al_u4665_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4666 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/n212 [26]),
    .d(addr_ex[26]),
    .o(_al_u4666_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4667 (
    .a(_al_u4664_o),
    .b(_al_u4665_o),
    .c(_al_u4666_o),
    .o(_al_u4667_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4668 (
    .a(_al_u4667_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [26]),
    .o(\biu/maddress [26]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4669 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [89]),
    .d(\biu/cache_ctrl_logic/pa_temp [89]),
    .o(_al_u4669_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4670 (
    .a(_al_u4669_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[25]),
    .o(_al_u4670_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4671 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [89]),
    .d(addr_ex[25]),
    .o(_al_u4671_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4672 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [25]),
    .d(\biu/cache_ctrl_logic/n212 [25]),
    .o(_al_u4672_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4673 (
    .a(_al_u4670_o),
    .b(_al_u4671_o),
    .c(_al_u4672_o),
    .o(_al_u4673_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4674 (
    .a(_al_u4673_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [25]),
    .o(\biu/maddress [25]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4675 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [24]),
    .d(\biu/cache_ctrl_logic/l1i_pa [88]),
    .o(_al_u4675_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4676 (
    .a(_al_u4675_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[24]),
    .o(_al_u4676_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4677 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [24]),
    .d(\biu/cache_ctrl_logic/l1d_pa [88]),
    .o(_al_u4677_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4678 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [88]),
    .d(addr_ex[24]),
    .o(_al_u4678_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4679 (
    .a(_al_u4676_o),
    .b(_al_u4677_o),
    .c(_al_u4678_o),
    .o(_al_u4679_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4680 (
    .a(_al_u4679_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [24]),
    .o(\biu/maddress [24]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4681 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [87]),
    .d(addr_ex[23]),
    .o(_al_u4681_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4682 (
    .a(_al_u4681_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[23]),
    .o(_al_u4682_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4683 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [23]),
    .d(\biu/cache_ctrl_logic/n212 [23]),
    .o(_al_u4683_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4684 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [87]),
    .d(\biu/cache_ctrl_logic/pa_temp [87]),
    .o(_al_u4684_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4685 (
    .a(_al_u4682_o),
    .b(_al_u4683_o),
    .c(_al_u4684_o),
    .o(_al_u4685_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4686 (
    .a(_al_u4685_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [23]),
    .o(\biu/maddress [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4687 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [22]),
    .d(\biu/cache_ctrl_logic/l1i_pa [86]),
    .o(_al_u4687_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4688 (
    .a(_al_u4687_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[22]),
    .o(_al_u4688_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4689 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [22]),
    .d(addr_ex[22]),
    .o(_al_u4689_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4690 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [86]),
    .d(\biu/cache_ctrl_logic/pa_temp [86]),
    .o(_al_u4690_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4691 (
    .a(_al_u4688_o),
    .b(_al_u4689_o),
    .c(_al_u4690_o),
    .o(_al_u4691_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4692 (
    .a(_al_u4691_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [22]),
    .o(\biu/maddress [22]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4693 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [21]),
    .d(\biu/cache_ctrl_logic/l1i_pa [85]),
    .o(_al_u4693_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4694 (
    .a(_al_u4693_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[21]),
    .o(_al_u4694_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4695 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [21]),
    .d(\biu/cache_ctrl_logic/l1d_pa [85]),
    .o(_al_u4695_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4696 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [85]),
    .d(addr_ex[21]),
    .o(_al_u4696_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4697 (
    .a(_al_u4694_o),
    .b(_al_u4695_o),
    .c(_al_u4696_o),
    .o(_al_u4697_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4698 (
    .a(_al_u4697_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [21]),
    .o(\biu/maddress [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4699 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [20]),
    .d(\biu/cache_ctrl_logic/l1i_pa [84]),
    .o(_al_u4699_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4700 (
    .a(_al_u4699_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[20]),
    .o(_al_u4700_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4701 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [20]),
    .d(addr_ex[20]),
    .o(_al_u4701_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4702 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [84]),
    .d(\biu/cache_ctrl_logic/pa_temp [84]),
    .o(_al_u4702_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4703 (
    .a(_al_u4700_o),
    .b(_al_u4701_o),
    .c(_al_u4702_o),
    .o(_al_u4703_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4704 (
    .a(_al_u4703_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [20]),
    .o(\biu/maddress [20]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4705 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [19]),
    .d(addr_ex[19]),
    .o(_al_u4705_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4706 (
    .a(_al_u4705_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[19]),
    .o(_al_u4706_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4707 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/n212 [19]),
    .d(\biu/cache_ctrl_logic/l1d_pa [83]),
    .o(_al_u4707_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4708 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [83]),
    .d(\biu/cache_ctrl_logic/pa_temp [83]),
    .o(_al_u4708_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4709 (
    .a(_al_u4706_o),
    .b(_al_u4707_o),
    .c(_al_u4708_o),
    .o(_al_u4709_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4710 (
    .a(_al_u4709_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [19]),
    .o(\biu/maddress [19]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4711 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [82]),
    .d(addr_ex[18]),
    .o(_al_u4711_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4712 (
    .a(_al_u4711_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[18]),
    .o(_al_u4712_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4713 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [18]),
    .d(\biu/cache_ctrl_logic/n212 [18]),
    .o(_al_u4713_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4714 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [82]),
    .d(\biu/cache_ctrl_logic/pa_temp [82]),
    .o(_al_u4714_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4715 (
    .a(_al_u4712_o),
    .b(_al_u4713_o),
    .c(_al_u4714_o),
    .o(_al_u4715_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4716 (
    .a(_al_u4715_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [18]),
    .o(\biu/maddress [18]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4717 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [17]),
    .d(\biu/cache_ctrl_logic/l1i_pa [81]),
    .o(_al_u4717_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4718 (
    .a(_al_u4717_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[17]),
    .o(_al_u4718_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4719 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [17]),
    .d(\biu/cache_ctrl_logic/l1d_pa [81]),
    .o(_al_u4719_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4720 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [81]),
    .d(addr_ex[17]),
    .o(_al_u4720_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4721 (
    .a(_al_u4718_o),
    .b(_al_u4719_o),
    .c(_al_u4720_o),
    .o(_al_u4721_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4722 (
    .a(_al_u4721_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [17]),
    .o(\biu/maddress [17]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4723 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [16]),
    .d(\biu/cache_ctrl_logic/l1i_pa [80]),
    .o(_al_u4723_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4724 (
    .a(_al_u4723_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[16]),
    .o(_al_u4724_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4725 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [16]),
    .d(\biu/cache_ctrl_logic/l1d_pa [80]),
    .o(_al_u4725_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4726 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [80]),
    .d(addr_ex[16]),
    .o(_al_u4726_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4727 (
    .a(_al_u4724_o),
    .b(_al_u4725_o),
    .c(_al_u4726_o),
    .o(_al_u4727_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4728 (
    .a(_al_u4727_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [16]),
    .o(\biu/maddress [16]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4729 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [79]),
    .d(\biu/cache_ctrl_logic/pa_temp [79]),
    .o(_al_u4729_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4730 (
    .a(_al_u4729_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[15]),
    .o(_al_u4730_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4731 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [15]),
    .d(\biu/cache_ctrl_logic/l1i_pa [79]),
    .o(_al_u4731_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4732 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/n212 [15]),
    .d(addr_ex[15]),
    .o(_al_u4732_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4733 (
    .a(_al_u4730_o),
    .b(_al_u4731_o),
    .c(_al_u4732_o),
    .o(_al_u4733_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4734 (
    .a(_al_u4733_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [15]),
    .o(\biu/maddress [15]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4735 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [78]),
    .d(\biu/cache_ctrl_logic/pa_temp [78]),
    .o(_al_u4735_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4736 (
    .a(_al_u4735_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[14]),
    .o(_al_u4736_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4737 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [14]),
    .d(\biu/cache_ctrl_logic/l1i_pa [78]),
    .o(_al_u4737_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4738 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [14]),
    .d(addr_ex[14]),
    .o(_al_u4738_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4739 (
    .a(_al_u4736_o),
    .b(_al_u4737_o),
    .c(_al_u4738_o),
    .o(_al_u4739_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4740 (
    .a(_al_u4739_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [14]),
    .o(\biu/maddress [14]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4741 (
    .a(_al_u3950_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [13]),
    .d(\biu/cache_ctrl_logic/l1i_pa [77]),
    .o(_al_u4741_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4742 (
    .a(_al_u4741_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[13]),
    .o(_al_u4742_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4743 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [77]),
    .d(addr_ex[13]),
    .o(_al_u4743_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4744 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/n212 [13]),
    .d(\biu/cache_ctrl_logic/pa_temp [77]),
    .o(_al_u4744_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4745 (
    .a(_al_u4742_o),
    .b(_al_u4743_o),
    .c(_al_u4744_o),
    .o(_al_u4745_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4746 (
    .a(_al_u4745_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [13]),
    .o(\biu/maddress [13]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4747 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [12]),
    .d(\biu/cache_ctrl_logic/n212 [12]),
    .o(_al_u4747_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4748 (
    .a(_al_u4747_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[12]),
    .o(_al_u4748_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4749 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [76]),
    .d(addr_ex[12]),
    .o(_al_u4749_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4750 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [76]),
    .d(\biu/cache_ctrl_logic/pa_temp [76]),
    .o(_al_u4750_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4751 (
    .a(_al_u4748_o),
    .b(_al_u4749_o),
    .c(_al_u4750_o),
    .o(_al_u4751_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4752 (
    .a(_al_u4751_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [12]),
    .o(\biu/maddress [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4753 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/n212 [11]),
    .d(\biu/cache_ctrl_logic/l1i_pa [75]),
    .o(_al_u4753_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4754 (
    .a(_al_u4753_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[11]),
    .o(_al_u4754_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4755 (
    .a(_al_u3947_o),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [11]),
    .d(\biu/cache_ctrl_logic/l1d_pa [75]),
    .o(_al_u4755_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4756 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/pa_temp [75]),
    .d(addr_ex[11]),
    .o(_al_u4756_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4757 (
    .a(_al_u4754_o),
    .b(_al_u4755_o),
    .c(_al_u4756_o),
    .o(_al_u4757_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4758 (
    .a(_al_u4757_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [11]),
    .o(\biu/maddress [11]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4759 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [74]),
    .d(\biu/cache_ctrl_logic/pa_temp [74]),
    .o(_al_u4759_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4760 (
    .a(_al_u4759_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .c(addr_if[10]),
    .o(_al_u4760_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4761 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [74]),
    .d(addr_ex[10]),
    .o(_al_u4761_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4762 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [10]),
    .d(\biu/cache_ctrl_logic/n212 [10]),
    .o(_al_u4762_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u4763 (
    .a(_al_u4760_o),
    .b(_al_u4761_o),
    .c(_al_u4762_o),
    .o(_al_u4763_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u4764 (
    .a(_al_u4763_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [10]),
    .o(\biu/maddress [10]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4765 (
    .a(hresp_pad),
    .b(\biu/bus_unit/mux11_b4_sel_is_2_o ),
    .o(_al_u4765_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C)*~(A)+~(D*~B)*C*~(A)+~(~(D*~B))*C*A+~(D*~B)*C*A)"),
    .INIT(16'he4f5))
    _al_u4766 (
    .a(_al_u3404_o),
    .b(_al_u3407_o),
    .c(_al_u4099_o),
    .d(\biu/bus_unit/statu [2]),
    .o(_al_u4766_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u4767 (
    .a(_al_u4765_o),
    .b(_al_u4766_o),
    .o(\biu/bus_unit/n35 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4768 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [7]),
    .d(\biu/cache_ctrl_logic/pte_temp [7]),
    .o(_al_u4768_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4769 (
    .a(_al_u2705_o),
    .b(_al_u4768_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [7]),
    .o(_al_u4769_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4770 (
    .a(\exu/lsu/n1 [7]),
    .b(_al_u4769_o),
    .c(_al_u3222_o),
    .o(_al_u4770_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4771 (
    .a(_al_u4770_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [7]),
    .o(hwdata_pad[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4772 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [6]),
    .d(\biu/cache_ctrl_logic/l1d_pte [6]),
    .o(_al_u4772_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4773 (
    .a(_al_u2705_o),
    .b(_al_u4772_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [6]),
    .o(_al_u4773_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4774 (
    .a(\exu/lsu/n1 [6]),
    .b(_al_u4773_o),
    .c(_al_u3222_o),
    .o(_al_u4774_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4775 (
    .a(_al_u4774_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [6]),
    .o(hwdata_pad[6]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4776 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [5]),
    .d(\biu/cache_ctrl_logic/l1d_pte [5]),
    .o(_al_u4776_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4777 (
    .a(_al_u2705_o),
    .b(_al_u4776_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [5]),
    .o(_al_u4777_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4778 (
    .a(\exu/lsu/n1 [5]),
    .b(_al_u4777_o),
    .c(_al_u3222_o),
    .o(_al_u4778_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4779 (
    .a(_al_u4778_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [5]),
    .o(hwdata_pad[5]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4780 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [4]),
    .d(\biu/cache_ctrl_logic/l1d_pte [4]),
    .o(_al_u4780_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4781 (
    .a(_al_u2705_o),
    .b(_al_u4780_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [4]),
    .o(_al_u4781_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4782 (
    .a(\exu/lsu/n1 [4]),
    .b(_al_u4781_o),
    .c(_al_u3222_o),
    .o(_al_u4782_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4783 (
    .a(_al_u4782_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [4]),
    .o(hwdata_pad[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4784 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [3]),
    .d(\biu/cache_ctrl_logic/l1d_pte [3]),
    .o(_al_u4784_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4785 (
    .a(_al_u2705_o),
    .b(_al_u4784_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [3]),
    .o(_al_u4785_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4786 (
    .a(\exu/lsu/n1 [3]),
    .b(_al_u4785_o),
    .c(_al_u3222_o),
    .o(_al_u4786_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4787 (
    .a(_al_u4786_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [3]),
    .o(hwdata_pad[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4788 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [2]),
    .d(\biu/cache_ctrl_logic/l1d_pte [2]),
    .o(_al_u4788_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4789 (
    .a(_al_u2705_o),
    .b(_al_u4788_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [2]),
    .o(_al_u4789_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4790 (
    .a(\exu/lsu/n1 [2]),
    .b(_al_u4789_o),
    .c(_al_u3222_o),
    .o(_al_u4790_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4791 (
    .a(_al_u4790_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [2]),
    .o(hwdata_pad[2]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4792 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [1]),
    .d(\biu/cache_ctrl_logic/l1d_pte [1]),
    .o(_al_u4792_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4793 (
    .a(_al_u2705_o),
    .b(_al_u4792_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [1]),
    .o(_al_u4793_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4794 (
    .a(\exu/lsu/n1 [1]),
    .b(_al_u4793_o),
    .c(_al_u3222_o),
    .o(_al_u4794_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4795 (
    .a(_al_u4794_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [1]),
    .o(hwdata_pad[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4796 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [0]),
    .d(\biu/cache_ctrl_logic/pte_temp [0]),
    .o(_al_u4796_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4797 (
    .a(_al_u4796_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [0]),
    .o(_al_u4797_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4798 (
    .a(\exu/lsu/n1 [0]),
    .b(_al_u4797_o),
    .c(_al_u3222_o),
    .o(_al_u4798_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u4799 (
    .a(_al_u4798_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [0]),
    .o(hwdata_pad[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u4800 (
    .a(_al_u4092_o),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .d(_al_u3384_o),
    .o(\ins_dec/ins_srli ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u4801 (
    .a(_al_u3925_o),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .d(_al_u3384_o),
    .o(_al_u4801_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(~C*~B)))"),
    .INIT(16'h0155))
    _al_u4802 (
    .a(\ins_dec/ins_srli ),
    .b(\ins_dec/funct7_0_lutinv ),
    .c(\ins_dec/funct7_32_lutinv ),
    .d(_al_u4801_o),
    .o(_al_u4802_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u4803 (
    .a(\ins_dec/op_32_imm_lutinv ),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .d(_al_u3384_o),
    .o(\ins_dec/n38 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u4804 (
    .a(id_ins[26]),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .d(_al_u3384_o),
    .o(_al_u4804_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u4805 (
    .a(\ins_dec/funct5_8_lutinv ),
    .b(_al_u3927_o),
    .c(_al_u4804_o),
    .d(_al_u3928_o),
    .o(\ins_dec/ins_srai ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u4806 (
    .a(\ins_dec/n38 ),
    .b(\ins_dec/ins_srai ),
    .c(\ins_dec/funct7_32_lutinv ),
    .o(_al_u4806_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u4807 (
    .a(_al_u4802_o),
    .b(_al_u4806_o),
    .c(\ins_dec/funct7_0_lutinv ),
    .d(\ins_dec/n38 ),
    .o(\ins_dec/n232 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4808 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [2]),
    .d(\biu/cache_ctrl_logic/n212 [2]),
    .o(_al_u4808_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4809 (
    .a(_al_u4808_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [66]),
    .o(_al_u4809_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4810 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [66]),
    .d(\biu/cache_ctrl_logic/pa_temp [66]),
    .o(_al_u4810_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4811 (
    .a(_al_u2705_o),
    .b(_al_u4810_o),
    .c(\biu/cache_ctrl_logic/n75_lutinv ),
    .d(addr_ex[2]),
    .o(_al_u4811_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u4812 (
    .a(_al_u4809_o),
    .b(_al_u4811_o),
    .c(\biu/bus_unit/mmu/n19_lutinv ),
    .d(addr_if[2]),
    .o(_al_u4812_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4813 (
    .a(_al_u4812_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [2]),
    .o(_al_u4813_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4814 (
    .a(_al_u4813_o),
    .b(_al_u2705_o),
    .c(\biu/paddress [66]),
    .o(haddr_pad[2]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4815 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [1]),
    .d(addr_ex[1]),
    .o(_al_u4815_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4816 (
    .a(_al_u4815_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [65]),
    .o(_al_u4816_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4817 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pa [65]),
    .d(\biu/cache_ctrl_logic/pa_temp [65]),
    .o(_al_u4817_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4818 (
    .a(_al_u2705_o),
    .b(_al_u4817_o),
    .c(\biu/cache_ctrl_logic/n97_lutinv ),
    .d(\biu/cache_ctrl_logic/n212 [1]),
    .o(_al_u4818_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u4819 (
    .a(_al_u4816_o),
    .b(_al_u4818_o),
    .c(\biu/bus_unit/mmu/n19_lutinv ),
    .d(addr_if[1]),
    .o(_al_u4819_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4820 (
    .a(_al_u4819_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [1]),
    .o(_al_u4820_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4821 (
    .a(_al_u4820_o),
    .b(_al_u2705_o),
    .c(\biu/paddress [65]),
    .o(haddr_pad[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4822 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n209 [0]),
    .d(addr_ex[0]),
    .o(_al_u4822_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u4823 (
    .a(_al_u4822_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pa [64]),
    .o(_al_u4823_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u4824 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u3945_o),
    .c(\biu/cache_ctrl_logic/n212 [0]),
    .d(\biu/cache_ctrl_logic/pa_temp [64]),
    .o(_al_u4824_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4825 (
    .a(_al_u2705_o),
    .b(_al_u4824_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pa [64]),
    .o(_al_u4825_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u4826 (
    .a(_al_u4823_o),
    .b(_al_u4825_o),
    .c(\biu/bus_unit/mmu/n19_lutinv ),
    .d(addr_if[0]),
    .o(_al_u4826_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u4827 (
    .a(_al_u4826_o),
    .b(_al_u4403_o),
    .c(\biu/cache_ctrl_logic/n207 [0]),
    .o(_al_u4827_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4828 (
    .a(_al_u4827_o),
    .b(_al_u2705_o),
    .c(\biu/paddress [64]),
    .o(haddr_pad[0]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u4829 (
    .a(_al_u2890_o),
    .b(_al_u3404_o),
    .c(_al_u4099_o),
    .o(_al_u4829_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~C*~B))"),
    .INIT(16'ha8aa))
    _al_u4830 (
    .a(_al_u4829_o),
    .b(_al_u2890_o),
    .c(_al_u3407_o),
    .d(\biu/bus_unit/statu [1]),
    .o(_al_u4830_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u4831 (
    .a(_al_u4830_o),
    .b(_al_u3403_o),
    .c(_al_u3404_o),
    .d(hresp_pad),
    .o(_al_u4831_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4832 (
    .a(_al_u4831_o),
    .b(_al_u3403_o),
    .c(_al_u4099_o),
    .o(_al_u4832_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u4833 (
    .a(_al_u4832_o),
    .b(_al_u2952_o),
    .o(_al_u4833_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u4834 (
    .a(_al_u2847_o),
    .b(\biu/cache_ctrl_logic/statu [2]),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(_al_u4834_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u4835 (
    .a(_al_u4834_o),
    .b(_al_u2847_o),
    .c(_al_u3944_o),
    .o(_al_u4835_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(~C*B))"),
    .INIT(8'h5d))
    _al_u4836 (
    .a(_al_u4833_o),
    .b(_al_u4194_o),
    .c(_al_u4835_o),
    .o(\biu/bus_unit/n35 [1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4837 (
    .a(wb_jmp),
    .b(wb_system),
    .c(wb_int_acc),
    .o(_al_u4837_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u4838 (
    .a(_al_u4837_o),
    .b(wb_m_ret),
    .c(wb_s_ret),
    .o(_al_u4838_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u4839 (
    .a(_al_u4134_o),
    .b(_al_u4136_o),
    .c(_al_u4838_o),
    .d(wb_valid),
    .o(ex_nop));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4840 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [15]),
    .d(\biu/cache_ctrl_logic/l1d_pte [15]),
    .o(_al_u4840_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4841 (
    .a(_al_u2705_o),
    .b(_al_u4840_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [15]),
    .o(_al_u4841_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4842 (
    .a(\exu/lsu/n4 [15]),
    .b(_al_u4841_o),
    .c(_al_u3222_o),
    .o(_al_u4842_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4843 (
    .a(_al_u4842_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [15]),
    .o(hwdata_pad[15]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4844 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [14]),
    .d(\biu/cache_ctrl_logic/pte_temp [14]),
    .o(_al_u4844_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4845 (
    .a(_al_u2705_o),
    .b(_al_u4844_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [14]),
    .o(_al_u4845_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4846 (
    .a(\exu/lsu/n4 [14]),
    .b(_al_u4845_o),
    .c(_al_u3222_o),
    .o(_al_u4846_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4847 (
    .a(_al_u4846_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [14]),
    .o(hwdata_pad[14]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4848 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [13]),
    .d(\biu/cache_ctrl_logic/l1d_pte [13]),
    .o(_al_u4848_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4849 (
    .a(_al_u2705_o),
    .b(_al_u4848_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [13]),
    .o(_al_u4849_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4850 (
    .a(\exu/lsu/n4 [13]),
    .b(_al_u4849_o),
    .c(_al_u3222_o),
    .o(_al_u4850_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4851 (
    .a(_al_u4850_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [13]),
    .o(hwdata_pad[13]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4852 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [12]),
    .d(\biu/cache_ctrl_logic/l1d_pte [12]),
    .o(_al_u4852_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4853 (
    .a(_al_u2705_o),
    .b(_al_u4852_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [12]),
    .o(_al_u4853_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4854 (
    .a(\exu/lsu/n4 [12]),
    .b(_al_u4853_o),
    .c(_al_u3222_o),
    .o(_al_u4854_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4855 (
    .a(_al_u4854_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [12]),
    .o(hwdata_pad[12]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4856 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [11]),
    .d(\biu/cache_ctrl_logic/pte_temp [11]),
    .o(_al_u4856_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4857 (
    .a(_al_u2705_o),
    .b(_al_u4856_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [11]),
    .o(_al_u4857_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4858 (
    .a(\exu/lsu/n4 [11]),
    .b(_al_u4857_o),
    .c(_al_u3222_o),
    .o(_al_u4858_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4859 (
    .a(_al_u4858_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [11]),
    .o(hwdata_pad[11]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4860 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [10]),
    .d(\biu/cache_ctrl_logic/l1d_pte [10]),
    .o(_al_u4860_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4861 (
    .a(_al_u2705_o),
    .b(_al_u4860_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [10]),
    .o(_al_u4861_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4862 (
    .a(\exu/lsu/n4 [10]),
    .b(_al_u4861_o),
    .c(_al_u3222_o),
    .o(_al_u4862_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4863 (
    .a(_al_u4862_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [10]),
    .o(hwdata_pad[10]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4864 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [9]),
    .d(\biu/cache_ctrl_logic/pte_temp [9]),
    .o(_al_u4864_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4865 (
    .a(_al_u2705_o),
    .b(_al_u4864_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [9]),
    .o(_al_u4865_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4866 (
    .a(\exu/lsu/n4 [9]),
    .b(_al_u4865_o),
    .c(_al_u3222_o),
    .o(_al_u4866_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4867 (
    .a(_al_u4866_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [9]),
    .o(hwdata_pad[9]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u4868 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [8]),
    .d(\biu/cache_ctrl_logic/pte_temp [8]),
    .o(_al_u4868_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u4869 (
    .a(_al_u2705_o),
    .b(_al_u4868_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [8]),
    .o(_al_u4869_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u4870 (
    .a(\exu/lsu/n4 [8]),
    .b(_al_u4869_o),
    .c(_al_u3222_o),
    .o(_al_u4870_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u4871 (
    .a(_al_u4870_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [8]),
    .o(hwdata_pad[8]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u4872 (
    .a(id_rs1_index[2]),
    .b(id_rs1_index[1]),
    .c(id_rs1_index[0]),
    .o(_al_u4872_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u4873 (
    .a(_al_u4872_o),
    .b(id_rs1_index[4]),
    .c(id_rs1_index[3]),
    .o(\cu_ru/n45_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4874 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_009 ),
    .c(\cu_ru/al_ram_gpr_do_i1_009 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[9]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u4875 (
    .a(_al_u3214_o),
    .b(_al_u4064_o),
    .o(_al_u4875_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4876 (
    .a(rs1_data[9]),
    .b(_al_u4875_o),
    .c(id_ins_pc[9]),
    .o(\ins_dec/n286 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4877 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_008 ),
    .c(\cu_ru/al_ram_gpr_do_i1_008 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4878 (
    .a(rs1_data[8]),
    .b(_al_u4875_o),
    .c(id_ins_pc[8]),
    .o(\ins_dec/n286 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4879 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_007 ),
    .c(\cu_ru/al_ram_gpr_do_i1_007 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4880 (
    .a(rs1_data[7]),
    .b(_al_u4875_o),
    .c(id_ins_pc[7]),
    .o(\ins_dec/n286 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4881 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_063 ),
    .c(\cu_ru/al_ram_gpr_do_i1_063 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[63]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4882 (
    .a(rs1_data[63]),
    .b(_al_u4875_o),
    .c(id_ins_pc[63]),
    .o(\ins_dec/n286 [63]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4883 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_062 ),
    .c(\cu_ru/al_ram_gpr_do_i1_062 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[62]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4884 (
    .a(rs1_data[62]),
    .b(_al_u4875_o),
    .c(id_ins_pc[62]),
    .o(\ins_dec/n286 [62]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4885 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_061 ),
    .c(\cu_ru/al_ram_gpr_do_i1_061 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[61]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4886 (
    .a(rs1_data[61]),
    .b(_al_u4875_o),
    .c(id_ins_pc[61]),
    .o(\ins_dec/n286 [61]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4887 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_060 ),
    .c(\cu_ru/al_ram_gpr_do_i1_060 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[60]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4888 (
    .a(rs1_data[60]),
    .b(_al_u4875_o),
    .c(id_ins_pc[60]),
    .o(\ins_dec/n286 [60]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4889 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_006 ),
    .c(\cu_ru/al_ram_gpr_do_i1_006 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4890 (
    .a(rs1_data[6]),
    .b(_al_u4875_o),
    .c(id_ins_pc[6]),
    .o(\ins_dec/n286 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4891 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_059 ),
    .c(\cu_ru/al_ram_gpr_do_i1_059 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[59]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4892 (
    .a(rs1_data[59]),
    .b(_al_u4875_o),
    .c(id_ins_pc[59]),
    .o(\ins_dec/n286 [59]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4893 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_058 ),
    .c(\cu_ru/al_ram_gpr_do_i1_058 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[58]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4894 (
    .a(rs1_data[58]),
    .b(_al_u4875_o),
    .c(id_ins_pc[58]),
    .o(\ins_dec/n286 [58]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4895 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_057 ),
    .c(\cu_ru/al_ram_gpr_do_i1_057 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[57]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4896 (
    .a(rs1_data[57]),
    .b(_al_u4875_o),
    .c(id_ins_pc[57]),
    .o(\ins_dec/n286 [57]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4897 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_056 ),
    .c(\cu_ru/al_ram_gpr_do_i1_056 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[56]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4898 (
    .a(rs1_data[56]),
    .b(_al_u4875_o),
    .c(id_ins_pc[56]),
    .o(\ins_dec/n286 [56]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4899 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_055 ),
    .c(\cu_ru/al_ram_gpr_do_i1_055 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[55]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4900 (
    .a(rs1_data[55]),
    .b(_al_u4875_o),
    .c(id_ins_pc[55]),
    .o(\ins_dec/n286 [55]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4901 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_054 ),
    .c(\cu_ru/al_ram_gpr_do_i1_054 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[54]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4902 (
    .a(rs1_data[54]),
    .b(_al_u4875_o),
    .c(id_ins_pc[54]),
    .o(\ins_dec/n286 [54]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4903 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_053 ),
    .c(\cu_ru/al_ram_gpr_do_i1_053 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[53]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4904 (
    .a(rs1_data[53]),
    .b(_al_u4875_o),
    .c(id_ins_pc[53]),
    .o(\ins_dec/n286 [53]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4905 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_052 ),
    .c(\cu_ru/al_ram_gpr_do_i1_052 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[52]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4906 (
    .a(rs1_data[52]),
    .b(_al_u4875_o),
    .c(id_ins_pc[52]),
    .o(\ins_dec/n286 [52]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4907 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_051 ),
    .c(\cu_ru/al_ram_gpr_do_i1_051 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[51]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4908 (
    .a(rs1_data[51]),
    .b(_al_u4875_o),
    .c(id_ins_pc[51]),
    .o(\ins_dec/n286 [51]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4909 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_050 ),
    .c(\cu_ru/al_ram_gpr_do_i1_050 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[50]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4910 (
    .a(rs1_data[50]),
    .b(_al_u4875_o),
    .c(id_ins_pc[50]),
    .o(\ins_dec/n286 [50]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4911 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_005 ),
    .c(\cu_ru/al_ram_gpr_do_i1_005 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4912 (
    .a(rs1_data[5]),
    .b(_al_u4875_o),
    .c(id_ins_pc[5]),
    .o(\ins_dec/n286 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4913 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_049 ),
    .c(\cu_ru/al_ram_gpr_do_i1_049 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[49]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4914 (
    .a(rs1_data[49]),
    .b(_al_u4875_o),
    .c(id_ins_pc[49]),
    .o(\ins_dec/n286 [49]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4915 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_048 ),
    .c(\cu_ru/al_ram_gpr_do_i1_048 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[48]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4916 (
    .a(rs1_data[48]),
    .b(_al_u4875_o),
    .c(id_ins_pc[48]),
    .o(\ins_dec/n286 [48]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4917 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_047 ),
    .c(\cu_ru/al_ram_gpr_do_i1_047 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[47]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4918 (
    .a(rs1_data[47]),
    .b(_al_u4875_o),
    .c(id_ins_pc[47]),
    .o(\ins_dec/n286 [47]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4919 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_046 ),
    .c(\cu_ru/al_ram_gpr_do_i1_046 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[46]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4920 (
    .a(rs1_data[46]),
    .b(_al_u4875_o),
    .c(id_ins_pc[46]),
    .o(\ins_dec/n286 [46]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4921 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_045 ),
    .c(\cu_ru/al_ram_gpr_do_i1_045 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[45]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4922 (
    .a(rs1_data[45]),
    .b(_al_u4875_o),
    .c(id_ins_pc[45]),
    .o(\ins_dec/n286 [45]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4923 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_044 ),
    .c(\cu_ru/al_ram_gpr_do_i1_044 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[44]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4924 (
    .a(rs1_data[44]),
    .b(_al_u4875_o),
    .c(id_ins_pc[44]),
    .o(\ins_dec/n286 [44]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4925 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_043 ),
    .c(\cu_ru/al_ram_gpr_do_i1_043 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[43]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4926 (
    .a(rs1_data[43]),
    .b(_al_u4875_o),
    .c(id_ins_pc[43]),
    .o(\ins_dec/n286 [43]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4927 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_042 ),
    .c(\cu_ru/al_ram_gpr_do_i1_042 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[42]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4928 (
    .a(rs1_data[42]),
    .b(_al_u4875_o),
    .c(id_ins_pc[42]),
    .o(\ins_dec/n286 [42]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4929 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_041 ),
    .c(\cu_ru/al_ram_gpr_do_i1_041 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[41]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4930 (
    .a(rs1_data[41]),
    .b(_al_u4875_o),
    .c(id_ins_pc[41]),
    .o(\ins_dec/n286 [41]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4931 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_040 ),
    .c(\cu_ru/al_ram_gpr_do_i1_040 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[40]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4932 (
    .a(rs1_data[40]),
    .b(_al_u4875_o),
    .c(id_ins_pc[40]),
    .o(\ins_dec/n286 [40]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4933 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_004 ),
    .c(\cu_ru/al_ram_gpr_do_i1_004 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4934 (
    .a(rs1_data[4]),
    .b(_al_u4875_o),
    .c(id_ins_pc[4]),
    .o(\ins_dec/n286 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4935 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_039 ),
    .c(\cu_ru/al_ram_gpr_do_i1_039 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[39]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4936 (
    .a(rs1_data[39]),
    .b(_al_u4875_o),
    .c(id_ins_pc[39]),
    .o(\ins_dec/n286 [39]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4937 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_038 ),
    .c(\cu_ru/al_ram_gpr_do_i1_038 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[38]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4938 (
    .a(rs1_data[38]),
    .b(_al_u4875_o),
    .c(id_ins_pc[38]),
    .o(\ins_dec/n286 [38]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4939 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_037 ),
    .c(\cu_ru/al_ram_gpr_do_i1_037 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[37]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4940 (
    .a(rs1_data[37]),
    .b(_al_u4875_o),
    .c(id_ins_pc[37]),
    .o(\ins_dec/n286 [37]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4941 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_036 ),
    .c(\cu_ru/al_ram_gpr_do_i1_036 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[36]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4942 (
    .a(rs1_data[36]),
    .b(_al_u4875_o),
    .c(id_ins_pc[36]),
    .o(\ins_dec/n286 [36]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4943 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_035 ),
    .c(\cu_ru/al_ram_gpr_do_i1_035 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[35]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4944 (
    .a(rs1_data[35]),
    .b(_al_u4875_o),
    .c(id_ins_pc[35]),
    .o(\ins_dec/n286 [35]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4945 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_034 ),
    .c(\cu_ru/al_ram_gpr_do_i1_034 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[34]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4946 (
    .a(rs1_data[34]),
    .b(_al_u4875_o),
    .c(id_ins_pc[34]),
    .o(\ins_dec/n286 [34]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4947 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_033 ),
    .c(\cu_ru/al_ram_gpr_do_i1_033 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[33]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4948 (
    .a(rs1_data[33]),
    .b(_al_u4875_o),
    .c(id_ins_pc[33]),
    .o(\ins_dec/n286 [33]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4949 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_032 ),
    .c(\cu_ru/al_ram_gpr_do_i1_032 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[32]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4950 (
    .a(rs1_data[32]),
    .b(_al_u4875_o),
    .c(id_ins_pc[32]),
    .o(\ins_dec/n286 [32]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4951 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_031 ),
    .c(\cu_ru/al_ram_gpr_do_i1_031 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4952 (
    .a(rs1_data[31]),
    .b(_al_u4875_o),
    .c(id_ins_pc[31]),
    .o(\ins_dec/n286 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4953 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_030 ),
    .c(\cu_ru/al_ram_gpr_do_i1_030 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4954 (
    .a(rs1_data[30]),
    .b(_al_u4875_o),
    .c(id_ins_pc[30]),
    .o(\ins_dec/n286 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4955 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_003 ),
    .c(\cu_ru/al_ram_gpr_do_i1_003 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4956 (
    .a(rs1_data[3]),
    .b(_al_u4875_o),
    .c(id_ins_pc[3]),
    .o(\ins_dec/n286 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4957 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_029 ),
    .c(\cu_ru/al_ram_gpr_do_i1_029 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[29]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4958 (
    .a(rs1_data[29]),
    .b(_al_u4875_o),
    .c(id_ins_pc[29]),
    .o(\ins_dec/n286 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4959 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_028 ),
    .c(\cu_ru/al_ram_gpr_do_i1_028 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[28]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4960 (
    .a(rs1_data[28]),
    .b(_al_u4875_o),
    .c(id_ins_pc[28]),
    .o(\ins_dec/n286 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4961 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_027 ),
    .c(\cu_ru/al_ram_gpr_do_i1_027 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[27]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4962 (
    .a(rs1_data[27]),
    .b(_al_u4875_o),
    .c(id_ins_pc[27]),
    .o(\ins_dec/n286 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4963 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_026 ),
    .c(\cu_ru/al_ram_gpr_do_i1_026 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[26]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4964 (
    .a(rs1_data[26]),
    .b(_al_u4875_o),
    .c(id_ins_pc[26]),
    .o(\ins_dec/n286 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4965 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_025 ),
    .c(\cu_ru/al_ram_gpr_do_i1_025 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[25]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4966 (
    .a(rs1_data[25]),
    .b(_al_u4875_o),
    .c(id_ins_pc[25]),
    .o(\ins_dec/n286 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4967 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_024 ),
    .c(\cu_ru/al_ram_gpr_do_i1_024 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[24]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4968 (
    .a(rs1_data[24]),
    .b(_al_u4875_o),
    .c(id_ins_pc[24]),
    .o(\ins_dec/n286 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4969 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_023 ),
    .c(\cu_ru/al_ram_gpr_do_i1_023 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[23]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4970 (
    .a(rs1_data[23]),
    .b(_al_u4875_o),
    .c(id_ins_pc[23]),
    .o(\ins_dec/n286 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4971 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_022 ),
    .c(\cu_ru/al_ram_gpr_do_i1_022 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[22]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4972 (
    .a(rs1_data[22]),
    .b(_al_u4875_o),
    .c(id_ins_pc[22]),
    .o(\ins_dec/n286 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4973 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_021 ),
    .c(\cu_ru/al_ram_gpr_do_i1_021 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[21]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4974 (
    .a(rs1_data[21]),
    .b(_al_u4875_o),
    .c(id_ins_pc[21]),
    .o(\ins_dec/n286 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4975 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_020 ),
    .c(\cu_ru/al_ram_gpr_do_i1_020 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[20]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4976 (
    .a(rs1_data[20]),
    .b(_al_u4875_o),
    .c(id_ins_pc[20]),
    .o(\ins_dec/n286 [20]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4977 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_002 ),
    .c(\cu_ru/al_ram_gpr_do_i1_002 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4978 (
    .a(rs1_data[2]),
    .b(_al_u4875_o),
    .c(id_ins_pc[2]),
    .o(\ins_dec/n286 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4979 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_019 ),
    .c(\cu_ru/al_ram_gpr_do_i1_019 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4980 (
    .a(rs1_data[19]),
    .b(_al_u4875_o),
    .c(id_ins_pc[19]),
    .o(\ins_dec/n286 [19]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4981 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_018 ),
    .c(\cu_ru/al_ram_gpr_do_i1_018 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4982 (
    .a(rs1_data[18]),
    .b(_al_u4875_o),
    .c(id_ins_pc[18]),
    .o(\ins_dec/n286 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4983 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_017 ),
    .c(\cu_ru/al_ram_gpr_do_i1_017 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4984 (
    .a(rs1_data[17]),
    .b(_al_u4875_o),
    .c(id_ins_pc[17]),
    .o(\ins_dec/n286 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4985 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_016 ),
    .c(\cu_ru/al_ram_gpr_do_i1_016 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4986 (
    .a(rs1_data[16]),
    .b(_al_u4875_o),
    .c(id_ins_pc[16]),
    .o(\ins_dec/n286 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4987 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_015 ),
    .c(\cu_ru/al_ram_gpr_do_i1_015 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4988 (
    .a(rs1_data[15]),
    .b(_al_u4875_o),
    .c(id_ins_pc[15]),
    .o(\ins_dec/n286 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4989 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_014 ),
    .c(\cu_ru/al_ram_gpr_do_i1_014 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4990 (
    .a(rs1_data[14]),
    .b(_al_u4875_o),
    .c(id_ins_pc[14]),
    .o(\ins_dec/n286 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4991 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_013 ),
    .c(\cu_ru/al_ram_gpr_do_i1_013 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4992 (
    .a(rs1_data[13]),
    .b(_al_u4875_o),
    .c(id_ins_pc[13]),
    .o(\ins_dec/n286 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4993 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_012 ),
    .c(\cu_ru/al_ram_gpr_do_i1_012 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4994 (
    .a(rs1_data[12]),
    .b(_al_u4875_o),
    .c(id_ins_pc[12]),
    .o(\ins_dec/n286 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4995 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_011 ),
    .c(\cu_ru/al_ram_gpr_do_i1_011 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4996 (
    .a(rs1_data[11]),
    .b(_al_u4875_o),
    .c(id_ins_pc[11]),
    .o(\ins_dec/n286 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4997 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_010 ),
    .c(\cu_ru/al_ram_gpr_do_i1_010 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u4998 (
    .a(rs1_data[10]),
    .b(_al_u4875_o),
    .c(id_ins_pc[10]),
    .o(\ins_dec/n286 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u4999 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_001 ),
    .c(\cu_ru/al_ram_gpr_do_i1_001 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u5000 (
    .a(rs1_data[1]),
    .b(_al_u4875_o),
    .c(id_ins_pc[1]),
    .o(\ins_dec/n286 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u5001 (
    .a(\cu_ru/n45_lutinv ),
    .b(\cu_ru/al_ram_gpr_do_i0_000 ),
    .c(\cu_ru/al_ram_gpr_do_i1_000 ),
    .d(\cu_ru/n46 [4]),
    .o(rs1_data[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u5002 (
    .a(rs1_data[0]),
    .b(_al_u4875_o),
    .c(id_ins_pc[0]),
    .o(\ins_dec/n286 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcf44))
    _al_u5003 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [63]),
    .o(_al_u5003_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u5004 (
    .a(\biu/maddress [63]),
    .b(_al_u5003_o),
    .c(_al_u2914_o),
    .d(_al_u2698_o),
    .o(\biu/bus_unit/mmu/n66 [63]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcf44))
    _al_u5005 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [62]),
    .o(_al_u5005_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u5006 (
    .a(\biu/maddress [62]),
    .b(_al_u5005_o),
    .c(_al_u2914_o),
    .d(_al_u2698_o),
    .o(\biu/bus_unit/mmu/n66 [62]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcf44))
    _al_u5007 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [61]),
    .o(_al_u5007_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u5008 (
    .a(\biu/maddress [61]),
    .b(_al_u5007_o),
    .c(_al_u2914_o),
    .d(_al_u2698_o),
    .o(\biu/bus_unit/mmu/n66 [61]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcf44))
    _al_u5009 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [60]),
    .o(_al_u5009_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u5010 (
    .a(\biu/maddress [60]),
    .b(_al_u5009_o),
    .c(_al_u2914_o),
    .d(_al_u2698_o),
    .o(\biu/bus_unit/mmu/n66 [60]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcf44))
    _al_u5011 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [59]),
    .o(_al_u5011_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u5012 (
    .a(\biu/maddress [59]),
    .b(_al_u5011_o),
    .c(_al_u2914_o),
    .d(_al_u2698_o),
    .o(\biu/bus_unit/mmu/n66 [59]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcf44))
    _al_u5013 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [58]),
    .o(_al_u5013_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u5014 (
    .a(\biu/maddress [58]),
    .b(_al_u5013_o),
    .c(_al_u2914_o),
    .d(_al_u2698_o),
    .o(\biu/bus_unit/mmu/n66 [58]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcf44))
    _al_u5015 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [57]),
    .o(_al_u5015_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u5016 (
    .a(\biu/maddress [57]),
    .b(_al_u5015_o),
    .c(_al_u2914_o),
    .d(_al_u2698_o),
    .o(\biu/bus_unit/mmu/n66 [57]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcf44))
    _al_u5017 (
    .a(_al_u2914_o),
    .b(_al_u2698_o),
    .c(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .d(\biu/paddress [56]),
    .o(_al_u5017_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u5018 (
    .a(\biu/maddress [56]),
    .b(_al_u5017_o),
    .c(_al_u2914_o),
    .d(_al_u2698_o),
    .o(\biu/bus_unit/mmu/n66 [56]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5019 (
    .a(\biu/maddress [55]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [55]),
    .o(_al_u5019_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5020 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [55]),
    .d(\biu/bus_unit/mmu_hwdata [53]),
    .o(_al_u5020_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5021 (
    .a(_al_u5019_o),
    .b(_al_u5020_o),
    .o(\biu/bus_unit/mmu/n66 [55]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5022 (
    .a(\biu/maddress [54]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [54]),
    .o(_al_u5022_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5023 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [54]),
    .d(\biu/bus_unit/mmu_hwdata [52]),
    .o(_al_u5023_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5024 (
    .a(_al_u5022_o),
    .b(_al_u5023_o),
    .o(\biu/bus_unit/mmu/n66 [54]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5025 (
    .a(\biu/maddress [53]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [53]),
    .o(_al_u5025_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5026 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [53]),
    .d(\biu/bus_unit/mmu_hwdata [51]),
    .o(_al_u5026_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5027 (
    .a(_al_u5025_o),
    .b(_al_u5026_o),
    .o(\biu/bus_unit/mmu/n66 [53]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5028 (
    .a(\biu/maddress [52]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [52]),
    .o(_al_u5028_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5029 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [52]),
    .d(\biu/bus_unit/mmu_hwdata [50]),
    .o(_al_u5029_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5030 (
    .a(_al_u5028_o),
    .b(_al_u5029_o),
    .o(\biu/bus_unit/mmu/n66 [52]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5031 (
    .a(\biu/maddress [51]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [51]),
    .o(_al_u5031_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5032 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [51]),
    .d(\biu/bus_unit/mmu_hwdata [49]),
    .o(_al_u5032_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5033 (
    .a(_al_u5031_o),
    .b(_al_u5032_o),
    .o(\biu/bus_unit/mmu/n66 [51]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5034 (
    .a(\biu/maddress [50]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [50]),
    .o(_al_u5034_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5035 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [50]),
    .d(\biu/bus_unit/mmu_hwdata [48]),
    .o(_al_u5035_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5036 (
    .a(_al_u5034_o),
    .b(_al_u5035_o),
    .o(\biu/bus_unit/mmu/n66 [50]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5037 (
    .a(\biu/maddress [49]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [49]),
    .o(_al_u5037_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5038 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [49]),
    .d(\biu/bus_unit/mmu_hwdata [47]),
    .o(_al_u5038_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5039 (
    .a(_al_u5037_o),
    .b(_al_u5038_o),
    .o(\biu/bus_unit/mmu/n66 [49]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5040 (
    .a(\biu/maddress [48]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [48]),
    .o(_al_u5040_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5041 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [48]),
    .d(\biu/bus_unit/mmu_hwdata [46]),
    .o(_al_u5041_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5042 (
    .a(_al_u5040_o),
    .b(_al_u5041_o),
    .o(\biu/bus_unit/mmu/n66 [48]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5043 (
    .a(\biu/maddress [47]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [47]),
    .o(_al_u5043_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5044 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [47]),
    .d(\biu/bus_unit/mmu_hwdata [45]),
    .o(_al_u5044_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5045 (
    .a(_al_u5043_o),
    .b(_al_u5044_o),
    .o(\biu/bus_unit/mmu/n66 [47]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5046 (
    .a(\biu/maddress [46]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [46]),
    .o(_al_u5046_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5047 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [46]),
    .d(\biu/bus_unit/mmu_hwdata [44]),
    .o(_al_u5047_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5048 (
    .a(_al_u5046_o),
    .b(_al_u5047_o),
    .o(\biu/bus_unit/mmu/n66 [46]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5049 (
    .a(\biu/maddress [45]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [45]),
    .o(_al_u5049_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5050 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [45]),
    .d(\biu/bus_unit/mmu_hwdata [43]),
    .o(_al_u5050_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5051 (
    .a(_al_u5049_o),
    .b(_al_u5050_o),
    .o(\biu/bus_unit/mmu/n66 [45]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5052 (
    .a(\biu/maddress [44]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [44]),
    .o(_al_u5052_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5053 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [44]),
    .d(\biu/bus_unit/mmu_hwdata [42]),
    .o(_al_u5053_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5054 (
    .a(_al_u5052_o),
    .b(_al_u5053_o),
    .o(\biu/bus_unit/mmu/n66 [44]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5055 (
    .a(\biu/maddress [43]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [43]),
    .o(_al_u5055_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5056 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [43]),
    .d(\biu/bus_unit/mmu_hwdata [41]),
    .o(_al_u5056_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5057 (
    .a(_al_u5055_o),
    .b(_al_u5056_o),
    .o(\biu/bus_unit/mmu/n66 [43]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5058 (
    .a(\biu/maddress [42]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [42]),
    .o(_al_u5058_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5059 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [42]),
    .d(\biu/bus_unit/mmu_hwdata [40]),
    .o(_al_u5059_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5060 (
    .a(_al_u5058_o),
    .b(_al_u5059_o),
    .o(\biu/bus_unit/mmu/n66 [42]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5061 (
    .a(\biu/maddress [41]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [41]),
    .o(_al_u5061_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5062 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [41]),
    .d(\biu/bus_unit/mmu_hwdata [39]),
    .o(_al_u5062_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5063 (
    .a(_al_u5061_o),
    .b(_al_u5062_o),
    .o(\biu/bus_unit/mmu/n66 [41]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5064 (
    .a(\biu/maddress [40]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [40]),
    .o(_al_u5064_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5065 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [40]),
    .d(\biu/bus_unit/mmu_hwdata [38]),
    .o(_al_u5065_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5066 (
    .a(_al_u5064_o),
    .b(_al_u5065_o),
    .o(\biu/bus_unit/mmu/n66 [40]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5067 (
    .a(\biu/maddress [39]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [39]),
    .o(_al_u5067_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5068 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [39]),
    .d(\biu/bus_unit/mmu_hwdata [37]),
    .o(_al_u5068_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5069 (
    .a(_al_u5067_o),
    .b(_al_u5068_o),
    .o(\biu/bus_unit/mmu/n66 [39]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5070 (
    .a(\biu/maddress [38]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [38]),
    .o(_al_u5070_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5071 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [38]),
    .d(\biu/bus_unit/mmu_hwdata [36]),
    .o(_al_u5071_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5072 (
    .a(_al_u5070_o),
    .b(_al_u5071_o),
    .o(\biu/bus_unit/mmu/n66 [38]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5073 (
    .a(\biu/maddress [37]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [37]),
    .o(_al_u5073_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5074 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [37]),
    .d(\biu/bus_unit/mmu_hwdata [35]),
    .o(_al_u5074_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5075 (
    .a(_al_u5073_o),
    .b(_al_u5074_o),
    .o(\biu/bus_unit/mmu/n66 [37]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5076 (
    .a(\biu/maddress [36]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [36]),
    .o(_al_u5076_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5077 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [36]),
    .d(\biu/bus_unit/mmu_hwdata [34]),
    .o(_al_u5077_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5078 (
    .a(_al_u5076_o),
    .b(_al_u5077_o),
    .o(\biu/bus_unit/mmu/n66 [36]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5079 (
    .a(\biu/maddress [35]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [35]),
    .o(_al_u5079_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5080 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [35]),
    .d(\biu/bus_unit/mmu_hwdata [33]),
    .o(_al_u5080_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5081 (
    .a(_al_u5079_o),
    .b(_al_u5080_o),
    .o(\biu/bus_unit/mmu/n66 [35]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5082 (
    .a(\biu/maddress [34]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [34]),
    .o(_al_u5082_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5083 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [34]),
    .d(\biu/bus_unit/mmu_hwdata [32]),
    .o(_al_u5083_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5084 (
    .a(_al_u5082_o),
    .b(_al_u5083_o),
    .o(\biu/bus_unit/mmu/n66 [34]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5085 (
    .a(\biu/maddress [33]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [33]),
    .o(_al_u5085_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5086 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [33]),
    .d(\biu/bus_unit/mmu_hwdata [31]),
    .o(_al_u5086_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5087 (
    .a(_al_u5085_o),
    .b(_al_u5086_o),
    .o(\biu/bus_unit/mmu/n66 [33]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5088 (
    .a(\biu/maddress [32]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [32]),
    .o(_al_u5088_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5089 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [32]),
    .d(\biu/bus_unit/mmu_hwdata [30]),
    .o(_al_u5089_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5090 (
    .a(_al_u5088_o),
    .b(_al_u5089_o),
    .o(\biu/bus_unit/mmu/n66 [32]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5091 (
    .a(\biu/maddress [31]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [31]),
    .o(_al_u5091_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5092 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [31]),
    .d(\biu/bus_unit/mmu_hwdata [29]),
    .o(_al_u5092_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5093 (
    .a(_al_u5091_o),
    .b(_al_u5092_o),
    .o(\biu/bus_unit/mmu/n66 [31]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5094 (
    .a(\biu/maddress [30]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [30]),
    .o(_al_u5094_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5095 (
    .a(_al_u2698_o),
    .b(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .c(\biu/paddress [30]),
    .d(\biu/bus_unit/mmu_hwdata [28]),
    .o(_al_u5095_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5096 (
    .a(_al_u5094_o),
    .b(_al_u5095_o),
    .o(\biu/bus_unit/mmu/n66 [30]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u5097 (
    .a(ex_nop),
    .b(rst_pad),
    .o(\exu/n86 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5098 (
    .a(_al_u4137_o),
    .b(wb_int_acc),
    .o(_al_u5098_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(C*~B)))"),
    .INIT(16'h1055))
    _al_u5099 (
    .a(\cu_ru/medeleg_exc_ctrl/iaf_target_m_lutinv ),
    .b(priv[3]),
    .c(\cu_ru/medeleg [12]),
    .d(wb_ins_page_fault),
    .o(_al_u5099_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(C*~B)))"),
    .INIT(16'h1055))
    _al_u5100 (
    .a(\cu_ru/medeleg_exc_ctrl/lam_target_m_lutinv ),
    .b(priv[3]),
    .c(\cu_ru/medeleg [3]),
    .d(wb_ebreak),
    .o(_al_u5100_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(C*~B)))"),
    .INIT(16'h1055))
    _al_u5101 (
    .a(\cu_ru/medeleg_exc_ctrl/spf_target_m_lutinv ),
    .b(priv[3]),
    .c(\cu_ru/medeleg [6]),
    .d(wb_st_addr_mis),
    .o(_al_u5101_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5102 (
    .a(_al_u5099_o),
    .b(_al_u5100_o),
    .c(_al_u5101_o),
    .o(_al_u5102_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u5103 (
    .a(priv[0]),
    .b(\cu_ru/medeleg [8]),
    .c(wb_ecall),
    .o(\cu_ru/medeleg_exc_ctrl/ecu_target_m ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*A))"),
    .INIT(16'h0301))
    _al_u5104 (
    .a(_al_u4229_o),
    .b(\cu_ru/medeleg_exc_ctrl/iam_target_m_lutinv ),
    .c(\cu_ru/medeleg_exc_ctrl/ecu_target_m ),
    .d(\cu_ru/medeleg [9]),
    .o(_al_u5104_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(C*~B)))"),
    .INIT(16'h1055))
    _al_u5105 (
    .a(\cu_ru/medeleg_exc_ctrl/saf_target_m_lutinv ),
    .b(priv[3]),
    .c(\cu_ru/medeleg [13]),
    .d(wb_ld_page_fault),
    .o(_al_u5105_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(C*~B)))"),
    .INIT(16'h1055))
    _al_u5106 (
    .a(\cu_ru/medeleg_exc_ctrl/laf_target_m_lutinv ),
    .b(priv[3]),
    .c(\cu_ru/medeleg [2]),
    .d(wb_ill_ins),
    .o(_al_u5106_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5107 (
    .a(_al_u5104_o),
    .b(_al_u5105_o),
    .c(_al_u5106_o),
    .o(_al_u5107_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(B*~A))"),
    .INIT(16'hb000))
    _al_u5108 (
    .a(\cu_ru/mideleg_int_ctrl/n28_lutinv ),
    .b(_al_u5098_o),
    .c(_al_u5102_o),
    .d(_al_u5107_o),
    .o(_al_u5108_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u5109 (
    .a(_al_u5108_o),
    .b(wb_valid),
    .o(\cu_ru/trap_target_m ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5110 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [17]),
    .d(\biu/cache_ctrl_logic/l1d_pte [17]),
    .o(_al_u5110_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5111 (
    .a(_al_u2705_o),
    .b(_al_u5110_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [17]),
    .o(_al_u5111_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5112 (
    .a(_al_u4205_o),
    .b(_al_u5111_o),
    .c(_al_u3222_o),
    .o(_al_u5112_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5113 (
    .a(_al_u5112_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [17]),
    .o(hwdata_pad[17]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5114 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [16]),
    .d(\biu/cache_ctrl_logic/pte_temp [16]),
    .o(_al_u5114_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5115 (
    .a(_al_u2705_o),
    .b(_al_u5114_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [16]),
    .o(_al_u5115_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5116 (
    .a(_al_u4208_o),
    .b(_al_u5115_o),
    .c(_al_u3222_o),
    .o(_al_u5116_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5117 (
    .a(_al_u5116_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [16]),
    .o(hwdata_pad[16]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5118 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [23]),
    .d(\biu/cache_ctrl_logic/pte_temp [23]),
    .o(_al_u5118_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5119 (
    .a(_al_u2705_o),
    .b(_al_u5118_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [23]),
    .o(_al_u5119_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5120 (
    .a(_al_u4211_o),
    .b(_al_u5119_o),
    .c(_al_u3222_o),
    .o(_al_u5120_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5121 (
    .a(_al_u5120_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [23]),
    .o(hwdata_pad[23]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5122 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [22]),
    .d(\biu/cache_ctrl_logic/l1d_pte [22]),
    .o(_al_u5122_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5123 (
    .a(_al_u2705_o),
    .b(_al_u5122_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [22]),
    .o(_al_u5123_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5124 (
    .a(_al_u4214_o),
    .b(_al_u5123_o),
    .c(_al_u3222_o),
    .o(_al_u5124_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5125 (
    .a(_al_u5124_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [22]),
    .o(hwdata_pad[22]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5126 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [21]),
    .d(\biu/cache_ctrl_logic/pte_temp [21]),
    .o(_al_u5126_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5127 (
    .a(_al_u2705_o),
    .b(_al_u5126_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [21]),
    .o(_al_u5127_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5128 (
    .a(_al_u4217_o),
    .b(_al_u5127_o),
    .c(_al_u3222_o),
    .o(_al_u5128_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5129 (
    .a(_al_u5128_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [21]),
    .o(hwdata_pad[21]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5130 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [20]),
    .d(\biu/cache_ctrl_logic/l1d_pte [20]),
    .o(_al_u5130_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5131 (
    .a(_al_u2705_o),
    .b(_al_u5130_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [20]),
    .o(_al_u5131_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5132 (
    .a(_al_u4220_o),
    .b(_al_u5131_o),
    .c(_al_u3222_o),
    .o(_al_u5132_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5133 (
    .a(_al_u5132_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [20]),
    .o(hwdata_pad[20]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5134 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [19]),
    .d(\biu/cache_ctrl_logic/l1d_pte [19]),
    .o(_al_u5134_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5135 (
    .a(_al_u2705_o),
    .b(_al_u5134_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [19]),
    .o(_al_u5135_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5136 (
    .a(_al_u4223_o),
    .b(_al_u5135_o),
    .c(_al_u3222_o),
    .o(_al_u5136_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5137 (
    .a(_al_u5136_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [19]),
    .o(hwdata_pad[19]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5138 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [18]),
    .d(\biu/cache_ctrl_logic/pte_temp [18]),
    .o(_al_u5138_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5139 (
    .a(_al_u2705_o),
    .b(_al_u5138_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [18]),
    .o(_al_u5139_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5140 (
    .a(_al_u4226_o),
    .b(_al_u5139_o),
    .c(_al_u3222_o),
    .o(_al_u5140_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5141 (
    .a(_al_u5140_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [18]),
    .o(hwdata_pad[18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u5142 (
    .a(id_ins[22]),
    .b(id_ins[20]),
    .c(_al_u3392_o),
    .o(_al_u5142_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5143 (
    .a(_al_u5142_o),
    .b(id_ins[21]),
    .o(_al_u5143_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5144 (
    .a(_al_u4086_o),
    .b(_al_u5143_o),
    .o(_al_u5144_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5145 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_007 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_007 ),
    .d(\cu_ru/n49 [4]),
    .o(\ins_dec/op_count_decode [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5146 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_006 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_006 ),
    .d(\cu_ru/n49 [4]),
    .o(\ins_dec/op_count_decode [6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u5147 (
    .a(\cu_ru/mideleg_int_ctrl/n28_lutinv ),
    .b(_al_u3250_o),
    .c(_al_u5098_o),
    .o(_al_u5147_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u5148 (
    .a(priv[0]),
    .b(\cu_ru/medeleg [8]),
    .c(wb_ecall),
    .o(\cu_ru/medeleg_exc_ctrl/ecu_target_s ));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u5149 (
    .a(\cu_ru/medeleg_exc_ctrl/iam_target_s ),
    .b(_al_u4229_o),
    .c(\cu_ru/medeleg_exc_ctrl/ecu_target_s ),
    .d(\cu_ru/medeleg [9]),
    .o(_al_u5149_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u5150 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(\cu_ru/medeleg [2]),
    .c(wb_ill_ins),
    .o(\cu_ru/medeleg_exc_ctrl/ii_target_s ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*~(D*C)))"),
    .INIT(16'h5444))
    _al_u5151 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(_al_u4108_o),
    .c(\cu_ru/medeleg [13]),
    .d(wb_ld_page_fault),
    .o(_al_u5151_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u5152 (
    .a(_al_u5149_o),
    .b(\cu_ru/medeleg_exc_ctrl/laf_target_s ),
    .c(\cu_ru/medeleg_exc_ctrl/ii_target_s ),
    .d(_al_u5151_o),
    .o(_al_u5152_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u5153 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(\cu_ru/medeleg [6]),
    .c(wb_st_addr_mis),
    .o(\cu_ru/medeleg_exc_ctrl/sam_target_s ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*~(D*C)))"),
    .INIT(16'h5444))
    _al_u5154 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(_al_u4119_o),
    .c(\cu_ru/medeleg [12]),
    .d(wb_ins_page_fault),
    .o(_al_u5154_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*~(D*C)))"),
    .INIT(16'h5444))
    _al_u5155 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(_al_u4123_o),
    .c(\cu_ru/medeleg [3]),
    .d(wb_ebreak),
    .o(_al_u5155_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u5156 (
    .a(\cu_ru/medeleg_exc_ctrl/sam_target_s ),
    .b(\cu_ru/medeleg_exc_ctrl/spf_target_s ),
    .c(_al_u5154_o),
    .d(_al_u5155_o),
    .o(_al_u5156_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u5157 (
    .a(_al_u5147_o),
    .b(_al_u5152_o),
    .c(_al_u5156_o),
    .d(wb_valid),
    .o(_al_u5157_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5158 (
    .a(_al_u3420_o),
    .b(_al_u3184_o),
    .o(_al_u5158_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5159 (
    .a(_al_u5158_o),
    .b(_al_u3204_o),
    .o(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5160 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [9]),
    .c(data_csr[9]),
    .o(_al_u5160_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5161 (
    .a(_al_u4133_o),
    .b(wb_ebreak),
    .o(_al_u5161_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5162 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[9]),
    .c(wb_exc_code[9]),
    .o(\cu_ru/m_s_tval/n3 [9]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5163 (
    .a(_al_u5157_o),
    .b(_al_u5160_o),
    .c(\cu_ru/m_s_tval/n3 [9]),
    .o(\cu_ru/m_s_tval/n9 [9]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5164 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [8]),
    .c(data_csr[8]),
    .o(_al_u5164_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5165 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[8]),
    .c(wb_exc_code[8]),
    .o(\cu_ru/m_s_tval/n3 [8]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5166 (
    .a(_al_u5157_o),
    .b(_al_u5164_o),
    .c(\cu_ru/m_s_tval/n3 [8]),
    .o(\cu_ru/m_s_tval/n9 [8]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5167 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [7]),
    .c(data_csr[7]),
    .o(_al_u5167_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5168 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[7]),
    .c(wb_exc_code[7]),
    .o(\cu_ru/m_s_tval/n3 [7]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5169 (
    .a(_al_u5157_o),
    .b(_al_u5167_o),
    .c(\cu_ru/m_s_tval/n3 [7]),
    .o(\cu_ru/m_s_tval/n9 [7]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5170 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [63]),
    .c(data_csr[63]),
    .o(_al_u5170_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5171 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[63]),
    .c(wb_exc_code[63]),
    .o(\cu_ru/m_s_tval/n3 [63]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5172 (
    .a(_al_u5157_o),
    .b(_al_u5170_o),
    .c(\cu_ru/m_s_tval/n3 [63]),
    .o(\cu_ru/m_s_tval/n9 [63]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5173 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [62]),
    .c(data_csr[62]),
    .o(_al_u5173_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5174 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[62]),
    .c(wb_exc_code[62]),
    .o(\cu_ru/m_s_tval/n3 [62]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5175 (
    .a(_al_u5157_o),
    .b(_al_u5173_o),
    .c(\cu_ru/m_s_tval/n3 [62]),
    .o(\cu_ru/m_s_tval/n9 [62]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5176 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [61]),
    .c(data_csr[61]),
    .o(_al_u5176_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5177 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[61]),
    .c(wb_exc_code[61]),
    .o(\cu_ru/m_s_tval/n3 [61]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5178 (
    .a(_al_u5157_o),
    .b(_al_u5176_o),
    .c(\cu_ru/m_s_tval/n3 [61]),
    .o(\cu_ru/m_s_tval/n9 [61]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5179 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [60]),
    .c(data_csr[60]),
    .o(_al_u5179_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5180 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[60]),
    .c(wb_exc_code[60]),
    .o(\cu_ru/m_s_tval/n3 [60]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5181 (
    .a(_al_u5157_o),
    .b(_al_u5179_o),
    .c(\cu_ru/m_s_tval/n3 [60]),
    .o(\cu_ru/m_s_tval/n9 [60]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5182 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [6]),
    .c(data_csr[6]),
    .o(_al_u5182_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5183 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[6]),
    .c(wb_exc_code[6]),
    .o(\cu_ru/m_s_tval/n3 [6]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5184 (
    .a(_al_u5157_o),
    .b(_al_u5182_o),
    .c(\cu_ru/m_s_tval/n3 [6]),
    .o(\cu_ru/m_s_tval/n9 [6]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5185 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [59]),
    .c(data_csr[59]),
    .o(_al_u5185_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5186 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[59]),
    .c(wb_exc_code[59]),
    .o(\cu_ru/m_s_tval/n3 [59]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5187 (
    .a(_al_u5157_o),
    .b(_al_u5185_o),
    .c(\cu_ru/m_s_tval/n3 [59]),
    .o(\cu_ru/m_s_tval/n9 [59]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5188 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [58]),
    .c(data_csr[58]),
    .o(_al_u5188_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5189 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[58]),
    .c(wb_exc_code[58]),
    .o(\cu_ru/m_s_tval/n3 [58]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5190 (
    .a(_al_u5157_o),
    .b(_al_u5188_o),
    .c(\cu_ru/m_s_tval/n3 [58]),
    .o(\cu_ru/m_s_tval/n9 [58]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5191 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [57]),
    .c(data_csr[57]),
    .o(_al_u5191_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5192 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[57]),
    .c(wb_exc_code[57]),
    .o(\cu_ru/m_s_tval/n3 [57]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5193 (
    .a(_al_u5157_o),
    .b(_al_u5191_o),
    .c(\cu_ru/m_s_tval/n3 [57]),
    .o(\cu_ru/m_s_tval/n9 [57]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5194 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [56]),
    .c(data_csr[56]),
    .o(_al_u5194_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5195 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[56]),
    .c(wb_exc_code[56]),
    .o(\cu_ru/m_s_tval/n3 [56]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5196 (
    .a(_al_u5157_o),
    .b(_al_u5194_o),
    .c(\cu_ru/m_s_tval/n3 [56]),
    .o(\cu_ru/m_s_tval/n9 [56]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5197 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [55]),
    .c(data_csr[55]),
    .o(_al_u5197_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5198 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[55]),
    .c(wb_exc_code[55]),
    .o(\cu_ru/m_s_tval/n3 [55]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5199 (
    .a(_al_u5157_o),
    .b(_al_u5197_o),
    .c(\cu_ru/m_s_tval/n3 [55]),
    .o(\cu_ru/m_s_tval/n9 [55]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5200 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [54]),
    .c(data_csr[54]),
    .o(_al_u5200_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5201 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[54]),
    .c(wb_exc_code[54]),
    .o(\cu_ru/m_s_tval/n3 [54]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5202 (
    .a(_al_u5157_o),
    .b(_al_u5200_o),
    .c(\cu_ru/m_s_tval/n3 [54]),
    .o(\cu_ru/m_s_tval/n9 [54]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5203 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [53]),
    .c(data_csr[53]),
    .o(_al_u5203_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5204 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[53]),
    .c(wb_exc_code[53]),
    .o(\cu_ru/m_s_tval/n3 [53]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5205 (
    .a(_al_u5157_o),
    .b(_al_u5203_o),
    .c(\cu_ru/m_s_tval/n3 [53]),
    .o(\cu_ru/m_s_tval/n9 [53]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5206 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [52]),
    .c(data_csr[52]),
    .o(_al_u5206_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5207 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[52]),
    .c(wb_exc_code[52]),
    .o(\cu_ru/m_s_tval/n3 [52]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5208 (
    .a(_al_u5157_o),
    .b(_al_u5206_o),
    .c(\cu_ru/m_s_tval/n3 [52]),
    .o(\cu_ru/m_s_tval/n9 [52]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5209 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [51]),
    .c(data_csr[51]),
    .o(_al_u5209_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5210 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[51]),
    .c(wb_exc_code[51]),
    .o(\cu_ru/m_s_tval/n3 [51]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5211 (
    .a(_al_u5157_o),
    .b(_al_u5209_o),
    .c(\cu_ru/m_s_tval/n3 [51]),
    .o(\cu_ru/m_s_tval/n9 [51]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5212 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [50]),
    .c(data_csr[50]),
    .o(_al_u5212_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5213 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[50]),
    .c(wb_exc_code[50]),
    .o(\cu_ru/m_s_tval/n3 [50]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5214 (
    .a(_al_u5157_o),
    .b(_al_u5212_o),
    .c(\cu_ru/m_s_tval/n3 [50]),
    .o(\cu_ru/m_s_tval/n9 [50]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5215 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [5]),
    .c(data_csr[5]),
    .o(_al_u5215_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5216 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[5]),
    .c(wb_exc_code[5]),
    .o(\cu_ru/m_s_tval/n3 [5]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5217 (
    .a(_al_u5157_o),
    .b(_al_u5215_o),
    .c(\cu_ru/m_s_tval/n3 [5]),
    .o(\cu_ru/m_s_tval/n9 [5]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5218 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [49]),
    .c(data_csr[49]),
    .o(_al_u5218_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5219 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[49]),
    .c(wb_exc_code[49]),
    .o(\cu_ru/m_s_tval/n3 [49]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5220 (
    .a(_al_u5157_o),
    .b(_al_u5218_o),
    .c(\cu_ru/m_s_tval/n3 [49]),
    .o(\cu_ru/m_s_tval/n9 [49]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5221 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [48]),
    .c(data_csr[48]),
    .o(_al_u5221_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5222 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[48]),
    .c(wb_exc_code[48]),
    .o(\cu_ru/m_s_tval/n3 [48]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5223 (
    .a(_al_u5157_o),
    .b(_al_u5221_o),
    .c(\cu_ru/m_s_tval/n3 [48]),
    .o(\cu_ru/m_s_tval/n9 [48]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5224 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [47]),
    .c(data_csr[47]),
    .o(_al_u5224_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5225 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[47]),
    .c(wb_exc_code[47]),
    .o(\cu_ru/m_s_tval/n3 [47]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5226 (
    .a(_al_u5157_o),
    .b(_al_u5224_o),
    .c(\cu_ru/m_s_tval/n3 [47]),
    .o(\cu_ru/m_s_tval/n9 [47]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5227 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [46]),
    .c(data_csr[46]),
    .o(_al_u5227_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5228 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[46]),
    .c(wb_exc_code[46]),
    .o(\cu_ru/m_s_tval/n3 [46]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5229 (
    .a(_al_u5157_o),
    .b(_al_u5227_o),
    .c(\cu_ru/m_s_tval/n3 [46]),
    .o(\cu_ru/m_s_tval/n9 [46]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5230 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [45]),
    .c(data_csr[45]),
    .o(_al_u5230_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5231 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[45]),
    .c(wb_exc_code[45]),
    .o(\cu_ru/m_s_tval/n3 [45]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5232 (
    .a(_al_u5157_o),
    .b(_al_u5230_o),
    .c(\cu_ru/m_s_tval/n3 [45]),
    .o(\cu_ru/m_s_tval/n9 [45]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5233 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [44]),
    .c(data_csr[44]),
    .o(_al_u5233_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5234 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[44]),
    .c(wb_exc_code[44]),
    .o(\cu_ru/m_s_tval/n3 [44]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5235 (
    .a(_al_u5157_o),
    .b(_al_u5233_o),
    .c(\cu_ru/m_s_tval/n3 [44]),
    .o(\cu_ru/m_s_tval/n9 [44]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5236 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [43]),
    .c(data_csr[43]),
    .o(_al_u5236_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5237 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[43]),
    .c(wb_exc_code[43]),
    .o(\cu_ru/m_s_tval/n3 [43]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5238 (
    .a(_al_u5157_o),
    .b(_al_u5236_o),
    .c(\cu_ru/m_s_tval/n3 [43]),
    .o(\cu_ru/m_s_tval/n9 [43]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5239 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [42]),
    .c(data_csr[42]),
    .o(_al_u5239_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5240 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[42]),
    .c(wb_exc_code[42]),
    .o(\cu_ru/m_s_tval/n3 [42]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5241 (
    .a(_al_u5157_o),
    .b(_al_u5239_o),
    .c(\cu_ru/m_s_tval/n3 [42]),
    .o(\cu_ru/m_s_tval/n9 [42]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5242 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [41]),
    .c(data_csr[41]),
    .o(_al_u5242_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5243 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[41]),
    .c(wb_exc_code[41]),
    .o(\cu_ru/m_s_tval/n3 [41]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5244 (
    .a(_al_u5157_o),
    .b(_al_u5242_o),
    .c(\cu_ru/m_s_tval/n3 [41]),
    .o(\cu_ru/m_s_tval/n9 [41]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5245 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [40]),
    .c(data_csr[40]),
    .o(_al_u5245_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5246 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[40]),
    .c(wb_exc_code[40]),
    .o(\cu_ru/m_s_tval/n3 [40]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5247 (
    .a(_al_u5157_o),
    .b(_al_u5245_o),
    .c(\cu_ru/m_s_tval/n3 [40]),
    .o(\cu_ru/m_s_tval/n9 [40]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5248 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [4]),
    .c(data_csr[4]),
    .o(_al_u5248_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5249 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[4]),
    .c(wb_exc_code[4]),
    .o(\cu_ru/m_s_tval/n3 [4]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5250 (
    .a(_al_u5157_o),
    .b(_al_u5248_o),
    .c(\cu_ru/m_s_tval/n3 [4]),
    .o(\cu_ru/m_s_tval/n9 [4]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5251 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [39]),
    .c(data_csr[39]),
    .o(_al_u5251_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5252 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[39]),
    .c(wb_exc_code[39]),
    .o(\cu_ru/m_s_tval/n3 [39]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5253 (
    .a(_al_u5157_o),
    .b(_al_u5251_o),
    .c(\cu_ru/m_s_tval/n3 [39]),
    .o(\cu_ru/m_s_tval/n9 [39]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5254 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [38]),
    .c(data_csr[38]),
    .o(_al_u5254_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5255 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[38]),
    .c(wb_exc_code[38]),
    .o(\cu_ru/m_s_tval/n3 [38]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5256 (
    .a(_al_u5157_o),
    .b(_al_u5254_o),
    .c(\cu_ru/m_s_tval/n3 [38]),
    .o(\cu_ru/m_s_tval/n9 [38]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5257 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [37]),
    .c(data_csr[37]),
    .o(_al_u5257_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5258 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[37]),
    .c(wb_exc_code[37]),
    .o(\cu_ru/m_s_tval/n3 [37]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5259 (
    .a(_al_u5157_o),
    .b(_al_u5257_o),
    .c(\cu_ru/m_s_tval/n3 [37]),
    .o(\cu_ru/m_s_tval/n9 [37]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5260 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [36]),
    .c(data_csr[36]),
    .o(_al_u5260_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5261 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[36]),
    .c(wb_exc_code[36]),
    .o(\cu_ru/m_s_tval/n3 [36]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5262 (
    .a(_al_u5157_o),
    .b(_al_u5260_o),
    .c(\cu_ru/m_s_tval/n3 [36]),
    .o(\cu_ru/m_s_tval/n9 [36]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5263 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [35]),
    .c(data_csr[35]),
    .o(_al_u5263_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5264 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[35]),
    .c(wb_exc_code[35]),
    .o(\cu_ru/m_s_tval/n3 [35]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5265 (
    .a(_al_u5157_o),
    .b(_al_u5263_o),
    .c(\cu_ru/m_s_tval/n3 [35]),
    .o(\cu_ru/m_s_tval/n9 [35]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5266 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [34]),
    .c(data_csr[34]),
    .o(_al_u5266_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5267 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[34]),
    .c(wb_exc_code[34]),
    .o(\cu_ru/m_s_tval/n3 [34]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5268 (
    .a(_al_u5157_o),
    .b(_al_u5266_o),
    .c(\cu_ru/m_s_tval/n3 [34]),
    .o(\cu_ru/m_s_tval/n9 [34]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5269 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [33]),
    .c(data_csr[33]),
    .o(_al_u5269_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5270 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[33]),
    .c(wb_exc_code[33]),
    .o(\cu_ru/m_s_tval/n3 [33]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5271 (
    .a(_al_u5157_o),
    .b(_al_u5269_o),
    .c(\cu_ru/m_s_tval/n3 [33]),
    .o(\cu_ru/m_s_tval/n9 [33]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5272 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [32]),
    .c(data_csr[32]),
    .o(_al_u5272_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5273 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[32]),
    .c(wb_exc_code[32]),
    .o(\cu_ru/m_s_tval/n3 [32]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5274 (
    .a(_al_u5157_o),
    .b(_al_u5272_o),
    .c(\cu_ru/m_s_tval/n3 [32]),
    .o(\cu_ru/m_s_tval/n9 [32]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5275 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [31]),
    .c(data_csr[31]),
    .o(_al_u5275_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5276 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[31]),
    .c(wb_exc_code[31]),
    .o(\cu_ru/m_s_tval/n3 [31]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5277 (
    .a(_al_u5157_o),
    .b(_al_u5275_o),
    .c(\cu_ru/m_s_tval/n3 [31]),
    .o(\cu_ru/m_s_tval/n9 [31]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5278 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [30]),
    .c(data_csr[30]),
    .o(_al_u5278_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5279 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[30]),
    .c(wb_exc_code[30]),
    .o(\cu_ru/m_s_tval/n3 [30]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5280 (
    .a(_al_u5157_o),
    .b(_al_u5278_o),
    .c(\cu_ru/m_s_tval/n3 [30]),
    .o(\cu_ru/m_s_tval/n9 [30]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5281 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [3]),
    .c(data_csr[3]),
    .o(_al_u5281_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5282 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[3]),
    .c(wb_exc_code[3]),
    .o(\cu_ru/m_s_tval/n3 [3]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5283 (
    .a(_al_u5157_o),
    .b(_al_u5281_o),
    .c(\cu_ru/m_s_tval/n3 [3]),
    .o(\cu_ru/m_s_tval/n9 [3]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5284 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [29]),
    .c(data_csr[29]),
    .o(_al_u5284_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5285 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[29]),
    .c(wb_exc_code[29]),
    .o(\cu_ru/m_s_tval/n3 [29]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5286 (
    .a(_al_u5157_o),
    .b(_al_u5284_o),
    .c(\cu_ru/m_s_tval/n3 [29]),
    .o(\cu_ru/m_s_tval/n9 [29]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5287 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [28]),
    .c(data_csr[28]),
    .o(_al_u5287_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5288 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[28]),
    .c(wb_exc_code[28]),
    .o(\cu_ru/m_s_tval/n3 [28]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5289 (
    .a(_al_u5157_o),
    .b(_al_u5287_o),
    .c(\cu_ru/m_s_tval/n3 [28]),
    .o(\cu_ru/m_s_tval/n9 [28]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5290 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [27]),
    .c(data_csr[27]),
    .o(_al_u5290_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5291 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[27]),
    .c(wb_exc_code[27]),
    .o(\cu_ru/m_s_tval/n3 [27]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5292 (
    .a(_al_u5157_o),
    .b(_al_u5290_o),
    .c(\cu_ru/m_s_tval/n3 [27]),
    .o(\cu_ru/m_s_tval/n9 [27]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5293 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [26]),
    .c(data_csr[26]),
    .o(_al_u5293_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5294 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[26]),
    .c(wb_exc_code[26]),
    .o(\cu_ru/m_s_tval/n3 [26]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5295 (
    .a(_al_u5157_o),
    .b(_al_u5293_o),
    .c(\cu_ru/m_s_tval/n3 [26]),
    .o(\cu_ru/m_s_tval/n9 [26]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5296 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [25]),
    .c(data_csr[25]),
    .o(_al_u5296_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5297 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[25]),
    .c(wb_exc_code[25]),
    .o(\cu_ru/m_s_tval/n3 [25]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5298 (
    .a(_al_u5157_o),
    .b(_al_u5296_o),
    .c(\cu_ru/m_s_tval/n3 [25]),
    .o(\cu_ru/m_s_tval/n9 [25]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5299 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [24]),
    .c(data_csr[24]),
    .o(_al_u5299_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5300 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[24]),
    .c(wb_exc_code[24]),
    .o(\cu_ru/m_s_tval/n3 [24]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5301 (
    .a(_al_u5157_o),
    .b(_al_u5299_o),
    .c(\cu_ru/m_s_tval/n3 [24]),
    .o(\cu_ru/m_s_tval/n9 [24]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5302 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [23]),
    .c(data_csr[23]),
    .o(_al_u5302_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5303 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[23]),
    .c(wb_exc_code[23]),
    .o(\cu_ru/m_s_tval/n3 [23]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5304 (
    .a(_al_u5157_o),
    .b(_al_u5302_o),
    .c(\cu_ru/m_s_tval/n3 [23]),
    .o(\cu_ru/m_s_tval/n9 [23]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5305 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [22]),
    .c(data_csr[22]),
    .o(_al_u5305_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5306 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[22]),
    .c(wb_exc_code[22]),
    .o(\cu_ru/m_s_tval/n3 [22]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5307 (
    .a(_al_u5157_o),
    .b(_al_u5305_o),
    .c(\cu_ru/m_s_tval/n3 [22]),
    .o(\cu_ru/m_s_tval/n9 [22]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5308 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [21]),
    .c(data_csr[21]),
    .o(_al_u5308_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5309 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[21]),
    .c(wb_exc_code[21]),
    .o(\cu_ru/m_s_tval/n3 [21]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5310 (
    .a(_al_u5157_o),
    .b(_al_u5308_o),
    .c(\cu_ru/m_s_tval/n3 [21]),
    .o(\cu_ru/m_s_tval/n9 [21]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5311 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [20]),
    .c(data_csr[20]),
    .o(_al_u5311_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5312 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[20]),
    .c(wb_exc_code[20]),
    .o(\cu_ru/m_s_tval/n3 [20]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5313 (
    .a(_al_u5157_o),
    .b(_al_u5311_o),
    .c(\cu_ru/m_s_tval/n3 [20]),
    .o(\cu_ru/m_s_tval/n9 [20]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5314 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [2]),
    .c(data_csr[2]),
    .o(_al_u5314_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5315 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[2]),
    .c(wb_exc_code[2]),
    .o(\cu_ru/m_s_tval/n3 [2]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5316 (
    .a(_al_u5157_o),
    .b(_al_u5314_o),
    .c(\cu_ru/m_s_tval/n3 [2]),
    .o(\cu_ru/m_s_tval/n9 [2]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5317 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [19]),
    .c(data_csr[19]),
    .o(_al_u5317_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5318 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[19]),
    .c(wb_exc_code[19]),
    .o(\cu_ru/m_s_tval/n3 [19]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5319 (
    .a(_al_u5157_o),
    .b(_al_u5317_o),
    .c(\cu_ru/m_s_tval/n3 [19]),
    .o(\cu_ru/m_s_tval/n9 [19]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5320 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [18]),
    .c(data_csr[18]),
    .o(_al_u5320_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5321 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[18]),
    .c(wb_exc_code[18]),
    .o(\cu_ru/m_s_tval/n3 [18]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5322 (
    .a(_al_u5157_o),
    .b(_al_u5320_o),
    .c(\cu_ru/m_s_tval/n3 [18]),
    .o(\cu_ru/m_s_tval/n9 [18]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5323 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [17]),
    .c(data_csr[17]),
    .o(_al_u5323_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5324 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[17]),
    .c(wb_exc_code[17]),
    .o(\cu_ru/m_s_tval/n3 [17]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5325 (
    .a(_al_u5157_o),
    .b(_al_u5323_o),
    .c(\cu_ru/m_s_tval/n3 [17]),
    .o(\cu_ru/m_s_tval/n9 [17]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5326 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [16]),
    .c(data_csr[16]),
    .o(_al_u5326_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5327 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[16]),
    .c(wb_exc_code[16]),
    .o(\cu_ru/m_s_tval/n3 [16]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5328 (
    .a(_al_u5157_o),
    .b(_al_u5326_o),
    .c(\cu_ru/m_s_tval/n3 [16]),
    .o(\cu_ru/m_s_tval/n9 [16]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5329 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [15]),
    .c(data_csr[15]),
    .o(_al_u5329_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5330 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[15]),
    .c(wb_exc_code[15]),
    .o(\cu_ru/m_s_tval/n3 [15]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5331 (
    .a(_al_u5157_o),
    .b(_al_u5329_o),
    .c(\cu_ru/m_s_tval/n3 [15]),
    .o(\cu_ru/m_s_tval/n9 [15]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5332 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [14]),
    .c(data_csr[14]),
    .o(_al_u5332_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5333 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[14]),
    .c(wb_exc_code[14]),
    .o(\cu_ru/m_s_tval/n3 [14]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5334 (
    .a(_al_u5157_o),
    .b(_al_u5332_o),
    .c(\cu_ru/m_s_tval/n3 [14]),
    .o(\cu_ru/m_s_tval/n9 [14]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5335 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [13]),
    .c(data_csr[13]),
    .o(_al_u5335_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5336 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[13]),
    .c(wb_exc_code[13]),
    .o(\cu_ru/m_s_tval/n3 [13]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5337 (
    .a(_al_u5157_o),
    .b(_al_u5335_o),
    .c(\cu_ru/m_s_tval/n3 [13]),
    .o(\cu_ru/m_s_tval/n9 [13]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5338 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [12]),
    .c(data_csr[12]),
    .o(_al_u5338_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5339 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[12]),
    .c(wb_exc_code[12]),
    .o(\cu_ru/m_s_tval/n3 [12]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5340 (
    .a(_al_u5157_o),
    .b(_al_u5338_o),
    .c(\cu_ru/m_s_tval/n3 [12]),
    .o(\cu_ru/m_s_tval/n9 [12]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5341 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [11]),
    .c(data_csr[11]),
    .o(_al_u5341_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5342 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[11]),
    .c(wb_exc_code[11]),
    .o(\cu_ru/m_s_tval/n3 [11]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5343 (
    .a(_al_u5157_o),
    .b(_al_u5341_o),
    .c(\cu_ru/m_s_tval/n3 [11]),
    .o(\cu_ru/m_s_tval/n9 [11]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5344 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [10]),
    .c(data_csr[10]),
    .o(_al_u5344_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5345 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[10]),
    .c(wb_exc_code[10]),
    .o(\cu_ru/m_s_tval/n3 [10]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5346 (
    .a(_al_u5157_o),
    .b(_al_u5344_o),
    .c(\cu_ru/m_s_tval/n3 [10]),
    .o(\cu_ru/m_s_tval/n9 [10]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5347 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [1]),
    .c(data_csr[1]),
    .o(_al_u5347_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5348 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[1]),
    .c(wb_exc_code[1]),
    .o(\cu_ru/m_s_tval/n3 [1]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5349 (
    .a(_al_u5157_o),
    .b(_al_u5347_o),
    .c(\cu_ru/m_s_tval/n3 [1]),
    .o(\cu_ru/m_s_tval/n9 [1]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5350 (
    .a(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .b(\cu_ru/stval [0]),
    .c(data_csr[0]),
    .o(_al_u5350_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u5351 (
    .a(_al_u5161_o),
    .b(wb_ins_pc[0]),
    .c(wb_exc_code[0]),
    .o(\cu_ru/m_s_tval/n3 [0]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5352 (
    .a(_al_u5157_o),
    .b(_al_u5350_o),
    .c(\cu_ru/m_s_tval/n3 [0]),
    .o(\cu_ru/m_s_tval/n9 [0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5353 (
    .a(int_req),
    .b(wb_ebreak),
    .o(_al_u5353_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5354 (
    .a(\cu_ru/m_s_epc/n0 [7]),
    .b(pc_jmp),
    .c(new_pc[9]),
    .o(_al_u5354_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5355 (
    .a(_al_u5353_o),
    .b(_al_u5354_o),
    .c(wb_ins_pc[9]),
    .o(\cu_ru/m_s_epc/n2 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u5356 (
    .a(_al_u5158_o),
    .b(_al_u3200_o),
    .c(csr_index[1]),
    .d(csr_index[2]),
    .o(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5357 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [9]),
    .c(data_csr[9]),
    .o(_al_u5357_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5358 (
    .a(\cu_ru/m_s_epc/n2 [9]),
    .b(_al_u5157_o),
    .c(_al_u5357_o),
    .o(\cu_ru/m_s_epc/n8 [9]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5359 (
    .a(\cu_ru/m_s_epc/n0 [6]),
    .b(pc_jmp),
    .c(new_pc[8]),
    .o(_al_u5359_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5360 (
    .a(_al_u5353_o),
    .b(_al_u5359_o),
    .c(wb_ins_pc[8]),
    .o(\cu_ru/m_s_epc/n2 [8]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5361 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [8]),
    .c(data_csr[8]),
    .o(_al_u5361_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5362 (
    .a(\cu_ru/m_s_epc/n2 [8]),
    .b(_al_u5157_o),
    .c(_al_u5361_o),
    .o(\cu_ru/m_s_epc/n8 [8]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5363 (
    .a(\cu_ru/m_s_epc/n0 [5]),
    .b(pc_jmp),
    .c(new_pc[7]),
    .o(_al_u5363_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5364 (
    .a(_al_u5353_o),
    .b(_al_u5363_o),
    .c(wb_ins_pc[7]),
    .o(\cu_ru/m_s_epc/n2 [7]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5365 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [7]),
    .c(data_csr[7]),
    .o(_al_u5365_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5366 (
    .a(\cu_ru/m_s_epc/n2 [7]),
    .b(_al_u5157_o),
    .c(_al_u5365_o),
    .o(\cu_ru/m_s_epc/n8 [7]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5367 (
    .a(\cu_ru/m_s_epc/n0 [61]),
    .b(pc_jmp),
    .c(new_pc[63]),
    .o(_al_u5367_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5368 (
    .a(_al_u5353_o),
    .b(_al_u5367_o),
    .c(wb_ins_pc[63]),
    .o(\cu_ru/m_s_epc/n2 [63]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5369 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [63]),
    .c(data_csr[63]),
    .o(_al_u5369_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5370 (
    .a(\cu_ru/m_s_epc/n2 [63]),
    .b(_al_u5157_o),
    .c(_al_u5369_o),
    .o(\cu_ru/m_s_epc/n8 [63]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5371 (
    .a(\cu_ru/m_s_epc/n0 [60]),
    .b(pc_jmp),
    .c(new_pc[62]),
    .o(_al_u5371_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5372 (
    .a(_al_u5353_o),
    .b(_al_u5371_o),
    .c(wb_ins_pc[62]),
    .o(\cu_ru/m_s_epc/n2 [62]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5373 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [62]),
    .c(data_csr[62]),
    .o(_al_u5373_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5374 (
    .a(\cu_ru/m_s_epc/n2 [62]),
    .b(_al_u5157_o),
    .c(_al_u5373_o),
    .o(\cu_ru/m_s_epc/n8 [62]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5375 (
    .a(\cu_ru/m_s_epc/n0 [59]),
    .b(pc_jmp),
    .c(new_pc[61]),
    .o(_al_u5375_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5376 (
    .a(_al_u5353_o),
    .b(_al_u5375_o),
    .c(wb_ins_pc[61]),
    .o(\cu_ru/m_s_epc/n2 [61]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5377 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [61]),
    .c(data_csr[61]),
    .o(_al_u5377_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5378 (
    .a(\cu_ru/m_s_epc/n2 [61]),
    .b(_al_u5157_o),
    .c(_al_u5377_o),
    .o(\cu_ru/m_s_epc/n8 [61]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5379 (
    .a(\cu_ru/m_s_epc/n0 [58]),
    .b(pc_jmp),
    .c(new_pc[60]),
    .o(_al_u5379_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5380 (
    .a(_al_u5353_o),
    .b(_al_u5379_o),
    .c(wb_ins_pc[60]),
    .o(\cu_ru/m_s_epc/n2 [60]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5381 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [60]),
    .c(data_csr[60]),
    .o(_al_u5381_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5382 (
    .a(\cu_ru/m_s_epc/n2 [60]),
    .b(_al_u5157_o),
    .c(_al_u5381_o),
    .o(\cu_ru/m_s_epc/n8 [60]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5383 (
    .a(\cu_ru/m_s_epc/n0 [4]),
    .b(pc_jmp),
    .c(new_pc[6]),
    .o(_al_u5383_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5384 (
    .a(_al_u5353_o),
    .b(_al_u5383_o),
    .c(wb_ins_pc[6]),
    .o(\cu_ru/m_s_epc/n2 [6]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5385 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [6]),
    .c(data_csr[6]),
    .o(_al_u5385_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5386 (
    .a(\cu_ru/m_s_epc/n2 [6]),
    .b(_al_u5157_o),
    .c(_al_u5385_o),
    .o(\cu_ru/m_s_epc/n8 [6]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5387 (
    .a(\cu_ru/m_s_epc/n0 [57]),
    .b(pc_jmp),
    .c(new_pc[59]),
    .o(_al_u5387_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5388 (
    .a(_al_u5353_o),
    .b(_al_u5387_o),
    .c(wb_ins_pc[59]),
    .o(\cu_ru/m_s_epc/n2 [59]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5389 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [59]),
    .c(data_csr[59]),
    .o(_al_u5389_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5390 (
    .a(\cu_ru/m_s_epc/n2 [59]),
    .b(_al_u5157_o),
    .c(_al_u5389_o),
    .o(\cu_ru/m_s_epc/n8 [59]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5391 (
    .a(\cu_ru/m_s_epc/n0 [56]),
    .b(pc_jmp),
    .c(new_pc[58]),
    .o(_al_u5391_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5392 (
    .a(_al_u5353_o),
    .b(_al_u5391_o),
    .c(wb_ins_pc[58]),
    .o(\cu_ru/m_s_epc/n2 [58]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5393 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [58]),
    .c(data_csr[58]),
    .o(_al_u5393_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5394 (
    .a(\cu_ru/m_s_epc/n2 [58]),
    .b(_al_u5157_o),
    .c(_al_u5393_o),
    .o(\cu_ru/m_s_epc/n8 [58]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5395 (
    .a(\cu_ru/m_s_epc/n0 [55]),
    .b(pc_jmp),
    .c(new_pc[57]),
    .o(_al_u5395_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5396 (
    .a(_al_u5353_o),
    .b(_al_u5395_o),
    .c(wb_ins_pc[57]),
    .o(\cu_ru/m_s_epc/n2 [57]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5397 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [57]),
    .c(data_csr[57]),
    .o(_al_u5397_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5398 (
    .a(\cu_ru/m_s_epc/n2 [57]),
    .b(_al_u5157_o),
    .c(_al_u5397_o),
    .o(\cu_ru/m_s_epc/n8 [57]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5399 (
    .a(\cu_ru/m_s_epc/n0 [54]),
    .b(pc_jmp),
    .c(new_pc[56]),
    .o(_al_u5399_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5400 (
    .a(_al_u5353_o),
    .b(_al_u5399_o),
    .c(wb_ins_pc[56]),
    .o(\cu_ru/m_s_epc/n2 [56]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5401 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [56]),
    .c(data_csr[56]),
    .o(_al_u5401_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5402 (
    .a(\cu_ru/m_s_epc/n2 [56]),
    .b(_al_u5157_o),
    .c(_al_u5401_o),
    .o(\cu_ru/m_s_epc/n8 [56]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5403 (
    .a(\cu_ru/m_s_epc/n0 [53]),
    .b(pc_jmp),
    .c(new_pc[55]),
    .o(_al_u5403_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5404 (
    .a(_al_u5353_o),
    .b(_al_u5403_o),
    .c(wb_ins_pc[55]),
    .o(\cu_ru/m_s_epc/n2 [55]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5405 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [55]),
    .c(data_csr[55]),
    .o(_al_u5405_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5406 (
    .a(\cu_ru/m_s_epc/n2 [55]),
    .b(_al_u5157_o),
    .c(_al_u5405_o),
    .o(\cu_ru/m_s_epc/n8 [55]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5407 (
    .a(\cu_ru/m_s_epc/n0 [52]),
    .b(pc_jmp),
    .c(new_pc[54]),
    .o(_al_u5407_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5408 (
    .a(_al_u5353_o),
    .b(_al_u5407_o),
    .c(wb_ins_pc[54]),
    .o(\cu_ru/m_s_epc/n2 [54]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5409 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [54]),
    .c(data_csr[54]),
    .o(_al_u5409_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5410 (
    .a(\cu_ru/m_s_epc/n2 [54]),
    .b(_al_u5157_o),
    .c(_al_u5409_o),
    .o(\cu_ru/m_s_epc/n8 [54]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5411 (
    .a(\cu_ru/m_s_epc/n0 [51]),
    .b(pc_jmp),
    .c(new_pc[53]),
    .o(_al_u5411_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5412 (
    .a(_al_u5353_o),
    .b(_al_u5411_o),
    .c(wb_ins_pc[53]),
    .o(\cu_ru/m_s_epc/n2 [53]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5413 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [53]),
    .c(data_csr[53]),
    .o(_al_u5413_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5414 (
    .a(\cu_ru/m_s_epc/n2 [53]),
    .b(_al_u5157_o),
    .c(_al_u5413_o),
    .o(\cu_ru/m_s_epc/n8 [53]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5415 (
    .a(\cu_ru/m_s_epc/n0 [50]),
    .b(pc_jmp),
    .c(new_pc[52]),
    .o(_al_u5415_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5416 (
    .a(_al_u5353_o),
    .b(_al_u5415_o),
    .c(wb_ins_pc[52]),
    .o(\cu_ru/m_s_epc/n2 [52]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5417 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [52]),
    .c(data_csr[52]),
    .o(_al_u5417_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5418 (
    .a(\cu_ru/m_s_epc/n2 [52]),
    .b(_al_u5157_o),
    .c(_al_u5417_o),
    .o(\cu_ru/m_s_epc/n8 [52]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5419 (
    .a(\cu_ru/m_s_epc/n0 [49]),
    .b(pc_jmp),
    .c(new_pc[51]),
    .o(_al_u5419_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5420 (
    .a(_al_u5353_o),
    .b(_al_u5419_o),
    .c(wb_ins_pc[51]),
    .o(\cu_ru/m_s_epc/n2 [51]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5421 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [51]),
    .c(data_csr[51]),
    .o(_al_u5421_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5422 (
    .a(\cu_ru/m_s_epc/n2 [51]),
    .b(_al_u5157_o),
    .c(_al_u5421_o),
    .o(\cu_ru/m_s_epc/n8 [51]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5423 (
    .a(\cu_ru/m_s_epc/n0 [48]),
    .b(pc_jmp),
    .c(new_pc[50]),
    .o(_al_u5423_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5424 (
    .a(_al_u5353_o),
    .b(_al_u5423_o),
    .c(wb_ins_pc[50]),
    .o(\cu_ru/m_s_epc/n2 [50]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5425 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [50]),
    .c(data_csr[50]),
    .o(_al_u5425_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5426 (
    .a(\cu_ru/m_s_epc/n2 [50]),
    .b(_al_u5157_o),
    .c(_al_u5425_o),
    .o(\cu_ru/m_s_epc/n8 [50]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5427 (
    .a(\cu_ru/m_s_epc/n0 [3]),
    .b(pc_jmp),
    .c(new_pc[5]),
    .o(_al_u5427_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5428 (
    .a(_al_u5353_o),
    .b(_al_u5427_o),
    .c(wb_ins_pc[5]),
    .o(\cu_ru/m_s_epc/n2 [5]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5429 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [5]),
    .c(data_csr[5]),
    .o(_al_u5429_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5430 (
    .a(\cu_ru/m_s_epc/n2 [5]),
    .b(_al_u5157_o),
    .c(_al_u5429_o),
    .o(\cu_ru/m_s_epc/n8 [5]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5431 (
    .a(\cu_ru/m_s_epc/n0 [47]),
    .b(pc_jmp),
    .c(new_pc[49]),
    .o(_al_u5431_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5432 (
    .a(_al_u5353_o),
    .b(_al_u5431_o),
    .c(wb_ins_pc[49]),
    .o(\cu_ru/m_s_epc/n2 [49]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5433 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [49]),
    .c(data_csr[49]),
    .o(_al_u5433_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5434 (
    .a(\cu_ru/m_s_epc/n2 [49]),
    .b(_al_u5157_o),
    .c(_al_u5433_o),
    .o(\cu_ru/m_s_epc/n8 [49]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5435 (
    .a(\cu_ru/m_s_epc/n0 [46]),
    .b(pc_jmp),
    .c(new_pc[48]),
    .o(_al_u5435_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5436 (
    .a(_al_u5353_o),
    .b(_al_u5435_o),
    .c(wb_ins_pc[48]),
    .o(\cu_ru/m_s_epc/n2 [48]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5437 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [48]),
    .c(data_csr[48]),
    .o(_al_u5437_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5438 (
    .a(\cu_ru/m_s_epc/n2 [48]),
    .b(_al_u5157_o),
    .c(_al_u5437_o),
    .o(\cu_ru/m_s_epc/n8 [48]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5439 (
    .a(\cu_ru/m_s_epc/n0 [45]),
    .b(pc_jmp),
    .c(new_pc[47]),
    .o(_al_u5439_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5440 (
    .a(_al_u5353_o),
    .b(_al_u5439_o),
    .c(wb_ins_pc[47]),
    .o(\cu_ru/m_s_epc/n2 [47]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5441 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [47]),
    .c(data_csr[47]),
    .o(_al_u5441_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5442 (
    .a(\cu_ru/m_s_epc/n2 [47]),
    .b(_al_u5157_o),
    .c(_al_u5441_o),
    .o(\cu_ru/m_s_epc/n8 [47]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5443 (
    .a(\cu_ru/m_s_epc/n0 [44]),
    .b(pc_jmp),
    .c(new_pc[46]),
    .o(_al_u5443_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5444 (
    .a(_al_u5353_o),
    .b(_al_u5443_o),
    .c(wb_ins_pc[46]),
    .o(\cu_ru/m_s_epc/n2 [46]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5445 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [46]),
    .c(data_csr[46]),
    .o(_al_u5445_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5446 (
    .a(\cu_ru/m_s_epc/n2 [46]),
    .b(_al_u5157_o),
    .c(_al_u5445_o),
    .o(\cu_ru/m_s_epc/n8 [46]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5447 (
    .a(\cu_ru/m_s_epc/n0 [43]),
    .b(pc_jmp),
    .c(new_pc[45]),
    .o(_al_u5447_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5448 (
    .a(_al_u5353_o),
    .b(_al_u5447_o),
    .c(wb_ins_pc[45]),
    .o(\cu_ru/m_s_epc/n2 [45]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5449 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [45]),
    .c(data_csr[45]),
    .o(_al_u5449_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5450 (
    .a(\cu_ru/m_s_epc/n2 [45]),
    .b(_al_u5157_o),
    .c(_al_u5449_o),
    .o(\cu_ru/m_s_epc/n8 [45]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5451 (
    .a(\cu_ru/m_s_epc/n0 [42]),
    .b(pc_jmp),
    .c(new_pc[44]),
    .o(_al_u5451_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5452 (
    .a(_al_u5353_o),
    .b(_al_u5451_o),
    .c(wb_ins_pc[44]),
    .o(\cu_ru/m_s_epc/n2 [44]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5453 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [44]),
    .c(data_csr[44]),
    .o(_al_u5453_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5454 (
    .a(\cu_ru/m_s_epc/n2 [44]),
    .b(_al_u5157_o),
    .c(_al_u5453_o),
    .o(\cu_ru/m_s_epc/n8 [44]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5455 (
    .a(\cu_ru/m_s_epc/n0 [41]),
    .b(pc_jmp),
    .c(new_pc[43]),
    .o(_al_u5455_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5456 (
    .a(_al_u5353_o),
    .b(_al_u5455_o),
    .c(wb_ins_pc[43]),
    .o(\cu_ru/m_s_epc/n2 [43]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5457 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [43]),
    .c(data_csr[43]),
    .o(_al_u5457_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5458 (
    .a(\cu_ru/m_s_epc/n2 [43]),
    .b(_al_u5157_o),
    .c(_al_u5457_o),
    .o(\cu_ru/m_s_epc/n8 [43]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5459 (
    .a(\cu_ru/m_s_epc/n0 [40]),
    .b(pc_jmp),
    .c(new_pc[42]),
    .o(_al_u5459_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5460 (
    .a(_al_u5353_o),
    .b(_al_u5459_o),
    .c(wb_ins_pc[42]),
    .o(\cu_ru/m_s_epc/n2 [42]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5461 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [42]),
    .c(data_csr[42]),
    .o(_al_u5461_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5462 (
    .a(\cu_ru/m_s_epc/n2 [42]),
    .b(_al_u5157_o),
    .c(_al_u5461_o),
    .o(\cu_ru/m_s_epc/n8 [42]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5463 (
    .a(\cu_ru/m_s_epc/n0 [39]),
    .b(pc_jmp),
    .c(new_pc[41]),
    .o(_al_u5463_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5464 (
    .a(_al_u5353_o),
    .b(_al_u5463_o),
    .c(wb_ins_pc[41]),
    .o(\cu_ru/m_s_epc/n2 [41]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5465 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [41]),
    .c(data_csr[41]),
    .o(_al_u5465_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5466 (
    .a(\cu_ru/m_s_epc/n2 [41]),
    .b(_al_u5157_o),
    .c(_al_u5465_o),
    .o(\cu_ru/m_s_epc/n8 [41]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5467 (
    .a(\cu_ru/m_s_epc/n0 [38]),
    .b(pc_jmp),
    .c(new_pc[40]),
    .o(_al_u5467_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5468 (
    .a(_al_u5353_o),
    .b(_al_u5467_o),
    .c(wb_ins_pc[40]),
    .o(\cu_ru/m_s_epc/n2 [40]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5469 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [40]),
    .c(data_csr[40]),
    .o(_al_u5469_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5470 (
    .a(\cu_ru/m_s_epc/n2 [40]),
    .b(_al_u5157_o),
    .c(_al_u5469_o),
    .o(\cu_ru/m_s_epc/n8 [40]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5471 (
    .a(\cu_ru/m_s_epc/n0 [2]),
    .b(pc_jmp),
    .c(new_pc[4]),
    .o(_al_u5471_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5472 (
    .a(_al_u5353_o),
    .b(_al_u5471_o),
    .c(wb_ins_pc[4]),
    .o(\cu_ru/m_s_epc/n2 [4]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5473 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [4]),
    .c(data_csr[4]),
    .o(_al_u5473_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5474 (
    .a(\cu_ru/m_s_epc/n2 [4]),
    .b(_al_u5157_o),
    .c(_al_u5473_o),
    .o(\cu_ru/m_s_epc/n8 [4]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5475 (
    .a(\cu_ru/m_s_epc/n0 [37]),
    .b(pc_jmp),
    .c(new_pc[39]),
    .o(_al_u5475_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5476 (
    .a(_al_u5353_o),
    .b(_al_u5475_o),
    .c(wb_ins_pc[39]),
    .o(\cu_ru/m_s_epc/n2 [39]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5477 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [39]),
    .c(data_csr[39]),
    .o(_al_u5477_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5478 (
    .a(\cu_ru/m_s_epc/n2 [39]),
    .b(_al_u5157_o),
    .c(_al_u5477_o),
    .o(\cu_ru/m_s_epc/n8 [39]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5479 (
    .a(\cu_ru/m_s_epc/n0 [36]),
    .b(pc_jmp),
    .c(new_pc[38]),
    .o(_al_u5479_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5480 (
    .a(_al_u5353_o),
    .b(_al_u5479_o),
    .c(wb_ins_pc[38]),
    .o(\cu_ru/m_s_epc/n2 [38]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5481 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [38]),
    .c(data_csr[38]),
    .o(_al_u5481_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5482 (
    .a(\cu_ru/m_s_epc/n2 [38]),
    .b(_al_u5157_o),
    .c(_al_u5481_o),
    .o(\cu_ru/m_s_epc/n8 [38]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5483 (
    .a(\cu_ru/m_s_epc/n0 [35]),
    .b(pc_jmp),
    .c(new_pc[37]),
    .o(_al_u5483_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5484 (
    .a(_al_u5353_o),
    .b(_al_u5483_o),
    .c(wb_ins_pc[37]),
    .o(\cu_ru/m_s_epc/n2 [37]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5485 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [37]),
    .c(data_csr[37]),
    .o(_al_u5485_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5486 (
    .a(\cu_ru/m_s_epc/n2 [37]),
    .b(_al_u5157_o),
    .c(_al_u5485_o),
    .o(\cu_ru/m_s_epc/n8 [37]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5487 (
    .a(\cu_ru/m_s_epc/n0 [34]),
    .b(pc_jmp),
    .c(new_pc[36]),
    .o(_al_u5487_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5488 (
    .a(_al_u5353_o),
    .b(_al_u5487_o),
    .c(wb_ins_pc[36]),
    .o(\cu_ru/m_s_epc/n2 [36]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5489 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [36]),
    .c(data_csr[36]),
    .o(_al_u5489_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5490 (
    .a(\cu_ru/m_s_epc/n2 [36]),
    .b(_al_u5157_o),
    .c(_al_u5489_o),
    .o(\cu_ru/m_s_epc/n8 [36]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5491 (
    .a(\cu_ru/m_s_epc/n0 [33]),
    .b(pc_jmp),
    .c(new_pc[35]),
    .o(_al_u5491_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5492 (
    .a(_al_u5353_o),
    .b(_al_u5491_o),
    .c(wb_ins_pc[35]),
    .o(\cu_ru/m_s_epc/n2 [35]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5493 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [35]),
    .c(data_csr[35]),
    .o(_al_u5493_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5494 (
    .a(\cu_ru/m_s_epc/n2 [35]),
    .b(_al_u5157_o),
    .c(_al_u5493_o),
    .o(\cu_ru/m_s_epc/n8 [35]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5495 (
    .a(\cu_ru/m_s_epc/n0 [32]),
    .b(pc_jmp),
    .c(new_pc[34]),
    .o(_al_u5495_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5496 (
    .a(_al_u5353_o),
    .b(_al_u5495_o),
    .c(wb_ins_pc[34]),
    .o(\cu_ru/m_s_epc/n2 [34]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5497 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [34]),
    .c(data_csr[34]),
    .o(_al_u5497_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5498 (
    .a(\cu_ru/m_s_epc/n2 [34]),
    .b(_al_u5157_o),
    .c(_al_u5497_o),
    .o(\cu_ru/m_s_epc/n8 [34]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5499 (
    .a(\cu_ru/m_s_epc/n0 [31]),
    .b(pc_jmp),
    .c(new_pc[33]),
    .o(_al_u5499_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5500 (
    .a(_al_u5353_o),
    .b(_al_u5499_o),
    .c(wb_ins_pc[33]),
    .o(\cu_ru/m_s_epc/n2 [33]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5501 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [33]),
    .c(data_csr[33]),
    .o(_al_u5501_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5502 (
    .a(\cu_ru/m_s_epc/n2 [33]),
    .b(_al_u5157_o),
    .c(_al_u5501_o),
    .o(\cu_ru/m_s_epc/n8 [33]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5503 (
    .a(\cu_ru/m_s_epc/n0 [30]),
    .b(pc_jmp),
    .c(new_pc[32]),
    .o(_al_u5503_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5504 (
    .a(_al_u5353_o),
    .b(_al_u5503_o),
    .c(wb_ins_pc[32]),
    .o(\cu_ru/m_s_epc/n2 [32]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5505 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [32]),
    .c(data_csr[32]),
    .o(_al_u5505_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5506 (
    .a(\cu_ru/m_s_epc/n2 [32]),
    .b(_al_u5157_o),
    .c(_al_u5505_o),
    .o(\cu_ru/m_s_epc/n8 [32]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5507 (
    .a(\cu_ru/m_s_epc/n0 [29]),
    .b(pc_jmp),
    .c(new_pc[31]),
    .o(_al_u5507_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5508 (
    .a(_al_u5353_o),
    .b(_al_u5507_o),
    .c(wb_ins_pc[31]),
    .o(\cu_ru/m_s_epc/n2 [31]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5509 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [31]),
    .c(data_csr[31]),
    .o(_al_u5509_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5510 (
    .a(\cu_ru/m_s_epc/n2 [31]),
    .b(_al_u5157_o),
    .c(_al_u5509_o),
    .o(\cu_ru/m_s_epc/n8 [31]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5511 (
    .a(\cu_ru/m_s_epc/n0 [28]),
    .b(pc_jmp),
    .c(new_pc[30]),
    .o(_al_u5511_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5512 (
    .a(_al_u5353_o),
    .b(_al_u5511_o),
    .c(wb_ins_pc[30]),
    .o(\cu_ru/m_s_epc/n2 [30]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5513 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [30]),
    .c(data_csr[30]),
    .o(_al_u5513_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5514 (
    .a(\cu_ru/m_s_epc/n2 [30]),
    .b(_al_u5157_o),
    .c(_al_u5513_o),
    .o(\cu_ru/m_s_epc/n8 [30]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5515 (
    .a(\cu_ru/m_s_epc/n0 [1]),
    .b(pc_jmp),
    .c(new_pc[3]),
    .o(_al_u5515_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5516 (
    .a(_al_u5353_o),
    .b(_al_u5515_o),
    .c(wb_ins_pc[3]),
    .o(\cu_ru/m_s_epc/n2 [3]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5517 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [3]),
    .c(data_csr[3]),
    .o(_al_u5517_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5518 (
    .a(\cu_ru/m_s_epc/n2 [3]),
    .b(_al_u5157_o),
    .c(_al_u5517_o),
    .o(\cu_ru/m_s_epc/n8 [3]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5519 (
    .a(\cu_ru/m_s_epc/n0 [27]),
    .b(pc_jmp),
    .c(new_pc[29]),
    .o(_al_u5519_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5520 (
    .a(_al_u5353_o),
    .b(_al_u5519_o),
    .c(wb_ins_pc[29]),
    .o(\cu_ru/m_s_epc/n2 [29]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5521 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [29]),
    .c(data_csr[29]),
    .o(_al_u5521_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5522 (
    .a(\cu_ru/m_s_epc/n2 [29]),
    .b(_al_u5157_o),
    .c(_al_u5521_o),
    .o(\cu_ru/m_s_epc/n8 [29]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5523 (
    .a(\cu_ru/m_s_epc/n0 [26]),
    .b(pc_jmp),
    .c(new_pc[28]),
    .o(_al_u5523_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5524 (
    .a(_al_u5353_o),
    .b(_al_u5523_o),
    .c(wb_ins_pc[28]),
    .o(\cu_ru/m_s_epc/n2 [28]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5525 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [28]),
    .c(data_csr[28]),
    .o(_al_u5525_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5526 (
    .a(\cu_ru/m_s_epc/n2 [28]),
    .b(_al_u5157_o),
    .c(_al_u5525_o),
    .o(\cu_ru/m_s_epc/n8 [28]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5527 (
    .a(\cu_ru/m_s_epc/n0 [25]),
    .b(pc_jmp),
    .c(new_pc[27]),
    .o(_al_u5527_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5528 (
    .a(_al_u5353_o),
    .b(_al_u5527_o),
    .c(wb_ins_pc[27]),
    .o(\cu_ru/m_s_epc/n2 [27]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5529 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [27]),
    .c(data_csr[27]),
    .o(_al_u5529_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5530 (
    .a(\cu_ru/m_s_epc/n2 [27]),
    .b(_al_u5157_o),
    .c(_al_u5529_o),
    .o(\cu_ru/m_s_epc/n8 [27]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5531 (
    .a(\cu_ru/m_s_epc/n0 [24]),
    .b(pc_jmp),
    .c(new_pc[26]),
    .o(_al_u5531_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5532 (
    .a(_al_u5353_o),
    .b(_al_u5531_o),
    .c(wb_ins_pc[26]),
    .o(\cu_ru/m_s_epc/n2 [26]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5533 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [26]),
    .c(data_csr[26]),
    .o(_al_u5533_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5534 (
    .a(\cu_ru/m_s_epc/n2 [26]),
    .b(_al_u5157_o),
    .c(_al_u5533_o),
    .o(\cu_ru/m_s_epc/n8 [26]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5535 (
    .a(\cu_ru/m_s_epc/n0 [23]),
    .b(pc_jmp),
    .c(new_pc[25]),
    .o(_al_u5535_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5536 (
    .a(_al_u5353_o),
    .b(_al_u5535_o),
    .c(wb_ins_pc[25]),
    .o(\cu_ru/m_s_epc/n2 [25]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5537 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [25]),
    .c(data_csr[25]),
    .o(_al_u5537_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5538 (
    .a(\cu_ru/m_s_epc/n2 [25]),
    .b(_al_u5157_o),
    .c(_al_u5537_o),
    .o(\cu_ru/m_s_epc/n8 [25]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5539 (
    .a(\cu_ru/m_s_epc/n0 [22]),
    .b(pc_jmp),
    .c(new_pc[24]),
    .o(_al_u5539_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5540 (
    .a(_al_u5353_o),
    .b(_al_u5539_o),
    .c(wb_ins_pc[24]),
    .o(\cu_ru/m_s_epc/n2 [24]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5541 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [24]),
    .c(data_csr[24]),
    .o(_al_u5541_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5542 (
    .a(\cu_ru/m_s_epc/n2 [24]),
    .b(_al_u5157_o),
    .c(_al_u5541_o),
    .o(\cu_ru/m_s_epc/n8 [24]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5543 (
    .a(\cu_ru/m_s_epc/n0 [21]),
    .b(pc_jmp),
    .c(new_pc[23]),
    .o(_al_u5543_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5544 (
    .a(_al_u5353_o),
    .b(_al_u5543_o),
    .c(wb_ins_pc[23]),
    .o(\cu_ru/m_s_epc/n2 [23]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5545 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [23]),
    .c(data_csr[23]),
    .o(_al_u5545_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5546 (
    .a(\cu_ru/m_s_epc/n2 [23]),
    .b(_al_u5157_o),
    .c(_al_u5545_o),
    .o(\cu_ru/m_s_epc/n8 [23]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5547 (
    .a(\cu_ru/m_s_epc/n0 [20]),
    .b(pc_jmp),
    .c(new_pc[22]),
    .o(_al_u5547_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5548 (
    .a(_al_u5353_o),
    .b(_al_u5547_o),
    .c(wb_ins_pc[22]),
    .o(\cu_ru/m_s_epc/n2 [22]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5549 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [22]),
    .c(data_csr[22]),
    .o(_al_u5549_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5550 (
    .a(\cu_ru/m_s_epc/n2 [22]),
    .b(_al_u5157_o),
    .c(_al_u5549_o),
    .o(\cu_ru/m_s_epc/n8 [22]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5551 (
    .a(\cu_ru/m_s_epc/n0 [19]),
    .b(pc_jmp),
    .c(new_pc[21]),
    .o(_al_u5551_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5552 (
    .a(_al_u5353_o),
    .b(_al_u5551_o),
    .c(wb_ins_pc[21]),
    .o(\cu_ru/m_s_epc/n2 [21]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5553 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [21]),
    .c(data_csr[21]),
    .o(_al_u5553_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5554 (
    .a(\cu_ru/m_s_epc/n2 [21]),
    .b(_al_u5157_o),
    .c(_al_u5553_o),
    .o(\cu_ru/m_s_epc/n8 [21]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5555 (
    .a(\cu_ru/m_s_epc/n0 [18]),
    .b(pc_jmp),
    .c(new_pc[20]),
    .o(_al_u5555_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5556 (
    .a(_al_u5353_o),
    .b(_al_u5555_o),
    .c(wb_ins_pc[20]),
    .o(\cu_ru/m_s_epc/n2 [20]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5557 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [20]),
    .c(data_csr[20]),
    .o(_al_u5557_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5558 (
    .a(\cu_ru/m_s_epc/n2 [20]),
    .b(_al_u5157_o),
    .c(_al_u5557_o),
    .o(\cu_ru/m_s_epc/n8 [20]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5559 (
    .a(\cu_ru/m_s_epc/n0 [0]),
    .b(pc_jmp),
    .c(new_pc[2]),
    .o(_al_u5559_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5560 (
    .a(_al_u5353_o),
    .b(_al_u5559_o),
    .c(wb_ins_pc[2]),
    .o(\cu_ru/m_s_epc/n2 [2]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5561 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [2]),
    .c(data_csr[2]),
    .o(_al_u5561_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5562 (
    .a(\cu_ru/m_s_epc/n2 [2]),
    .b(_al_u5157_o),
    .c(_al_u5561_o),
    .o(\cu_ru/m_s_epc/n8 [2]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5563 (
    .a(\cu_ru/m_s_epc/n0 [17]),
    .b(pc_jmp),
    .c(new_pc[19]),
    .o(_al_u5563_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5564 (
    .a(_al_u5353_o),
    .b(_al_u5563_o),
    .c(wb_ins_pc[19]),
    .o(\cu_ru/m_s_epc/n2 [19]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5565 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [19]),
    .c(data_csr[19]),
    .o(_al_u5565_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5566 (
    .a(\cu_ru/m_s_epc/n2 [19]),
    .b(_al_u5157_o),
    .c(_al_u5565_o),
    .o(\cu_ru/m_s_epc/n8 [19]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5567 (
    .a(\cu_ru/m_s_epc/n0 [16]),
    .b(pc_jmp),
    .c(new_pc[18]),
    .o(_al_u5567_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5568 (
    .a(_al_u5353_o),
    .b(_al_u5567_o),
    .c(wb_ins_pc[18]),
    .o(\cu_ru/m_s_epc/n2 [18]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5569 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [18]),
    .c(data_csr[18]),
    .o(_al_u5569_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5570 (
    .a(\cu_ru/m_s_epc/n2 [18]),
    .b(_al_u5157_o),
    .c(_al_u5569_o),
    .o(\cu_ru/m_s_epc/n8 [18]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5571 (
    .a(\cu_ru/m_s_epc/n0 [15]),
    .b(pc_jmp),
    .c(new_pc[17]),
    .o(_al_u5571_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5572 (
    .a(_al_u5353_o),
    .b(_al_u5571_o),
    .c(wb_ins_pc[17]),
    .o(\cu_ru/m_s_epc/n2 [17]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5573 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [17]),
    .c(data_csr[17]),
    .o(_al_u5573_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5574 (
    .a(\cu_ru/m_s_epc/n2 [17]),
    .b(_al_u5157_o),
    .c(_al_u5573_o),
    .o(\cu_ru/m_s_epc/n8 [17]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5575 (
    .a(\cu_ru/m_s_epc/n0 [14]),
    .b(pc_jmp),
    .c(new_pc[16]),
    .o(_al_u5575_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5576 (
    .a(_al_u5353_o),
    .b(_al_u5575_o),
    .c(wb_ins_pc[16]),
    .o(\cu_ru/m_s_epc/n2 [16]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5577 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [16]),
    .c(data_csr[16]),
    .o(_al_u5577_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5578 (
    .a(\cu_ru/m_s_epc/n2 [16]),
    .b(_al_u5157_o),
    .c(_al_u5577_o),
    .o(\cu_ru/m_s_epc/n8 [16]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5579 (
    .a(\cu_ru/m_s_epc/n0 [13]),
    .b(pc_jmp),
    .c(new_pc[15]),
    .o(_al_u5579_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5580 (
    .a(_al_u5353_o),
    .b(_al_u5579_o),
    .c(wb_ins_pc[15]),
    .o(\cu_ru/m_s_epc/n2 [15]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5581 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [15]),
    .c(data_csr[15]),
    .o(_al_u5581_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5582 (
    .a(\cu_ru/m_s_epc/n2 [15]),
    .b(_al_u5157_o),
    .c(_al_u5581_o),
    .o(\cu_ru/m_s_epc/n8 [15]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5583 (
    .a(\cu_ru/m_s_epc/n0 [12]),
    .b(pc_jmp),
    .c(new_pc[14]),
    .o(_al_u5583_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5584 (
    .a(_al_u5353_o),
    .b(_al_u5583_o),
    .c(wb_ins_pc[14]),
    .o(\cu_ru/m_s_epc/n2 [14]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5585 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [14]),
    .c(data_csr[14]),
    .o(_al_u5585_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5586 (
    .a(\cu_ru/m_s_epc/n2 [14]),
    .b(_al_u5157_o),
    .c(_al_u5585_o),
    .o(\cu_ru/m_s_epc/n8 [14]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5587 (
    .a(\cu_ru/m_s_epc/n0 [11]),
    .b(pc_jmp),
    .c(new_pc[13]),
    .o(_al_u5587_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5588 (
    .a(_al_u5353_o),
    .b(_al_u5587_o),
    .c(wb_ins_pc[13]),
    .o(\cu_ru/m_s_epc/n2 [13]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5589 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [13]),
    .c(data_csr[13]),
    .o(_al_u5589_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5590 (
    .a(\cu_ru/m_s_epc/n2 [13]),
    .b(_al_u5157_o),
    .c(_al_u5589_o),
    .o(\cu_ru/m_s_epc/n8 [13]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5591 (
    .a(\cu_ru/m_s_epc/n0 [10]),
    .b(pc_jmp),
    .c(new_pc[12]),
    .o(_al_u5591_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5592 (
    .a(_al_u5353_o),
    .b(_al_u5591_o),
    .c(wb_ins_pc[12]),
    .o(\cu_ru/m_s_epc/n2 [12]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5593 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [12]),
    .c(data_csr[12]),
    .o(_al_u5593_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5594 (
    .a(\cu_ru/m_s_epc/n2 [12]),
    .b(_al_u5157_o),
    .c(_al_u5593_o),
    .o(\cu_ru/m_s_epc/n8 [12]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5595 (
    .a(\cu_ru/m_s_epc/n0 [9]),
    .b(pc_jmp),
    .c(new_pc[11]),
    .o(_al_u5595_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5596 (
    .a(_al_u5353_o),
    .b(_al_u5595_o),
    .c(wb_ins_pc[11]),
    .o(\cu_ru/m_s_epc/n2 [11]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5597 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [11]),
    .c(data_csr[11]),
    .o(_al_u5597_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5598 (
    .a(\cu_ru/m_s_epc/n2 [11]),
    .b(_al_u5157_o),
    .c(_al_u5597_o),
    .o(\cu_ru/m_s_epc/n8 [11]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5599 (
    .a(\cu_ru/m_s_epc/n0 [8]),
    .b(pc_jmp),
    .c(new_pc[10]),
    .o(_al_u5599_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'hb1))
    _al_u5600 (
    .a(_al_u5353_o),
    .b(_al_u5599_o),
    .c(wb_ins_pc[10]),
    .o(\cu_ru/m_s_epc/n2 [10]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5601 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [10]),
    .c(data_csr[10]),
    .o(_al_u5601_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5602 (
    .a(\cu_ru/m_s_epc/n2 [10]),
    .b(_al_u5157_o),
    .c(_al_u5601_o),
    .o(\cu_ru/m_s_epc/n8 [10]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((B*~A))+D*C*~((B*~A))+~(D)*C*(B*~A)+D*C*(B*~A))"),
    .INIT(16'hfb40))
    _al_u5603 (
    .a(_al_u5353_o),
    .b(pc_jmp),
    .c(new_pc[1]),
    .d(wb_ins_pc[1]),
    .o(\cu_ru/m_s_epc/n2 [1]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5604 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [1]),
    .c(data_csr[1]),
    .o(_al_u5604_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5605 (
    .a(\cu_ru/m_s_epc/n2 [1]),
    .b(_al_u5157_o),
    .c(_al_u5604_o),
    .o(\cu_ru/m_s_epc/n8 [1]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((B*~A))+D*C*~((B*~A))+~(D)*C*(B*~A)+D*C*(B*~A))"),
    .INIT(16'hfb40))
    _al_u5606 (
    .a(_al_u5353_o),
    .b(pc_jmp),
    .c(new_pc[0]),
    .d(wb_ins_pc[0]),
    .o(\cu_ru/m_s_epc/n2 [0]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5607 (
    .a(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/sepc [0]),
    .c(data_csr[0]),
    .o(_al_u5607_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5608 (
    .a(\cu_ru/m_s_epc/n2 [0]),
    .b(_al_u5157_o),
    .c(_al_u5607_o),
    .o(\cu_ru/m_s_epc/n8 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5609 (
    .a(_al_u5158_o),
    .b(_al_u3206_o),
    .o(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5610 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [9]),
    .d(data_csr[9]),
    .o(\cu_ru/m_s_cause/n5 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5611 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [8]),
    .d(data_csr[8]),
    .o(\cu_ru/m_s_cause/n5 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5612 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [7]),
    .d(data_csr[7]),
    .o(\cu_ru/m_s_cause/n5 [7]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5613 (
    .a(_al_u5157_o),
    .b(_al_u4234_o),
    .o(\cu_ru/n41 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5614 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [63]),
    .d(data_csr[63]),
    .o(_al_u5614_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5615 (
    .a(\cu_ru/n41 ),
    .b(_al_u5614_o),
    .o(\cu_ru/m_s_cause/n5 [63]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5616 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [62]),
    .d(data_csr[62]),
    .o(\cu_ru/m_s_cause/n5 [62]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5617 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [61]),
    .d(data_csr[61]),
    .o(\cu_ru/m_s_cause/n5 [61]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5618 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [60]),
    .d(data_csr[60]),
    .o(\cu_ru/m_s_cause/n5 [60]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5619 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [6]),
    .d(data_csr[6]),
    .o(\cu_ru/m_s_cause/n5 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5620 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [59]),
    .d(data_csr[59]),
    .o(\cu_ru/m_s_cause/n5 [59]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5621 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [58]),
    .d(data_csr[58]),
    .o(\cu_ru/m_s_cause/n5 [58]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5622 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [57]),
    .d(data_csr[57]),
    .o(\cu_ru/m_s_cause/n5 [57]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5623 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [56]),
    .d(data_csr[56]),
    .o(\cu_ru/m_s_cause/n5 [56]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5624 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [55]),
    .d(data_csr[55]),
    .o(\cu_ru/m_s_cause/n5 [55]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5625 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [54]),
    .d(data_csr[54]),
    .o(\cu_ru/m_s_cause/n5 [54]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5626 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [53]),
    .d(data_csr[53]),
    .o(\cu_ru/m_s_cause/n5 [53]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5627 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [52]),
    .d(data_csr[52]),
    .o(\cu_ru/m_s_cause/n5 [52]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5628 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [51]),
    .d(data_csr[51]),
    .o(\cu_ru/m_s_cause/n5 [51]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5629 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [50]),
    .d(data_csr[50]),
    .o(\cu_ru/m_s_cause/n5 [50]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5630 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [5]),
    .d(data_csr[5]),
    .o(\cu_ru/m_s_cause/n5 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5631 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [49]),
    .d(data_csr[49]),
    .o(\cu_ru/m_s_cause/n5 [49]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5632 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [48]),
    .d(data_csr[48]),
    .o(\cu_ru/m_s_cause/n5 [48]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5633 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [47]),
    .d(data_csr[47]),
    .o(\cu_ru/m_s_cause/n5 [47]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5634 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [46]),
    .d(data_csr[46]),
    .o(\cu_ru/m_s_cause/n5 [46]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5635 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [45]),
    .d(data_csr[45]),
    .o(\cu_ru/m_s_cause/n5 [45]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5636 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [44]),
    .d(data_csr[44]),
    .o(\cu_ru/m_s_cause/n5 [44]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5637 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [43]),
    .d(data_csr[43]),
    .o(\cu_ru/m_s_cause/n5 [43]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5638 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [42]),
    .d(data_csr[42]),
    .o(\cu_ru/m_s_cause/n5 [42]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5639 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [41]),
    .d(data_csr[41]),
    .o(\cu_ru/m_s_cause/n5 [41]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5640 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [40]),
    .d(data_csr[40]),
    .o(\cu_ru/m_s_cause/n5 [40]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5641 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [4]),
    .d(data_csr[4]),
    .o(\cu_ru/m_s_cause/n5 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5642 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [39]),
    .d(data_csr[39]),
    .o(\cu_ru/m_s_cause/n5 [39]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5643 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [38]),
    .d(data_csr[38]),
    .o(\cu_ru/m_s_cause/n5 [38]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5644 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [37]),
    .d(data_csr[37]),
    .o(\cu_ru/m_s_cause/n5 [37]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5645 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [36]),
    .d(data_csr[36]),
    .o(\cu_ru/m_s_cause/n5 [36]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5646 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [35]),
    .d(data_csr[35]),
    .o(\cu_ru/m_s_cause/n5 [35]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5647 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [34]),
    .d(data_csr[34]),
    .o(\cu_ru/m_s_cause/n5 [34]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5648 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [33]),
    .d(data_csr[33]),
    .o(\cu_ru/m_s_cause/n5 [33]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5649 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [32]),
    .d(data_csr[32]),
    .o(\cu_ru/m_s_cause/n5 [32]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5650 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [31]),
    .d(data_csr[31]),
    .o(\cu_ru/m_s_cause/n5 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5651 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [30]),
    .d(data_csr[30]),
    .o(\cu_ru/m_s_cause/n5 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5652 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [29]),
    .d(data_csr[29]),
    .o(\cu_ru/m_s_cause/n5 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5653 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [28]),
    .d(data_csr[28]),
    .o(\cu_ru/m_s_cause/n5 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5654 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [27]),
    .d(data_csr[27]),
    .o(\cu_ru/m_s_cause/n5 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5655 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [26]),
    .d(data_csr[26]),
    .o(\cu_ru/m_s_cause/n5 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5656 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [25]),
    .d(data_csr[25]),
    .o(\cu_ru/m_s_cause/n5 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5657 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [24]),
    .d(data_csr[24]),
    .o(\cu_ru/m_s_cause/n5 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5658 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [23]),
    .d(data_csr[23]),
    .o(\cu_ru/m_s_cause/n5 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5659 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [22]),
    .d(data_csr[22]),
    .o(\cu_ru/m_s_cause/n5 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5660 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [21]),
    .d(data_csr[21]),
    .o(\cu_ru/m_s_cause/n5 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5661 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [20]),
    .d(data_csr[20]),
    .o(\cu_ru/m_s_cause/n5 [20]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u5662 (
    .a(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .b(\cu_ru/scause [2]),
    .c(data_csr[2]),
    .o(_al_u5662_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u5663 (
    .a(\cu_ru/trap_cause [2]),
    .b(_al_u5157_o),
    .c(_al_u5662_o),
    .o(\cu_ru/m_s_cause/n5 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5664 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [19]),
    .d(data_csr[19]),
    .o(\cu_ru/m_s_cause/n5 [19]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5665 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [18]),
    .d(data_csr[18]),
    .o(\cu_ru/m_s_cause/n5 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5666 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [17]),
    .d(data_csr[17]),
    .o(\cu_ru/m_s_cause/n5 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5667 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [16]),
    .d(data_csr[16]),
    .o(\cu_ru/m_s_cause/n5 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5668 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [15]),
    .d(data_csr[15]),
    .o(\cu_ru/m_s_cause/n5 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5669 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [14]),
    .d(data_csr[14]),
    .o(\cu_ru/m_s_cause/n5 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5670 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [13]),
    .d(data_csr[13]),
    .o(\cu_ru/m_s_cause/n5 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5671 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [12]),
    .d(data_csr[12]),
    .o(\cu_ru/m_s_cause/n5 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5672 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [11]),
    .d(data_csr[11]),
    .o(\cu_ru/m_s_cause/n5 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u5673 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [10]),
    .d(data_csr[10]),
    .o(\cu_ru/m_s_cause/n5 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u5674 (
    .a(_al_u5157_o),
    .b(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .c(\cu_ru/scause [0]),
    .d(data_csr[0]),
    .o(_al_u5674_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u5675 (
    .a(_al_u4232_o),
    .b(\cu_ru/n41 ),
    .c(_al_u5674_o),
    .o(\cu_ru/m_s_cause/n5 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5676 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [63]),
    .d(\biu/cache_ctrl_logic/l1d_pte [63]),
    .o(_al_u5676_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5677 (
    .a(_al_u2705_o),
    .b(_al_u5676_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [63]),
    .o(_al_u5677_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5678 (
    .a(_al_u4238_o),
    .b(_al_u5677_o),
    .c(_al_u3222_o),
    .o(_al_u5678_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5679 (
    .a(_al_u5678_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [63]),
    .o(hwdata_pad[63]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5680 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [62]),
    .d(\biu/cache_ctrl_logic/l1d_pte [62]),
    .o(_al_u5680_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5681 (
    .a(_al_u2705_o),
    .b(_al_u5680_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [62]),
    .o(_al_u5681_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5682 (
    .a(_al_u4242_o),
    .b(_al_u5681_o),
    .c(_al_u3222_o),
    .o(_al_u5682_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5683 (
    .a(_al_u5682_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [62]),
    .o(hwdata_pad[62]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5684 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [61]),
    .d(\biu/cache_ctrl_logic/pte_temp [61]),
    .o(_al_u5684_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5685 (
    .a(_al_u2705_o),
    .b(_al_u5684_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [61]),
    .o(_al_u5685_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5686 (
    .a(_al_u4246_o),
    .b(_al_u5685_o),
    .c(_al_u3222_o),
    .o(_al_u5686_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5687 (
    .a(_al_u5686_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [61]),
    .o(hwdata_pad[61]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5688 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [60]),
    .d(\biu/cache_ctrl_logic/l1d_pte [60]),
    .o(_al_u5688_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5689 (
    .a(_al_u2705_o),
    .b(_al_u5688_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [60]),
    .o(_al_u5689_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5690 (
    .a(_al_u4250_o),
    .b(_al_u5689_o),
    .c(_al_u3222_o),
    .o(_al_u5690_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5691 (
    .a(_al_u5690_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [60]),
    .o(hwdata_pad[60]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5692 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [59]),
    .d(\biu/cache_ctrl_logic/l1d_pte [59]),
    .o(_al_u5692_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5693 (
    .a(_al_u2705_o),
    .b(_al_u5692_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [59]),
    .o(_al_u5693_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5694 (
    .a(_al_u4254_o),
    .b(_al_u5693_o),
    .c(_al_u3222_o),
    .o(_al_u5694_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5695 (
    .a(_al_u5694_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [59]),
    .o(hwdata_pad[59]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5696 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [58]),
    .d(\biu/cache_ctrl_logic/l1d_pte [58]),
    .o(_al_u5696_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5697 (
    .a(_al_u2705_o),
    .b(_al_u5696_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [58]),
    .o(_al_u5697_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5698 (
    .a(_al_u4258_o),
    .b(_al_u5697_o),
    .c(_al_u3222_o),
    .o(_al_u5698_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5699 (
    .a(_al_u5698_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [58]),
    .o(hwdata_pad[58]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5700 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [57]),
    .d(\biu/cache_ctrl_logic/pte_temp [57]),
    .o(_al_u5700_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5701 (
    .a(_al_u2705_o),
    .b(_al_u5700_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [57]),
    .o(_al_u5701_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5702 (
    .a(_al_u4262_o),
    .b(_al_u5701_o),
    .c(_al_u3222_o),
    .o(_al_u5702_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5703 (
    .a(_al_u5702_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [57]),
    .o(hwdata_pad[57]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5704 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [56]),
    .d(\biu/cache_ctrl_logic/l1d_pte [56]),
    .o(_al_u5704_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5705 (
    .a(_al_u2705_o),
    .b(_al_u5704_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [56]),
    .o(_al_u5705_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5706 (
    .a(_al_u4266_o),
    .b(_al_u5705_o),
    .c(_al_u3222_o),
    .o(_al_u5706_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5707 (
    .a(_al_u5706_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [56]),
    .o(hwdata_pad[56]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5708 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [55]),
    .d(\biu/cache_ctrl_logic/pte_temp [55]),
    .o(_al_u5708_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5709 (
    .a(_al_u2705_o),
    .b(_al_u5708_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [55]),
    .o(_al_u5709_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5710 (
    .a(_al_u4270_o),
    .b(_al_u5709_o),
    .c(_al_u3222_o),
    .o(_al_u5710_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5711 (
    .a(_al_u5710_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [55]),
    .o(hwdata_pad[55]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5712 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [54]),
    .d(\biu/cache_ctrl_logic/pte_temp [54]),
    .o(_al_u5712_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5713 (
    .a(_al_u2705_o),
    .b(_al_u5712_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [54]),
    .o(_al_u5713_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5714 (
    .a(_al_u4274_o),
    .b(_al_u5713_o),
    .c(_al_u3222_o),
    .o(_al_u5714_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5715 (
    .a(_al_u5714_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [54]),
    .o(hwdata_pad[54]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5716 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [53]),
    .d(\biu/cache_ctrl_logic/pte_temp [53]),
    .o(_al_u5716_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5717 (
    .a(_al_u2705_o),
    .b(_al_u5716_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [53]),
    .o(_al_u5717_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5718 (
    .a(_al_u4278_o),
    .b(_al_u5717_o),
    .c(_al_u3222_o),
    .o(_al_u5718_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5719 (
    .a(_al_u5718_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [53]),
    .o(hwdata_pad[53]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5720 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [52]),
    .d(\biu/cache_ctrl_logic/l1d_pte [52]),
    .o(_al_u5720_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5721 (
    .a(_al_u2705_o),
    .b(_al_u5720_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [52]),
    .o(_al_u5721_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5722 (
    .a(_al_u4282_o),
    .b(_al_u5721_o),
    .c(_al_u3222_o),
    .o(_al_u5722_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5723 (
    .a(_al_u5722_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [52]),
    .o(hwdata_pad[52]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5724 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [51]),
    .d(\biu/cache_ctrl_logic/pte_temp [51]),
    .o(_al_u5724_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5725 (
    .a(_al_u2705_o),
    .b(_al_u5724_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [51]),
    .o(_al_u5725_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5726 (
    .a(_al_u4286_o),
    .b(_al_u5725_o),
    .c(_al_u3222_o),
    .o(_al_u5726_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5727 (
    .a(_al_u5726_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [51]),
    .o(hwdata_pad[51]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5728 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [50]),
    .d(\biu/cache_ctrl_logic/pte_temp [50]),
    .o(_al_u5728_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5729 (
    .a(_al_u2705_o),
    .b(_al_u5728_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [50]),
    .o(_al_u5729_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5730 (
    .a(_al_u4290_o),
    .b(_al_u5729_o),
    .c(_al_u3222_o),
    .o(_al_u5730_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5731 (
    .a(_al_u5730_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [50]),
    .o(hwdata_pad[50]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5732 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [49]),
    .d(\biu/cache_ctrl_logic/l1d_pte [49]),
    .o(_al_u5732_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5733 (
    .a(_al_u2705_o),
    .b(_al_u5732_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [49]),
    .o(_al_u5733_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5734 (
    .a(_al_u4294_o),
    .b(_al_u5733_o),
    .c(_al_u3222_o),
    .o(_al_u5734_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5735 (
    .a(_al_u5734_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [49]),
    .o(hwdata_pad[49]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5736 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [48]),
    .d(\biu/cache_ctrl_logic/l1d_pte [48]),
    .o(_al_u5736_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5737 (
    .a(_al_u2705_o),
    .b(_al_u5736_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [48]),
    .o(_al_u5737_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5738 (
    .a(_al_u4298_o),
    .b(_al_u5737_o),
    .c(_al_u3222_o),
    .o(_al_u5738_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5739 (
    .a(_al_u5738_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [48]),
    .o(hwdata_pad[48]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5740 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [47]),
    .d(\biu/cache_ctrl_logic/pte_temp [47]),
    .o(_al_u5740_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5741 (
    .a(_al_u2705_o),
    .b(_al_u5740_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [47]),
    .o(_al_u5741_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5742 (
    .a(_al_u4302_o),
    .b(_al_u5741_o),
    .c(_al_u3222_o),
    .o(_al_u5742_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5743 (
    .a(_al_u5742_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [47]),
    .o(hwdata_pad[47]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5744 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [46]),
    .d(\biu/cache_ctrl_logic/l1d_pte [46]),
    .o(_al_u5744_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5745 (
    .a(_al_u2705_o),
    .b(_al_u5744_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [46]),
    .o(_al_u5745_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5746 (
    .a(_al_u4306_o),
    .b(_al_u5745_o),
    .c(_al_u3222_o),
    .o(_al_u5746_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5747 (
    .a(_al_u5746_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [46]),
    .o(hwdata_pad[46]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5748 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [45]),
    .d(\biu/cache_ctrl_logic/pte_temp [45]),
    .o(_al_u5748_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5749 (
    .a(_al_u2705_o),
    .b(_al_u5748_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [45]),
    .o(_al_u5749_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5750 (
    .a(_al_u4310_o),
    .b(_al_u5749_o),
    .c(_al_u3222_o),
    .o(_al_u5750_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5751 (
    .a(_al_u5750_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [45]),
    .o(hwdata_pad[45]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5752 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [44]),
    .d(\biu/cache_ctrl_logic/pte_temp [44]),
    .o(_al_u5752_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5753 (
    .a(_al_u2705_o),
    .b(_al_u5752_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [44]),
    .o(_al_u5753_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5754 (
    .a(_al_u4314_o),
    .b(_al_u5753_o),
    .c(_al_u3222_o),
    .o(_al_u5754_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5755 (
    .a(_al_u5754_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [44]),
    .o(hwdata_pad[44]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5756 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [43]),
    .d(\biu/cache_ctrl_logic/l1d_pte [43]),
    .o(_al_u5756_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5757 (
    .a(_al_u2705_o),
    .b(_al_u5756_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [43]),
    .o(_al_u5757_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5758 (
    .a(_al_u4318_o),
    .b(_al_u5757_o),
    .c(_al_u3222_o),
    .o(_al_u5758_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5759 (
    .a(_al_u5758_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [43]),
    .o(hwdata_pad[43]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5760 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [42]),
    .d(\biu/cache_ctrl_logic/l1d_pte [42]),
    .o(_al_u5760_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5761 (
    .a(_al_u2705_o),
    .b(_al_u5760_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [42]),
    .o(_al_u5761_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5762 (
    .a(_al_u4322_o),
    .b(_al_u5761_o),
    .c(_al_u3222_o),
    .o(_al_u5762_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5763 (
    .a(_al_u5762_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [42]),
    .o(hwdata_pad[42]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5764 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [41]),
    .d(\biu/cache_ctrl_logic/l1d_pte [41]),
    .o(_al_u5764_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5765 (
    .a(_al_u2705_o),
    .b(_al_u5764_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [41]),
    .o(_al_u5765_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5766 (
    .a(_al_u4326_o),
    .b(_al_u5765_o),
    .c(_al_u3222_o),
    .o(_al_u5766_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5767 (
    .a(_al_u5766_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [41]),
    .o(hwdata_pad[41]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5768 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [40]),
    .d(\biu/cache_ctrl_logic/pte_temp [40]),
    .o(_al_u5768_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5769 (
    .a(_al_u2705_o),
    .b(_al_u5768_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [40]),
    .o(_al_u5769_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5770 (
    .a(_al_u4330_o),
    .b(_al_u5769_o),
    .c(_al_u3222_o),
    .o(_al_u5770_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5771 (
    .a(_al_u5770_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [40]),
    .o(hwdata_pad[40]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5772 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [39]),
    .d(\biu/cache_ctrl_logic/l1d_pte [39]),
    .o(_al_u5772_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5773 (
    .a(_al_u2705_o),
    .b(_al_u5772_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [39]),
    .o(_al_u5773_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5774 (
    .a(_al_u4334_o),
    .b(_al_u5773_o),
    .c(_al_u3222_o),
    .o(_al_u5774_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5775 (
    .a(_al_u5774_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [39]),
    .o(hwdata_pad[39]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5776 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [38]),
    .d(\biu/cache_ctrl_logic/l1d_pte [38]),
    .o(_al_u5776_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5777 (
    .a(_al_u2705_o),
    .b(_al_u5776_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [38]),
    .o(_al_u5777_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5778 (
    .a(_al_u4338_o),
    .b(_al_u5777_o),
    .c(_al_u3222_o),
    .o(_al_u5778_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5779 (
    .a(_al_u5778_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [38]),
    .o(hwdata_pad[38]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5780 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [37]),
    .d(\biu/cache_ctrl_logic/l1d_pte [37]),
    .o(_al_u5780_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5781 (
    .a(_al_u2705_o),
    .b(_al_u5780_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [37]),
    .o(_al_u5781_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5782 (
    .a(_al_u4342_o),
    .b(_al_u5781_o),
    .c(_al_u3222_o),
    .o(_al_u5782_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5783 (
    .a(_al_u5782_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [37]),
    .o(hwdata_pad[37]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5784 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [36]),
    .d(\biu/cache_ctrl_logic/pte_temp [36]),
    .o(_al_u5784_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5785 (
    .a(_al_u2705_o),
    .b(_al_u5784_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [36]),
    .o(_al_u5785_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5786 (
    .a(_al_u4346_o),
    .b(_al_u5785_o),
    .c(_al_u3222_o),
    .o(_al_u5786_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5787 (
    .a(_al_u5786_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [36]),
    .o(hwdata_pad[36]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5788 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [35]),
    .d(\biu/cache_ctrl_logic/pte_temp [35]),
    .o(_al_u5788_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5789 (
    .a(_al_u2705_o),
    .b(_al_u5788_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [35]),
    .o(_al_u5789_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5790 (
    .a(_al_u4350_o),
    .b(_al_u5789_o),
    .c(_al_u3222_o),
    .o(_al_u5790_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5791 (
    .a(_al_u5790_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [35]),
    .o(hwdata_pad[35]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5792 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [34]),
    .d(\biu/cache_ctrl_logic/l1d_pte [34]),
    .o(_al_u5792_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5793 (
    .a(_al_u2705_o),
    .b(_al_u5792_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [34]),
    .o(_al_u5793_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5794 (
    .a(_al_u4354_o),
    .b(_al_u5793_o),
    .c(_al_u3222_o),
    .o(_al_u5794_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5795 (
    .a(_al_u5794_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [34]),
    .o(hwdata_pad[34]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5796 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [33]),
    .d(\biu/cache_ctrl_logic/l1d_pte [33]),
    .o(_al_u5796_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5797 (
    .a(_al_u2705_o),
    .b(_al_u5796_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [33]),
    .o(_al_u5797_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5798 (
    .a(_al_u4358_o),
    .b(_al_u5797_o),
    .c(_al_u3222_o),
    .o(_al_u5798_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5799 (
    .a(_al_u5798_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [33]),
    .o(hwdata_pad[33]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5800 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [32]),
    .d(\biu/cache_ctrl_logic/pte_temp [32]),
    .o(_al_u5800_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5801 (
    .a(_al_u2705_o),
    .b(_al_u5800_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [32]),
    .o(_al_u5801_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5802 (
    .a(_al_u4362_o),
    .b(_al_u5801_o),
    .c(_al_u3222_o),
    .o(_al_u5802_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5803 (
    .a(_al_u5802_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [32]),
    .o(hwdata_pad[32]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5804 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [31]),
    .d(\biu/cache_ctrl_logic/pte_temp [31]),
    .o(_al_u5804_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5805 (
    .a(_al_u2705_o),
    .b(_al_u5804_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [31]),
    .o(_al_u5805_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5806 (
    .a(_al_u4366_o),
    .b(_al_u5805_o),
    .c(_al_u3222_o),
    .o(_al_u5806_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5807 (
    .a(_al_u5806_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [31]),
    .o(hwdata_pad[31]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5808 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [30]),
    .d(\biu/cache_ctrl_logic/l1d_pte [30]),
    .o(_al_u5808_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5809 (
    .a(_al_u2705_o),
    .b(_al_u5808_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [30]),
    .o(_al_u5809_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5810 (
    .a(_al_u4370_o),
    .b(_al_u5809_o),
    .c(_al_u3222_o),
    .o(_al_u5810_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5811 (
    .a(_al_u5810_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [30]),
    .o(hwdata_pad[30]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5812 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [29]),
    .d(\biu/cache_ctrl_logic/l1d_pte [29]),
    .o(_al_u5812_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5813 (
    .a(_al_u2705_o),
    .b(_al_u5812_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [29]),
    .o(_al_u5813_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5814 (
    .a(_al_u4374_o),
    .b(_al_u5813_o),
    .c(_al_u3222_o),
    .o(_al_u5814_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5815 (
    .a(_al_u5814_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [29]),
    .o(hwdata_pad[29]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5816 (
    .a(_al_u3945_o),
    .b(_al_u3947_o),
    .c(\biu/cache_ctrl_logic/l1d_pte [28]),
    .d(\biu/cache_ctrl_logic/pte_temp [28]),
    .o(_al_u5816_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5817 (
    .a(_al_u2705_o),
    .b(_al_u5816_o),
    .c(_al_u3950_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [28]),
    .o(_al_u5817_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5818 (
    .a(_al_u4378_o),
    .b(_al_u5817_o),
    .c(_al_u3222_o),
    .o(_al_u5818_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5819 (
    .a(_al_u5818_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [28]),
    .o(hwdata_pad[28]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5820 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [27]),
    .d(\biu/cache_ctrl_logic/l1d_pte [27]),
    .o(_al_u5820_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5821 (
    .a(_al_u2705_o),
    .b(_al_u5820_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [27]),
    .o(_al_u5821_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5822 (
    .a(_al_u4382_o),
    .b(_al_u5821_o),
    .c(_al_u3222_o),
    .o(_al_u5822_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5823 (
    .a(_al_u5822_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [27]),
    .o(hwdata_pad[27]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5824 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [26]),
    .d(\biu/cache_ctrl_logic/pte_temp [26]),
    .o(_al_u5824_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5825 (
    .a(_al_u2705_o),
    .b(_al_u5824_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [26]),
    .o(_al_u5825_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5826 (
    .a(_al_u4386_o),
    .b(_al_u5825_o),
    .c(_al_u3222_o),
    .o(_al_u5826_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5827 (
    .a(_al_u5826_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [26]),
    .o(hwdata_pad[26]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5828 (
    .a(_al_u3945_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [25]),
    .d(\biu/cache_ctrl_logic/pte_temp [25]),
    .o(_al_u5828_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5829 (
    .a(_al_u2705_o),
    .b(_al_u5828_o),
    .c(_al_u3947_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [25]),
    .o(_al_u5829_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5830 (
    .a(_al_u4390_o),
    .b(_al_u5829_o),
    .c(_al_u3222_o),
    .o(_al_u5830_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5831 (
    .a(_al_u5830_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [25]),
    .o(hwdata_pad[25]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u5832 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [24]),
    .d(\biu/cache_ctrl_logic/l1d_pte [24]),
    .o(_al_u5832_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u5833 (
    .a(_al_u2705_o),
    .b(_al_u5832_o),
    .c(_al_u3945_o),
    .d(\biu/cache_ctrl_logic/pte_temp [24]),
    .o(_al_u5833_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u5834 (
    .a(_al_u4394_o),
    .b(_al_u5833_o),
    .c(_al_u3222_o),
    .o(_al_u5834_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u5835 (
    .a(_al_u5834_o),
    .b(_al_u2705_o),
    .c(\biu/bus_unit/mmu_hwdata [24]),
    .o(hwdata_pad[24]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u5836 (
    .a(_al_u4092_o),
    .b(\ins_dec/ins_srai ),
    .c(_al_u3217_o),
    .d(_al_u3384_o),
    .o(\ins_dec/n57_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5837 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_005 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_005 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5837_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u5838 (
    .a(\ins_dec/n57_neg_lutinv ),
    .b(_al_u5837_o),
    .c(id_ins[20]),
    .o(\ins_dec/op_count_decode [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5839 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_004 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_004 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5839_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u5840 (
    .a(\ins_dec/n57_neg_lutinv ),
    .b(_al_u5839_o),
    .c(id_ins[19]),
    .o(\ins_dec/op_count_decode [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5841 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_003 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_003 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5841_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u5842 (
    .a(\ins_dec/n57_neg_lutinv ),
    .b(_al_u5841_o),
    .c(id_ins[18]),
    .o(\ins_dec/op_count_decode [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5843 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_002 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_002 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5843_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u5844 (
    .a(\ins_dec/n57_neg_lutinv ),
    .b(_al_u5843_o),
    .c(id_ins[17]),
    .o(\ins_dec/op_count_decode [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5845 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_001 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_001 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5845_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u5846 (
    .a(\ins_dec/n57_neg_lutinv ),
    .b(_al_u5845_o),
    .c(id_ins[16]),
    .o(\ins_dec/op_count_decode [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5847 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_000 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_000 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5847_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u5848 (
    .a(\ins_dec/n57_neg_lutinv ),
    .b(_al_u5847_o),
    .c(id_ins[15]),
    .o(\ins_dec/op_count_decode [0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u5849 (
    .a(\ins_dec/n239 ),
    .b(_al_u3216_o),
    .o(\ins_dec/mux19_b10_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .INIT(16'h07f7))
    _al_u5850 (
    .a(rs1_data[9]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3927_o),
    .d(id_ins[29]),
    .o(_al_u5850_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u5851 (
    .a(_al_u5143_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_009 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_009 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5851_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u5852 (
    .a(_al_u5850_o),
    .b(_al_u5851_o),
    .c(_al_u4086_o),
    .o(\ins_dec/n284 [9]));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .INIT(16'h07f7))
    _al_u5853 (
    .a(rs1_data[8]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3927_o),
    .d(id_ins[28]),
    .o(_al_u5853_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u5854 (
    .a(_al_u5143_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_008 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_008 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5854_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u5855 (
    .a(_al_u5853_o),
    .b(_al_u5854_o),
    .c(_al_u4086_o),
    .o(\ins_dec/n284 [8]));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .INIT(16'h07f7))
    _al_u5856 (
    .a(rs1_data[7]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3927_o),
    .d(id_ins[27]),
    .o(_al_u5856_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5857 (
    .a(_al_u5856_o),
    .b(\ins_dec/op_count_decode [7]),
    .o(\ins_dec/n284 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5858 (
    .a(_al_u3955_o),
    .b(id_ins[31]),
    .o(_al_u5858_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5859 (
    .a(rs1_data[63]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u5859_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5860 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_063 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_063 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5860_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5861 (
    .a(_al_u5859_o),
    .b(_al_u5860_o),
    .o(\ins_dec/n284 [63]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5862 (
    .a(rs1_data[62]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u5862_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5863 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_062 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_062 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5863_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5864 (
    .a(_al_u5862_o),
    .b(_al_u5863_o),
    .o(\ins_dec/n284 [62]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5865 (
    .a(rs1_data[61]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u5865_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5866 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_061 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_061 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5866_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5867 (
    .a(_al_u5865_o),
    .b(_al_u5866_o),
    .o(\ins_dec/n284 [61]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5868 (
    .a(rs1_data[60]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u5868_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5869 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_060 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_060 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5869_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5870 (
    .a(_al_u5868_o),
    .b(_al_u5869_o),
    .o(\ins_dec/n284 [60]));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .INIT(16'h07f7))
    _al_u5871 (
    .a(rs1_data[6]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3927_o),
    .d(id_ins[26]),
    .o(_al_u5871_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5872 (
    .a(_al_u5871_o),
    .b(\ins_dec/op_count_decode [6]),
    .o(\ins_dec/n284 [6]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5873 (
    .a(rs1_data[59]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u5873_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5874 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_059 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_059 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5874_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5875 (
    .a(_al_u5873_o),
    .b(_al_u5874_o),
    .o(\ins_dec/n284 [59]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5876 (
    .a(rs1_data[58]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u5876_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5877 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_058 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_058 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5877_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5878 (
    .a(_al_u5876_o),
    .b(_al_u5877_o),
    .o(\ins_dec/n284 [58]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5879 (
    .a(rs1_data[57]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u5879_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5880 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_057 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_057 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5880_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5881 (
    .a(_al_u5879_o),
    .b(_al_u5880_o),
    .o(\ins_dec/n284 [57]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u5882 (
    .a(rs1_data[56]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u5882_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u5883 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_056 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_056 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5883_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5884 (
    .a(_al_u5882_o),
    .b(_al_u5883_o),
    .o(\ins_dec/n284 [56]));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .INIT(16'h07f7))
    _al_u5885 (
    .a(rs1_data[5]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3927_o),
    .d(id_ins[25]),
    .o(_al_u5885_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u5886 (
    .a(_al_u5885_o),
    .b(_al_u5837_o),
    .o(\ins_dec/n284 [5]));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .INIT(16'h07f7))
    _al_u5887 (
    .a(rs1_data[11]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3927_o),
    .d(id_ins[31]),
    .o(_al_u5887_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u5888 (
    .a(_al_u5143_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_011 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_011 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5888_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u5889 (
    .a(_al_u5887_o),
    .b(_al_u5888_o),
    .c(_al_u4086_o),
    .o(\ins_dec/n284 [11]));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .INIT(16'h07f7))
    _al_u5890 (
    .a(rs1_data[10]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3927_o),
    .d(id_ins[30]),
    .o(_al_u5890_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h5044))
    _al_u5891 (
    .a(_al_u5143_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_010 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_010 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u5891_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u5892 (
    .a(_al_u5890_o),
    .b(_al_u5891_o),
    .c(_al_u4086_o),
    .o(\ins_dec/n284 [10]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    _al_u5893 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [29]),
    .d(\biu/bus_unit/mmu_hwdata [27]),
    .o(_al_u5893_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5894 (
    .a(\biu/maddress [29]),
    .b(_al_u5893_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5894_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    .INIT(16'h2023))
    _al_u5895 (
    .a(_al_u5894_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [29]),
    .o(_al_u5895_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5896 (
    .a(\biu/maddress [29]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [29]),
    .o(_al_u5896_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5897 (
    .a(_al_u5895_o),
    .b(_al_u5896_o),
    .o(\biu/bus_unit/mmu/n66 [29]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    _al_u5898 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [28]),
    .d(\biu/bus_unit/mmu_hwdata [26]),
    .o(_al_u5898_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5899 (
    .a(\biu/maddress [28]),
    .b(_al_u5898_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5899_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    .INIT(16'h2023))
    _al_u5900 (
    .a(_al_u5899_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [28]),
    .o(_al_u5900_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5901 (
    .a(\biu/maddress [28]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [28]),
    .o(_al_u5901_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5902 (
    .a(_al_u5900_o),
    .b(_al_u5901_o),
    .o(\biu/bus_unit/mmu/n66 [28]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    _al_u5903 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [27]),
    .d(\biu/bus_unit/mmu_hwdata [25]),
    .o(_al_u5903_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5904 (
    .a(\biu/maddress [27]),
    .b(_al_u5903_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5904_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    .INIT(16'h2023))
    _al_u5905 (
    .a(_al_u5904_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [27]),
    .o(_al_u5905_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5906 (
    .a(\biu/maddress [27]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [27]),
    .o(_al_u5906_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5907 (
    .a(_al_u5905_o),
    .b(_al_u5906_o),
    .o(\biu/bus_unit/mmu/n66 [27]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    _al_u5908 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [26]),
    .d(\biu/bus_unit/mmu_hwdata [24]),
    .o(_al_u5908_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5909 (
    .a(\biu/maddress [26]),
    .b(_al_u5908_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5909_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    .INIT(16'h2023))
    _al_u5910 (
    .a(_al_u5909_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [26]),
    .o(_al_u5910_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5911 (
    .a(\biu/maddress [26]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [26]),
    .o(_al_u5911_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5912 (
    .a(_al_u5910_o),
    .b(_al_u5911_o),
    .o(\biu/bus_unit/mmu/n66 [26]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    _al_u5913 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [25]),
    .d(\biu/bus_unit/mmu_hwdata [23]),
    .o(_al_u5913_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5914 (
    .a(\biu/maddress [25]),
    .b(_al_u5913_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5914_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    .INIT(16'h2023))
    _al_u5915 (
    .a(_al_u5914_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [25]),
    .o(_al_u5915_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5916 (
    .a(\biu/maddress [25]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [25]),
    .o(_al_u5916_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5917 (
    .a(_al_u5915_o),
    .b(_al_u5916_o),
    .o(\biu/bus_unit/mmu/n66 [25]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    _al_u5918 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [24]),
    .d(\biu/bus_unit/mmu_hwdata [22]),
    .o(_al_u5918_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5919 (
    .a(\biu/maddress [24]),
    .b(_al_u5918_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5919_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    .INIT(16'h2023))
    _al_u5920 (
    .a(_al_u5919_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [24]),
    .o(_al_u5920_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5921 (
    .a(\biu/maddress [24]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [24]),
    .o(_al_u5921_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5922 (
    .a(_al_u5920_o),
    .b(_al_u5921_o),
    .o(\biu/bus_unit/mmu/n66 [24]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    _al_u5923 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [23]),
    .d(\biu/bus_unit/mmu_hwdata [21]),
    .o(_al_u5923_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5924 (
    .a(\biu/maddress [23]),
    .b(_al_u5923_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5924_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    .INIT(16'h2023))
    _al_u5925 (
    .a(_al_u5924_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [23]),
    .o(_al_u5925_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5926 (
    .a(\biu/maddress [23]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [23]),
    .o(_al_u5926_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5927 (
    .a(_al_u5925_o),
    .b(_al_u5926_o),
    .o(\biu/bus_unit/mmu/n66 [23]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    _al_u5928 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [22]),
    .d(\biu/bus_unit/mmu_hwdata [20]),
    .o(_al_u5928_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5929 (
    .a(\biu/maddress [22]),
    .b(_al_u5928_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5929_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    .INIT(16'h2023))
    _al_u5930 (
    .a(_al_u5929_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [22]),
    .o(_al_u5930_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5931 (
    .a(\biu/maddress [22]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [22]),
    .o(_al_u5931_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5932 (
    .a(_al_u5930_o),
    .b(_al_u5931_o),
    .o(\biu/bus_unit/mmu/n66 [22]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((C*A))*~(B)+D*(C*A)*~(B)+~(D)*(C*A)*B+D*(C*A)*B)"),
    .INIT(16'h4c7f))
    _al_u5933 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [21]),
    .d(\biu/bus_unit/mmu_hwdata [19]),
    .o(_al_u5933_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u5934 (
    .a(\biu/maddress [21]),
    .b(_al_u5933_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5934_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    .INIT(16'h2023))
    _al_u5935 (
    .a(_al_u5934_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [21]),
    .o(_al_u5935_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5936 (
    .a(\biu/maddress [21]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [21]),
    .o(_al_u5936_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5937 (
    .a(_al_u5935_o),
    .b(_al_u5936_o),
    .o(\biu/bus_unit/mmu/n66 [21]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5938 (
    .a(\biu/maddress [20]),
    .b(_al_u2914_o),
    .c(\biu/paddress [20]),
    .o(_al_u5938_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h6e7f))
    _al_u5939 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [20]),
    .d(\biu/bus_unit/mmu_hwdata [18]),
    .o(_al_u5939_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5940 (
    .a(_al_u2915_o),
    .b(_al_u5939_o),
    .o(_al_u5940_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*(D@C)))"),
    .INIT(16'hc44c))
    _al_u5941 (
    .a(\biu/maddress [20]),
    .b(_al_u5940_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5941_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5942 (
    .a(_al_u2915_o),
    .b(\biu/paddress [20]),
    .o(_al_u5942_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    .INIT(16'h5053))
    _al_u5943 (
    .a(_al_u5938_o),
    .b(_al_u5941_o),
    .c(_al_u2698_o),
    .d(_al_u5942_o),
    .o(\biu/bus_unit/mmu/n66 [20]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5944 (
    .a(\biu/maddress [19]),
    .b(_al_u2914_o),
    .c(\biu/paddress [19]),
    .o(_al_u5944_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h6e7f))
    _al_u5945 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [19]),
    .d(\biu/bus_unit/mmu_hwdata [17]),
    .o(_al_u5945_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5946 (
    .a(_al_u2915_o),
    .b(_al_u5945_o),
    .o(_al_u5946_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*(D@C)))"),
    .INIT(16'hc44c))
    _al_u5947 (
    .a(\biu/maddress [19]),
    .b(_al_u5946_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5947_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5948 (
    .a(_al_u2915_o),
    .b(\biu/paddress [19]),
    .o(_al_u5948_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    .INIT(16'h5053))
    _al_u5949 (
    .a(_al_u5944_o),
    .b(_al_u5947_o),
    .c(_al_u2698_o),
    .d(_al_u5948_o),
    .o(\biu/bus_unit/mmu/n66 [19]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5950 (
    .a(\biu/maddress [18]),
    .b(_al_u2914_o),
    .c(\biu/paddress [18]),
    .o(_al_u5950_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h6e7f))
    _al_u5951 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [18]),
    .d(\biu/bus_unit/mmu_hwdata [16]),
    .o(_al_u5951_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5952 (
    .a(_al_u2915_o),
    .b(_al_u5951_o),
    .o(_al_u5952_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*(D@C)))"),
    .INIT(16'hc44c))
    _al_u5953 (
    .a(\biu/maddress [18]),
    .b(_al_u5952_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5953_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5954 (
    .a(_al_u2915_o),
    .b(\biu/paddress [18]),
    .o(_al_u5954_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    .INIT(16'h5053))
    _al_u5955 (
    .a(_al_u5950_o),
    .b(_al_u5953_o),
    .c(_al_u2698_o),
    .d(_al_u5954_o),
    .o(\biu/bus_unit/mmu/n66 [18]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5956 (
    .a(\biu/maddress [17]),
    .b(_al_u2914_o),
    .c(\biu/paddress [17]),
    .o(_al_u5956_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h6e7f))
    _al_u5957 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [17]),
    .d(\biu/bus_unit/mmu_hwdata [15]),
    .o(_al_u5957_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5958 (
    .a(_al_u2915_o),
    .b(_al_u5957_o),
    .o(_al_u5958_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*(D@C)))"),
    .INIT(16'hc44c))
    _al_u5959 (
    .a(\biu/maddress [17]),
    .b(_al_u5958_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5959_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5960 (
    .a(_al_u2915_o),
    .b(\biu/paddress [17]),
    .o(_al_u5960_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    .INIT(16'h5053))
    _al_u5961 (
    .a(_al_u5956_o),
    .b(_al_u5959_o),
    .c(_al_u2698_o),
    .d(_al_u5960_o),
    .o(\biu/bus_unit/mmu/n66 [17]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5962 (
    .a(\biu/maddress [16]),
    .b(_al_u2914_o),
    .c(\biu/paddress [16]),
    .o(_al_u5962_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h6e7f))
    _al_u5963 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [16]),
    .d(\biu/bus_unit/mmu_hwdata [14]),
    .o(_al_u5963_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5964 (
    .a(_al_u2915_o),
    .b(_al_u5963_o),
    .o(_al_u5964_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*(D@C)))"),
    .INIT(16'hc44c))
    _al_u5965 (
    .a(\biu/maddress [16]),
    .b(_al_u5964_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5965_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5966 (
    .a(_al_u2915_o),
    .b(\biu/paddress [16]),
    .o(_al_u5966_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    .INIT(16'h5053))
    _al_u5967 (
    .a(_al_u5962_o),
    .b(_al_u5965_o),
    .c(_al_u2698_o),
    .d(_al_u5966_o),
    .o(\biu/bus_unit/mmu/n66 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h6e7f))
    _al_u5968 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [15]),
    .d(\biu/bus_unit/mmu_hwdata [13]),
    .o(_al_u5968_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5969 (
    .a(_al_u2915_o),
    .b(_al_u5968_o),
    .o(_al_u5969_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*(D@C)))"),
    .INIT(16'hc44c))
    _al_u5970 (
    .a(\biu/maddress [15]),
    .b(_al_u5969_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5970_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~A*~(~D*~C)))"),
    .INIT(16'h2223))
    _al_u5971 (
    .a(_al_u5970_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [15]),
    .o(_al_u5971_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5972 (
    .a(\biu/maddress [15]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [15]),
    .o(_al_u5972_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5973 (
    .a(_al_u5971_o),
    .b(_al_u5972_o),
    .o(\biu/bus_unit/mmu/n66 [15]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5974 (
    .a(\biu/maddress [14]),
    .b(_al_u2914_o),
    .c(\biu/paddress [14]),
    .o(_al_u5974_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h6e7f))
    _al_u5975 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [14]),
    .d(\biu/bus_unit/mmu_hwdata [12]),
    .o(_al_u5975_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5976 (
    .a(_al_u2915_o),
    .b(_al_u5975_o),
    .o(_al_u5976_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*(D@C)))"),
    .INIT(16'hc44c))
    _al_u5977 (
    .a(\biu/maddress [14]),
    .b(_al_u5976_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5977_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5978 (
    .a(_al_u2915_o),
    .b(\biu/paddress [14]),
    .o(_al_u5978_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    .INIT(16'h5053))
    _al_u5979 (
    .a(_al_u5974_o),
    .b(_al_u5977_o),
    .c(_al_u2698_o),
    .d(_al_u5978_o),
    .o(\biu/bus_unit/mmu/n66 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h6e7f))
    _al_u5980 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [13]),
    .d(\biu/bus_unit/mmu_hwdata [11]),
    .o(_al_u5980_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5981 (
    .a(_al_u2915_o),
    .b(_al_u5980_o),
    .o(_al_u5981_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*(D@C)))"),
    .INIT(16'hc44c))
    _al_u5982 (
    .a(\biu/maddress [13]),
    .b(_al_u5981_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5982_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~A*~(~D*~C)))"),
    .INIT(16'h2223))
    _al_u5983 (
    .a(_al_u5982_o),
    .b(_al_u2698_o),
    .c(_al_u2915_o),
    .d(\biu/paddress [13]),
    .o(_al_u5983_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    _al_u5984 (
    .a(\biu/maddress [13]),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(\biu/paddress [13]),
    .o(_al_u5984_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5985 (
    .a(_al_u5983_o),
    .b(_al_u5984_o),
    .o(\biu/bus_unit/mmu/n66 [13]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u5986 (
    .a(\biu/maddress [12]),
    .b(_al_u2914_o),
    .c(\biu/paddress [12]),
    .o(_al_u5986_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h6e7f))
    _al_u5987 (
    .a(\biu/bus_unit/mmu/i [0]),
    .b(\biu/bus_unit/mmu/i [1]),
    .c(\biu/paddress [12]),
    .d(\biu/bus_unit/mmu_hwdata [10]),
    .o(_al_u5987_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5988 (
    .a(_al_u2915_o),
    .b(_al_u5987_o),
    .o(_al_u5988_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*(D@C)))"),
    .INIT(16'hc44c))
    _al_u5989 (
    .a(\biu/maddress [12]),
    .b(_al_u5988_o),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u5989_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u5990 (
    .a(_al_u2915_o),
    .b(\biu/paddress [12]),
    .o(_al_u5990_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*~B)*~(A)*~(C)+~(~D*~B)*A*~(C)+~(~(~D*~B))*A*C+~(~D*~B)*A*C)"),
    .INIT(16'h5053))
    _al_u5991 (
    .a(_al_u5986_o),
    .b(_al_u5989_o),
    .c(_al_u2698_o),
    .d(_al_u5990_o),
    .o(\biu/bus_unit/mmu/n66 [12]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u5992 (
    .a(_al_u5157_o),
    .b(_al_u3190_o),
    .c(_al_u3184_o),
    .o(_al_u5992_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5993 (
    .a(_al_u5992_o),
    .b(_al_u3206_o),
    .o(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u5994 (
    .a(_al_u5157_o),
    .b(_al_u5108_o),
    .o(\cu_ru/m_s_status/u14_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u5995 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [9]),
    .d(\cu_ru/mtvec [9]),
    .o(\cu_ru/tvec [9]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u5996 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [8]),
    .d(\cu_ru/mtvec [8]),
    .o(\cu_ru/tvec [8]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u5997 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [7]),
    .d(\cu_ru/mtvec [7]),
    .o(\cu_ru/tvec [7]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u5998 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [63]),
    .d(\cu_ru/mtvec [63]),
    .o(\cu_ru/tvec [63]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u5999 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [62]),
    .d(\cu_ru/mtvec [62]),
    .o(\cu_ru/tvec [62]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6000 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [61]),
    .d(\cu_ru/mtvec [61]),
    .o(\cu_ru/tvec [61]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6001 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [60]),
    .d(\cu_ru/mtvec [60]),
    .o(\cu_ru/tvec [60]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6002 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [6]),
    .d(\cu_ru/mtvec [6]),
    .o(\cu_ru/tvec [6]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6003 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [59]),
    .d(\cu_ru/mtvec [59]),
    .o(\cu_ru/tvec [59]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6004 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [58]),
    .d(\cu_ru/mtvec [58]),
    .o(\cu_ru/tvec [58]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6005 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [57]),
    .d(\cu_ru/mtvec [57]),
    .o(\cu_ru/tvec [57]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6006 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [56]),
    .d(\cu_ru/mtvec [56]),
    .o(\cu_ru/tvec [56]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6007 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [55]),
    .d(\cu_ru/mtvec [55]),
    .o(\cu_ru/tvec [55]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6008 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [54]),
    .d(\cu_ru/mtvec [54]),
    .o(\cu_ru/tvec [54]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6009 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [53]),
    .d(\cu_ru/mtvec [53]),
    .o(\cu_ru/tvec [53]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6010 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [52]),
    .d(\cu_ru/mtvec [52]),
    .o(\cu_ru/tvec [52]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6011 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [51]),
    .d(\cu_ru/mtvec [51]),
    .o(\cu_ru/tvec [51]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6012 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [50]),
    .d(\cu_ru/mtvec [50]),
    .o(\cu_ru/tvec [50]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6013 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [5]),
    .d(\cu_ru/mtvec [5]),
    .o(\cu_ru/tvec [5]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6014 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [49]),
    .d(\cu_ru/mtvec [49]),
    .o(\cu_ru/tvec [49]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6015 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [48]),
    .d(\cu_ru/mtvec [48]),
    .o(\cu_ru/tvec [48]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6016 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [47]),
    .d(\cu_ru/mtvec [47]),
    .o(\cu_ru/tvec [47]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6017 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [46]),
    .d(\cu_ru/mtvec [46]),
    .o(\cu_ru/tvec [46]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6018 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [45]),
    .d(\cu_ru/mtvec [45]),
    .o(\cu_ru/tvec [45]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6019 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [44]),
    .d(\cu_ru/mtvec [44]),
    .o(\cu_ru/tvec [44]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6020 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [43]),
    .d(\cu_ru/mtvec [43]),
    .o(\cu_ru/tvec [43]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6021 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [42]),
    .d(\cu_ru/mtvec [42]),
    .o(\cu_ru/tvec [42]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6022 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [41]),
    .d(\cu_ru/mtvec [41]),
    .o(\cu_ru/tvec [41]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6023 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [40]),
    .d(\cu_ru/mtvec [40]),
    .o(\cu_ru/tvec [40]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6024 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [4]),
    .d(\cu_ru/mtvec [4]),
    .o(\cu_ru/tvec [4]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6025 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [39]),
    .d(\cu_ru/mtvec [39]),
    .o(\cu_ru/tvec [39]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6026 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [38]),
    .d(\cu_ru/mtvec [38]),
    .o(\cu_ru/tvec [38]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6027 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [37]),
    .d(\cu_ru/mtvec [37]),
    .o(\cu_ru/tvec [37]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6028 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [36]),
    .d(\cu_ru/mtvec [36]),
    .o(\cu_ru/tvec [36]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6029 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [35]),
    .d(\cu_ru/mtvec [35]),
    .o(\cu_ru/tvec [35]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6030 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [34]),
    .d(\cu_ru/mtvec [34]),
    .o(\cu_ru/tvec [34]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6031 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [33]),
    .d(\cu_ru/mtvec [33]),
    .o(\cu_ru/tvec [33]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6032 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [32]),
    .d(\cu_ru/mtvec [32]),
    .o(\cu_ru/tvec [32]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6033 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [31]),
    .d(\cu_ru/mtvec [31]),
    .o(\cu_ru/tvec [31]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6034 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [30]),
    .d(\cu_ru/mtvec [30]),
    .o(\cu_ru/tvec [30]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6035 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [29]),
    .d(\cu_ru/mtvec [29]),
    .o(\cu_ru/tvec [29]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6036 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [28]),
    .d(\cu_ru/mtvec [28]),
    .o(\cu_ru/tvec [28]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6037 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [27]),
    .d(\cu_ru/mtvec [27]),
    .o(\cu_ru/tvec [27]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6038 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [26]),
    .d(\cu_ru/mtvec [26]),
    .o(\cu_ru/tvec [26]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6039 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [25]),
    .d(\cu_ru/mtvec [25]),
    .o(\cu_ru/tvec [25]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6040 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [24]),
    .d(\cu_ru/mtvec [24]),
    .o(\cu_ru/tvec [24]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6041 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [23]),
    .d(\cu_ru/mtvec [23]),
    .o(\cu_ru/tvec [23]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6042 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [22]),
    .d(\cu_ru/mtvec [22]),
    .o(\cu_ru/tvec [22]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6043 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [21]),
    .d(\cu_ru/mtvec [21]),
    .o(\cu_ru/tvec [21]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6044 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [20]),
    .d(\cu_ru/mtvec [20]),
    .o(\cu_ru/tvec [20]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6045 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [19]),
    .d(\cu_ru/mtvec [19]),
    .o(\cu_ru/tvec [19]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6046 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [18]),
    .d(\cu_ru/mtvec [18]),
    .o(\cu_ru/tvec [18]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6047 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [17]),
    .d(\cu_ru/mtvec [17]),
    .o(\cu_ru/tvec [17]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6048 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [16]),
    .d(\cu_ru/mtvec [16]),
    .o(\cu_ru/tvec [16]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6049 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [15]),
    .d(\cu_ru/mtvec [15]),
    .o(\cu_ru/tvec [15]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6050 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [14]),
    .d(\cu_ru/mtvec [14]),
    .o(\cu_ru/tvec [14]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6051 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [13]),
    .d(\cu_ru/mtvec [13]),
    .o(\cu_ru/tvec [13]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6052 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [12]),
    .d(\cu_ru/mtvec [12]),
    .o(\cu_ru/tvec [12]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6053 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [11]),
    .d(\cu_ru/mtvec [11]),
    .o(\cu_ru/tvec [11]));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u6054 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [10]),
    .d(\cu_ru/mtvec [10]),
    .o(\cu_ru/tvec [10]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6055 (
    .a(\cu_ru/trap_target_m ),
    .b(_al_u5157_o),
    .o(_al_u6055_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u6056 (
    .a(_al_u6055_o),
    .b(pc_jmp),
    .o(pip_flush));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6057 (
    .a(\cu_ru/trap_target_m ),
    .b(rst_pad),
    .o(\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6058 (
    .a(_al_u3939_o),
    .b(id_ins[31]),
    .c(id_ins[30]),
    .o(_al_u6058_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u6059 (
    .a(\ins_dec/op_load ),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .d(_al_u3384_o),
    .o(_al_u6059_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u6060 (
    .a(_al_u4064_o),
    .b(_al_u3216_o),
    .c(_al_u3217_o),
    .d(_al_u6059_o),
    .o(\ins_dec/n198_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6061 (
    .a(\ins_dec/n198_lutinv ),
    .b(\ins_dec/funct7_32_lutinv ),
    .c(_al_u4801_o),
    .o(_al_u6061_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~B*A)"),
    .INIT(8'hdf))
    _al_u6062 (
    .a(_al_u4806_o),
    .b(_al_u6058_o),
    .c(_al_u6061_o),
    .o(\ins_dec/n206 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6063 (
    .a(rs1_data[55]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6063_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6064 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_055 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_055 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6064_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6065 (
    .a(_al_u3927_o),
    .b(id_ins[31]),
    .o(_al_u6065_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6066 (
    .a(_al_u6063_o),
    .b(_al_u6064_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [55]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6067 (
    .a(rs1_data[54]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6067_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6068 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_054 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_054 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6068_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6069 (
    .a(_al_u6067_o),
    .b(_al_u6068_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [54]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6070 (
    .a(rs1_data[53]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6070_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6071 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_053 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_053 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6071_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6072 (
    .a(_al_u6070_o),
    .b(_al_u6071_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [53]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6073 (
    .a(rs1_data[52]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6073_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6074 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_052 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_052 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6074_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6075 (
    .a(_al_u6073_o),
    .b(_al_u6074_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [52]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6076 (
    .a(rs1_data[51]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6076_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6077 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_051 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_051 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6077_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6078 (
    .a(_al_u6076_o),
    .b(_al_u6077_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [51]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6079 (
    .a(rs1_data[50]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6079_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6080 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_050 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_050 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6080_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6081 (
    .a(_al_u6079_o),
    .b(_al_u6080_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [50]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6082 (
    .a(rs1_data[49]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6082_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6083 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_049 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_049 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6083_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6084 (
    .a(_al_u6082_o),
    .b(_al_u6083_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [49]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6085 (
    .a(rs1_data[48]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6085_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6086 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_048 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_048 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6086_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6087 (
    .a(_al_u6085_o),
    .b(_al_u6086_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [48]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6088 (
    .a(rs1_data[47]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6088_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6089 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_047 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_047 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6089_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6090 (
    .a(_al_u6088_o),
    .b(_al_u6089_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [47]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6091 (
    .a(rs1_data[46]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6091_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6092 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_046 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_046 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6092_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6093 (
    .a(_al_u6091_o),
    .b(_al_u6092_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [46]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6094 (
    .a(rs1_data[45]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6094_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6095 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_045 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_045 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6095_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6096 (
    .a(_al_u6094_o),
    .b(_al_u6095_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [45]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6097 (
    .a(rs1_data[44]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6097_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6098 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_044 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_044 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6098_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6099 (
    .a(_al_u6097_o),
    .b(_al_u6098_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [44]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6100 (
    .a(rs1_data[43]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6100_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6101 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_043 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_043 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6101_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6102 (
    .a(_al_u6100_o),
    .b(_al_u6101_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [43]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6103 (
    .a(rs1_data[42]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6103_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6104 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_042 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_042 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6104_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6105 (
    .a(_al_u6103_o),
    .b(_al_u6104_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [42]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6106 (
    .a(rs1_data[41]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6106_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6107 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_041 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_041 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6107_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6108 (
    .a(_al_u6106_o),
    .b(_al_u6107_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [41]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6109 (
    .a(rs1_data[40]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6109_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6110 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_040 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_040 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6110_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6111 (
    .a(_al_u6109_o),
    .b(_al_u6110_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [40]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6112 (
    .a(\ins_dec/n239 ),
    .b(_al_u3216_o),
    .o(_al_u6112_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .INIT(16'h1d3f))
    _al_u6113 (
    .a(_al_u6112_o),
    .b(_al_u3927_o),
    .c(id_ins[24]),
    .d(id_ins[11]),
    .o(_al_u6113_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u6114 (
    .a(rs1_data[4]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u6113_o),
    .o(_al_u6114_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u6115 (
    .a(_al_u6114_o),
    .b(_al_u5839_o),
    .o(\ins_dec/n284 [4]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6116 (
    .a(rs1_data[39]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6116_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6117 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_039 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_039 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6117_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6118 (
    .a(_al_u6116_o),
    .b(_al_u6117_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [39]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6119 (
    .a(rs1_data[38]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6119_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6120 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_038 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_038 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6120_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6121 (
    .a(_al_u6119_o),
    .b(_al_u6120_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [38]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6122 (
    .a(rs1_data[37]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6122_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6123 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_037 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_037 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6123_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6124 (
    .a(_al_u6122_o),
    .b(_al_u6123_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [37]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6125 (
    .a(rs1_data[36]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6125_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6126 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_036 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_036 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6126_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6127 (
    .a(_al_u6125_o),
    .b(_al_u6126_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [36]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6128 (
    .a(rs1_data[35]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6128_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6129 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_035 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_035 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6129_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6130 (
    .a(_al_u6128_o),
    .b(_al_u6129_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [35]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6131 (
    .a(rs1_data[34]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6131_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6132 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_034 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_034 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6132_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6133 (
    .a(_al_u6131_o),
    .b(_al_u6132_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [34]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6134 (
    .a(rs1_data[33]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6134_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6135 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_033 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_033 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6135_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6136 (
    .a(_al_u6134_o),
    .b(_al_u6135_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [33]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6137 (
    .a(rs1_data[32]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6137_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6138 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_032 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_032 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6138_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6139 (
    .a(_al_u6137_o),
    .b(_al_u6138_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [32]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6140 (
    .a(rs1_data[31]),
    .b(_al_u5858_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6140_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6141 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_031 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_031 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6141_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6142 (
    .a(_al_u6140_o),
    .b(_al_u6141_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [31]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6143 (
    .a(rs1_data[30]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[30]),
    .o(_al_u6143_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6144 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_030 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_030 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6144_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6145 (
    .a(_al_u6143_o),
    .b(_al_u6144_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [30]));
  AL_MAP_LUT4 #(
    .EQN("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .INIT(16'h1d3f))
    _al_u6146 (
    .a(_al_u6112_o),
    .b(_al_u3927_o),
    .c(id_ins[23]),
    .d(id_ins[10]),
    .o(_al_u6146_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u6147 (
    .a(rs1_data[3]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u6146_o),
    .o(_al_u6147_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u6148 (
    .a(_al_u6147_o),
    .b(_al_u5841_o),
    .o(\ins_dec/n284 [3]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6149 (
    .a(rs1_data[29]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[29]),
    .o(_al_u6149_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6150 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_029 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_029 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6150_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6151 (
    .a(_al_u6149_o),
    .b(_al_u6150_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [29]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6152 (
    .a(rs1_data[28]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[28]),
    .o(_al_u6152_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6153 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_028 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_028 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6153_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6154 (
    .a(_al_u6152_o),
    .b(_al_u6153_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [28]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6155 (
    .a(rs1_data[27]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[27]),
    .o(_al_u6155_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6156 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_027 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_027 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6156_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6157 (
    .a(_al_u6155_o),
    .b(_al_u6156_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [27]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6158 (
    .a(rs1_data[26]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[26]),
    .o(_al_u6158_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6159 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_026 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_026 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6159_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6160 (
    .a(_al_u6158_o),
    .b(_al_u6159_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [26]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6161 (
    .a(rs1_data[25]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[25]),
    .o(_al_u6161_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6162 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_025 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_025 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6162_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6163 (
    .a(_al_u6161_o),
    .b(_al_u6162_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [25]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6164 (
    .a(rs1_data[24]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[24]),
    .o(_al_u6164_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6165 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_024 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_024 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6165_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6166 (
    .a(_al_u6164_o),
    .b(_al_u6165_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [24]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6167 (
    .a(rs1_data[23]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[23]),
    .o(_al_u6167_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6168 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_023 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_023 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6168_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6169 (
    .a(_al_u6167_o),
    .b(_al_u6168_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [23]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6170 (
    .a(rs1_data[22]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[22]),
    .o(_al_u6170_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6171 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_022 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_022 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6171_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6172 (
    .a(_al_u6170_o),
    .b(_al_u6171_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [22]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6173 (
    .a(rs1_data[21]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[21]),
    .o(_al_u6173_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6174 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_021 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_021 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6174_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6175 (
    .a(_al_u6173_o),
    .b(_al_u6174_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [21]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6176 (
    .a(rs1_data[20]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[20]),
    .o(_al_u6176_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6177 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_020 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_020 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6177_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6178 (
    .a(_al_u6176_o),
    .b(_al_u6177_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [20]));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~((~D*A))*~(B)+~C*(~D*A)*~(B)+~(~C)*(~D*A)*B+~C*(~D*A)*B)"),
    .INIT(16'hfc74))
    _al_u6179 (
    .a(rs1_data[2]),
    .b(\ins_dec/n239 ),
    .c(_al_u3955_o),
    .d(_al_u3216_o),
    .o(_al_u6179_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6180 (
    .a(_al_u6179_o),
    .b(_al_u6112_o),
    .c(id_ins[9]),
    .o(_al_u6180_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u6181 (
    .a(_al_u6180_o),
    .b(_al_u4086_o),
    .c(_al_u3927_o),
    .d(id_ins[22]),
    .o(_al_u6181_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u6182 (
    .a(_al_u6181_o),
    .b(_al_u5843_o),
    .o(\ins_dec/n284 [2]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6183 (
    .a(rs1_data[19]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[19]),
    .o(_al_u6183_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6184 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_019 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_019 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6184_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6185 (
    .a(_al_u6183_o),
    .b(_al_u6184_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [19]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6186 (
    .a(rs1_data[18]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[18]),
    .o(_al_u6186_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6187 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_018 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_018 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6187_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6188 (
    .a(_al_u6186_o),
    .b(_al_u6187_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [18]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6189 (
    .a(rs1_data[17]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[17]),
    .o(_al_u6189_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6190 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_017 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_017 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6190_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6191 (
    .a(_al_u6189_o),
    .b(_al_u6190_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [17]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6192 (
    .a(rs1_data[16]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[16]),
    .o(_al_u6192_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6193 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_016 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_016 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6193_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6194 (
    .a(_al_u6192_o),
    .b(_al_u6193_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [16]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6195 (
    .a(rs1_data[15]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(id_ins[15]),
    .o(_al_u6195_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6196 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_015 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_015 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6196_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6197 (
    .a(_al_u6195_o),
    .b(_al_u6196_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [15]));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(C)*~(D)+(B*A)*C*~(D)+~((B*A))*C*D+(B*A)*C*D)"),
    .INIT(16'h0f77))
    _al_u6198 (
    .a(rs1_data[14]),
    .b(\ins_dec/n239 ),
    .c(_al_u3955_o),
    .d(_al_u3216_o),
    .o(_al_u6198_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6199 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_014 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_014 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6199_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6200 (
    .a(_al_u6198_o),
    .b(_al_u6199_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [14]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6201 (
    .a(rs1_data[13]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(_al_u3217_o),
    .o(_al_u6201_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6202 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_013 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_013 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6202_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6203 (
    .a(_al_u6201_o),
    .b(_al_u6202_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [13]));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u6204 (
    .a(rs1_data[12]),
    .b(\ins_dec/mux19_b10_sel_is_2_o ),
    .c(_al_u3955_o),
    .d(_al_u3384_o),
    .o(_al_u6204_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u6205 (
    .a(_al_u5144_o),
    .b(\cu_ru/al_ram_gpr_al_u0_do_i0_012 ),
    .c(\cu_ru/al_ram_gpr_al_u0_do_i1_012 ),
    .d(\cu_ru/n49 [4]),
    .o(_al_u6205_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*A)"),
    .INIT(8'hfd))
    _al_u6206 (
    .a(_al_u6204_o),
    .b(_al_u6205_o),
    .c(_al_u6065_o),
    .o(\ins_dec/n284 [12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6207 (
    .a(_al_u4086_o),
    .b(_al_u3927_o),
    .c(id_ins[21]),
    .o(_al_u6207_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6208 (
    .a(_al_u6112_o),
    .b(_al_u6207_o),
    .c(id_ins[8]),
    .o(_al_u6208_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6209 (
    .a(rs1_data[1]),
    .b(_al_u6208_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6209_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u6210 (
    .a(_al_u6209_o),
    .b(_al_u5845_o),
    .c(_al_u4086_o),
    .o(\ins_dec/n284 [1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6211 (
    .a(_al_u4086_o),
    .b(_al_u3927_o),
    .c(id_ins[20]),
    .o(_al_u6211_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6212 (
    .a(_al_u6112_o),
    .b(_al_u6211_o),
    .c(id_ins[7]),
    .o(_al_u6212_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6213 (
    .a(rs1_data[0]),
    .b(_al_u6212_o),
    .c(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(_al_u6213_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u6214 (
    .a(_al_u6213_o),
    .b(_al_u5847_o),
    .c(_al_u4086_o),
    .o(\ins_dec/n284 [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6215 (
    .a(\biu/maddress [20]),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6215_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u6216 (
    .a(\biu/maddress [38]),
    .b(\biu/maddress [29]),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6216_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6217 (
    .a(_al_u6215_o),
    .b(_al_u6216_o),
    .c(_al_u3034_o),
    .d(\biu/paddress [75]),
    .o(\biu/bus_unit/mmu/n71 [11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6218 (
    .a(\biu/maddress [19]),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6218_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u6219 (
    .a(\biu/maddress [37]),
    .b(\biu/maddress [28]),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6219_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6220 (
    .a(_al_u6218_o),
    .b(_al_u6219_o),
    .c(_al_u3034_o),
    .d(\biu/paddress [74]),
    .o(\biu/bus_unit/mmu/n71 [10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6221 (
    .a(\biu/maddress [18]),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6221_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u6222 (
    .a(\biu/maddress [36]),
    .b(\biu/maddress [27]),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6222_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6223 (
    .a(_al_u6221_o),
    .b(_al_u6222_o),
    .c(_al_u3034_o),
    .d(\biu/paddress [73]),
    .o(\biu/bus_unit/mmu/n71 [9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6224 (
    .a(\biu/maddress [17]),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6224_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u6225 (
    .a(\biu/maddress [35]),
    .b(\biu/maddress [26]),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6225_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6226 (
    .a(_al_u6224_o),
    .b(_al_u6225_o),
    .c(_al_u3034_o),
    .d(\biu/paddress [72]),
    .o(\biu/bus_unit/mmu/n71 [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6227 (
    .a(\biu/maddress [16]),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6227_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u6228 (
    .a(\biu/maddress [34]),
    .b(\biu/maddress [25]),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6228_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6229 (
    .a(_al_u6227_o),
    .b(_al_u6228_o),
    .c(_al_u3034_o),
    .d(\biu/paddress [71]),
    .o(\biu/bus_unit/mmu/n71 [7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6230 (
    .a(\biu/maddress [15]),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6230_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u6231 (
    .a(\biu/maddress [33]),
    .b(\biu/maddress [24]),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6231_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6232 (
    .a(_al_u6230_o),
    .b(_al_u6231_o),
    .c(_al_u3034_o),
    .d(\biu/paddress [70]),
    .o(\biu/bus_unit/mmu/n71 [6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6233 (
    .a(\biu/maddress [14]),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6233_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u6234 (
    .a(\biu/maddress [32]),
    .b(\biu/maddress [23]),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6234_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6235 (
    .a(_al_u6233_o),
    .b(_al_u6234_o),
    .c(_al_u3034_o),
    .d(\biu/paddress [69]),
    .o(\biu/bus_unit/mmu/n71 [5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6236 (
    .a(\biu/maddress [13]),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6236_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u6237 (
    .a(\biu/maddress [31]),
    .b(\biu/maddress [22]),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6237_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6238 (
    .a(_al_u6236_o),
    .b(_al_u6237_o),
    .c(_al_u3034_o),
    .d(\biu/paddress [68]),
    .o(\biu/bus_unit/mmu/n71 [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6239 (
    .a(\biu/maddress [12]),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6239_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u6240 (
    .a(\biu/maddress [30]),
    .b(\biu/maddress [21]),
    .c(\biu/bus_unit/mmu/i [0]),
    .d(\biu/bus_unit/mmu/i [1]),
    .o(_al_u6240_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6241 (
    .a(_al_u6239_o),
    .b(_al_u6240_o),
    .c(_al_u3034_o),
    .d(\biu/paddress [67]),
    .o(\biu/bus_unit/mmu/n71 [3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u6242 (
    .a(\ins_dec/ins_fence ),
    .b(\ins_dec/op_store ),
    .c(_al_u4064_o),
    .o(\ins_dec/dec_gpr_write ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6243 (
    .a(\biu/cache_ctrl_logic/l1d_va [37]),
    .b(\biu/cache_ctrl_logic/l1d_va [56]),
    .c(addr_ex[37]),
    .d(addr_ex[56]),
    .o(_al_u6243_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u6244 (
    .a(_al_u6243_o),
    .b(\biu/cache_ctrl_logic/l1d_va [51]),
    .c(addr_ex[51]),
    .o(_al_u6244_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6245 (
    .a(\biu/cache_ctrl_logic/l1d_va [12]),
    .b(\biu/cache_ctrl_logic/l1d_va [20]),
    .c(addr_ex[12]),
    .d(addr_ex[20]),
    .o(_al_u6245_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u6246 (
    .a(_al_u6244_o),
    .b(_al_u6245_o),
    .c(\biu/cache_ctrl_logic/l1d_va [14]),
    .d(addr_ex[14]),
    .o(_al_u6246_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6247 (
    .a(\biu/cache_ctrl_logic/l1d_va [12]),
    .b(\biu/cache_ctrl_logic/l1d_va [20]),
    .c(addr_ex[12]),
    .d(addr_ex[20]),
    .o(_al_u6247_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u6248 (
    .a(_al_u6247_o),
    .b(\biu/cache_ctrl_logic/l1d_va [22]),
    .c(addr_ex[22]),
    .o(_al_u6248_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6249 (
    .a(\biu/cache_ctrl_logic/l1d_va [18]),
    .b(\biu/cache_ctrl_logic/l1d_va [36]),
    .c(addr_ex[18]),
    .d(addr_ex[36]),
    .o(_al_u6249_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6250 (
    .a(\biu/cache_ctrl_logic/l1d_va [46]),
    .b(\biu/cache_ctrl_logic/l1d_va [52]),
    .c(addr_ex[46]),
    .d(addr_ex[52]),
    .o(_al_u6250_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6251 (
    .a(_al_u6246_o),
    .b(_al_u6248_o),
    .c(_al_u6249_o),
    .d(_al_u6250_o),
    .o(_al_u6251_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*(D@B))"),
    .INIT(16'h0104))
    _al_u6252 (
    .a(\exu/main_state [0]),
    .b(\exu/main_state [1]),
    .c(\exu/main_state [2]),
    .d(\exu/main_state [3]),
    .o(\exu/n59_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6253 (
    .a(\exu/n59_lutinv ),
    .b(load),
    .o(read));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u6254 (
    .a(\exu/main_state [0]),
    .b(\exu/main_state [1]),
    .c(\exu/main_state [2]),
    .d(\exu/main_state [3]),
    .o(_al_u6254_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u6255 (
    .a(\exu/main_state [0]),
    .b(\exu/main_state [1]),
    .c(\exu/main_state [2]),
    .d(\exu/main_state [3]),
    .o(_al_u6255_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u6256 (
    .a(_al_u6254_o),
    .b(_al_u6255_o),
    .c(store),
    .o(write));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6257 (
    .a(read),
    .b(write),
    .o(_al_u6257_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6258 (
    .a(\biu/cache_ctrl_logic/l1d_value ),
    .b(\biu/cache_ctrl_logic/l1d_va [44]),
    .c(addr_ex[44]),
    .o(_al_u6258_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6259 (
    .a(\biu/cache_ctrl_logic/l1d_va [33]),
    .b(\biu/cache_ctrl_logic/l1d_va [60]),
    .c(addr_ex[33]),
    .d(addr_ex[60]),
    .o(_al_u6259_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u6260 (
    .a(_al_u6258_o),
    .b(_al_u6259_o),
    .c(\biu/cache_ctrl_logic/l1d_va [55]),
    .d(addr_ex[55]),
    .o(_al_u6260_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6261 (
    .a(\biu/cache_ctrl_logic/l1d_va [49]),
    .b(\biu/cache_ctrl_logic/l1d_va [63]),
    .c(addr_ex[49]),
    .d(addr_ex[63]),
    .o(_al_u6261_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6262 (
    .a(\biu/cache_ctrl_logic/l1d_va [62]),
    .b(\biu/cache_ctrl_logic/l1d_va [63]),
    .c(addr_ex[62]),
    .d(addr_ex[63]),
    .o(_al_u6262_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6263 (
    .a(\biu/cache_ctrl_logic/l1d_va [52]),
    .b(\biu/cache_ctrl_logic/l1d_va [57]),
    .c(addr_ex[52]),
    .d(addr_ex[57]),
    .o(_al_u6263_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6264 (
    .a(\biu/cache_ctrl_logic/l1d_va [49]),
    .b(\biu/cache_ctrl_logic/l1d_va [57]),
    .c(addr_ex[49]),
    .d(addr_ex[57]),
    .o(_al_u6264_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6265 (
    .a(_al_u6261_o),
    .b(_al_u6262_o),
    .c(_al_u6263_o),
    .d(_al_u6264_o),
    .o(_al_u6265_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u6266 (
    .a(\biu/cache_ctrl_logic/l1d_va [16]),
    .b(addr_ex[16]),
    .o(\biu/cache_ctrl_logic/eq1/xor_i0[4]_i1[4]_o_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6267 (
    .a(\biu/cache_ctrl_logic/l1d_va [31]),
    .b(\biu/cache_ctrl_logic/l1d_va [39]),
    .c(addr_ex[31]),
    .d(addr_ex[39]),
    .o(_al_u6267_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6268 (
    .a(\biu/cache_ctrl_logic/l1d_va [19]),
    .b(\biu/cache_ctrl_logic/l1d_va [29]),
    .c(addr_ex[19]),
    .d(addr_ex[29]),
    .o(_al_u6268_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6269 (
    .a(\biu/cache_ctrl_logic/l1d_va [21]),
    .b(\biu/cache_ctrl_logic/l1d_va [61]),
    .c(addr_ex[21]),
    .d(addr_ex[61]),
    .o(_al_u6269_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u6270 (
    .a(\biu/cache_ctrl_logic/eq1/xor_i0[4]_i1[4]_o_lutinv ),
    .b(_al_u6267_o),
    .c(_al_u6268_o),
    .d(_al_u6269_o),
    .o(_al_u6270_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6271 (
    .a(_al_u6260_o),
    .b(_al_u6265_o),
    .c(_al_u6270_o),
    .o(_al_u6271_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u6272 (
    .a(\biu/cache_ctrl_logic/l1d_va [27]),
    .b(addr_ex[27]),
    .o(_al_u6272_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6273 (
    .a(\biu/cache_ctrl_logic/l1d_va [15]),
    .b(\biu/cache_ctrl_logic/l1d_va [25]),
    .c(addr_ex[15]),
    .d(addr_ex[25]),
    .o(_al_u6273_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6274 (
    .a(\biu/cache_ctrl_logic/l1d_va [43]),
    .b(\biu/cache_ctrl_logic/l1d_va [46]),
    .c(addr_ex[43]),
    .d(addr_ex[46]),
    .o(_al_u6274_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6275 (
    .a(\biu/cache_ctrl_logic/l1d_va [42]),
    .b(\biu/cache_ctrl_logic/l1d_va [54]),
    .c(addr_ex[42]),
    .d(addr_ex[54]),
    .o(_al_u6275_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6276 (
    .a(_al_u6272_o),
    .b(_al_u6273_o),
    .c(_al_u6274_o),
    .d(_al_u6275_o),
    .o(_al_u6276_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6277 (
    .a(\biu/cache_ctrl_logic/l1d_va [34]),
    .b(\biu/cache_ctrl_logic/l1d_va [38]),
    .c(addr_ex[34]),
    .d(addr_ex[38]),
    .o(_al_u6277_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6278 (
    .a(\biu/cache_ctrl_logic/l1d_va [28]),
    .b(\biu/cache_ctrl_logic/l1d_va [32]),
    .c(addr_ex[28]),
    .d(addr_ex[32]),
    .o(_al_u6278_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6279 (
    .a(\biu/cache_ctrl_logic/l1d_va [23]),
    .b(\biu/cache_ctrl_logic/l1d_va [35]),
    .c(addr_ex[23]),
    .d(addr_ex[35]),
    .o(_al_u6279_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6280 (
    .a(_al_u6277_o),
    .b(_al_u6278_o),
    .c(_al_u6279_o),
    .o(_al_u6280_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6281 (
    .a(\biu/cache_ctrl_logic/l1d_va [18]),
    .b(\biu/cache_ctrl_logic/l1d_va [24]),
    .c(addr_ex[18]),
    .d(addr_ex[24]),
    .o(_al_u6281_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6282 (
    .a(\biu/cache_ctrl_logic/l1d_va [44]),
    .b(\biu/cache_ctrl_logic/l1d_va [56]),
    .c(addr_ex[44]),
    .d(addr_ex[56]),
    .o(_al_u6282_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6283 (
    .a(\biu/cache_ctrl_logic/l1d_va [48]),
    .b(\biu/cache_ctrl_logic/l1d_va [58]),
    .c(addr_ex[48]),
    .d(addr_ex[58]),
    .o(_al_u6283_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6284 (
    .a(\biu/cache_ctrl_logic/l1d_va [30]),
    .b(\biu/cache_ctrl_logic/l1d_va [48]),
    .c(addr_ex[30]),
    .d(addr_ex[48]),
    .o(_al_u6284_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6285 (
    .a(_al_u6281_o),
    .b(_al_u6282_o),
    .c(_al_u6283_o),
    .d(_al_u6284_o),
    .o(_al_u6285_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6286 (
    .a(\biu/cache_ctrl_logic/l1d_va [54]),
    .b(\biu/cache_ctrl_logic/l1d_va [58]),
    .c(addr_ex[54]),
    .d(addr_ex[58]),
    .o(_al_u6286_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6287 (
    .a(\biu/cache_ctrl_logic/l1d_va [43]),
    .b(\biu/cache_ctrl_logic/l1d_va [45]),
    .c(addr_ex[43]),
    .d(addr_ex[45]),
    .o(_al_u6287_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6288 (
    .a(\biu/cache_ctrl_logic/l1d_va [50]),
    .b(\biu/cache_ctrl_logic/l1d_va [59]),
    .c(addr_ex[50]),
    .d(addr_ex[59]),
    .o(_al_u6288_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6289 (
    .a(\biu/cache_ctrl_logic/l1d_va [45]),
    .b(\biu/cache_ctrl_logic/l1d_va [59]),
    .c(addr_ex[45]),
    .d(addr_ex[59]),
    .o(_al_u6289_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6290 (
    .a(_al_u6286_o),
    .b(_al_u6287_o),
    .c(_al_u6288_o),
    .d(_al_u6289_o),
    .o(_al_u6290_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6291 (
    .a(_al_u6276_o),
    .b(_al_u6280_o),
    .c(_al_u6285_o),
    .d(_al_u6290_o),
    .o(_al_u6291_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u6292 (
    .a(_al_u6257_o),
    .b(_al_u6271_o),
    .c(_al_u6291_o),
    .o(_al_u6292_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6293 (
    .a(\biu/cache_ctrl_logic/l1d_va [25]),
    .b(\biu/cache_ctrl_logic/l1d_va [53]),
    .c(addr_ex[25]),
    .d(addr_ex[53]),
    .o(_al_u6293_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u6294 (
    .a(_al_u6293_o),
    .b(\biu/cache_ctrl_logic/l1d_va [13]),
    .c(addr_ex[13]),
    .o(_al_u6294_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C@A))"),
    .INIT(16'h84a5))
    _al_u6295 (
    .a(\biu/cache_ctrl_logic/l1d_va [47]),
    .b(\biu/cache_ctrl_logic/l1d_va [53]),
    .c(addr_ex[47]),
    .d(addr_ex[53]),
    .o(_al_u6295_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6296 (
    .a(\biu/cache_ctrl_logic/l1d_va [41]),
    .b(\biu/cache_ctrl_logic/l1d_va [62]),
    .c(addr_ex[41]),
    .d(addr_ex[62]),
    .o(_al_u6296_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6297 (
    .a(\biu/cache_ctrl_logic/l1d_va [15]),
    .b(\biu/cache_ctrl_logic/l1d_va [41]),
    .c(addr_ex[15]),
    .d(addr_ex[41]),
    .o(_al_u6297_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6298 (
    .a(_al_u6294_o),
    .b(_al_u6295_o),
    .c(_al_u6296_o),
    .d(_al_u6297_o),
    .o(_al_u6298_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6299 (
    .a(\biu/cache_ctrl_logic/l1d_va [24]),
    .b(\biu/cache_ctrl_logic/l1d_va [36]),
    .c(addr_ex[24]),
    .d(addr_ex[36]),
    .o(_al_u6299_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u6300 (
    .a(_al_u6299_o),
    .b(\biu/cache_ctrl_logic/l1d_va [40]),
    .c(addr_ex[40]),
    .o(_al_u6300_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6301 (
    .a(\biu/cache_ctrl_logic/l1d_va [17]),
    .b(\biu/cache_ctrl_logic/l1d_va [26]),
    .c(addr_ex[17]),
    .d(addr_ex[26]),
    .o(_al_u6301_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6302 (
    .a(\biu/cache_ctrl_logic/l1d_va [30]),
    .b(\biu/cache_ctrl_logic/l1d_va [37]),
    .c(addr_ex[30]),
    .d(addr_ex[37]),
    .o(_al_u6302_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6303 (
    .a(\biu/cache_ctrl_logic/l1d_va [32]),
    .b(\biu/cache_ctrl_logic/l1d_va [50]),
    .c(addr_ex[32]),
    .d(addr_ex[50]),
    .o(_al_u6303_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6304 (
    .a(\biu/cache_ctrl_logic/l1d_va [17]),
    .b(\biu/cache_ctrl_logic/l1d_va [26]),
    .c(addr_ex[17]),
    .d(addr_ex[26]),
    .o(_al_u6304_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6305 (
    .a(_al_u6301_o),
    .b(_al_u6302_o),
    .c(_al_u6303_o),
    .d(_al_u6304_o),
    .o(_al_u6305_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6306 (
    .a(\biu/cache_ctrl_logic/l1d_va [34]),
    .b(\biu/cache_ctrl_logic/l1d_va [42]),
    .c(addr_ex[34]),
    .d(addr_ex[42]),
    .o(_al_u6306_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6307 (
    .a(\biu/cache_ctrl_logic/l1d_va [28]),
    .b(\biu/cache_ctrl_logic/l1d_va [38]),
    .c(addr_ex[28]),
    .d(addr_ex[38]),
    .o(_al_u6307_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6308 (
    .a(_al_u6300_o),
    .b(_al_u6305_o),
    .c(_al_u6306_o),
    .d(_al_u6307_o),
    .o(_al_u6308_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6309 (
    .a(_al_u6251_o),
    .b(_al_u6292_o),
    .c(_al_u6298_o),
    .d(_al_u6308_o),
    .o(_al_u6309_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(D*C)))"),
    .INIT(16'ha888))
    _al_u6310 (
    .a(read),
    .b(\biu/cache_ctrl_logic/l1i_pte [1]),
    .c(\biu/cache_ctrl_logic/l1d_pte [3]),
    .d(mxr),
    .o(\biu/cache_ctrl_logic/n42 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6311 (
    .a(\biu/cache_ctrl_logic/n42 ),
    .b(write),
    .c(\biu/cache_ctrl_logic/l1d_pte [2]),
    .o(_al_u6311_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(D*C)))"),
    .INIT(16'ha888))
    _al_u6312 (
    .a(read),
    .b(\biu/cache_ctrl_logic/l1d_pte [1]),
    .c(\biu/cache_ctrl_logic/l1d_pte [3]),
    .d(mxr),
    .o(\biu/cache_ctrl_logic/n34 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6313 (
    .a(priv[1]),
    .b(priv[3]),
    .o(_al_u6313_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6314 (
    .a(_al_u6313_o),
    .b(priv[0]),
    .o(\biu/bus_unit/mmu/n7_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6315 (
    .a(\biu/bus_unit/mmu/n7_lutinv ),
    .b(\biu/cache_ctrl_logic/l1d_pte [4]),
    .o(\biu/cache_ctrl_logic/n30 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D*C)))"),
    .INIT(16'hc888))
    _al_u6316 (
    .a(\biu/cache_ctrl_logic/n34 ),
    .b(\biu/cache_ctrl_logic/n30 ),
    .c(write),
    .d(\biu/cache_ctrl_logic/l1d_pte [2]),
    .o(\biu/cache_ctrl_logic/n36 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u6317 (
    .a(priv[0]),
    .b(priv[1]),
    .c(priv[3]),
    .o(\biu/bus_unit/mmu/n8_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6318 (
    .a(\biu/bus_unit/mmu/n8_lutinv ),
    .b(\biu/cache_ctrl_logic/l1d_pte [4]),
    .c(sum),
    .o(\biu/cache_ctrl_logic/n40 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6319 (
    .a(\biu/bus_unit/mmu/n31_lutinv ),
    .b(\cu_ru/m_s_status/n5 [1]),
    .c(priv[3]),
    .o(_al_u6319_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(C*~A))"),
    .INIT(16'h2300))
    _al_u6320 (
    .a(_al_u6311_o),
    .b(\biu/cache_ctrl_logic/n36 ),
    .c(\biu/cache_ctrl_logic/n40 ),
    .d(_al_u6319_o),
    .o(_al_u6320_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6321 (
    .a(_al_u6309_o),
    .b(_al_u6320_o),
    .o(_al_u6321_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6322 (
    .a(_al_u2703_o),
    .b(hready_pad),
    .c(\biu/bus_unit/statu [1]),
    .d(\biu/bus_unit/statu [3]),
    .o(\biu/cache_write_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u6323 (
    .a(_al_u6321_o),
    .b(\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ),
    .c(write),
    .d(\biu/cache_write_lutinv ),
    .o(_al_u6323_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u6324 (
    .a(_al_u3415_o),
    .b(ex_size[2]),
    .c(ex_size[3]),
    .o(\biu/cache_ctrl_logic/n176_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u6325 (
    .a(ex_size[0]),
    .b(ex_size[1]),
    .c(ex_size[2]),
    .d(ex_size[3]),
    .o(\biu/cache_ctrl_logic/n174_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6326 (
    .a(\biu/cache_ctrl_logic/n176_lutinv ),
    .b(\biu/cache_ctrl_logic/n174_lutinv ),
    .o(_al_u6326_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u6327 (
    .a(_al_u6326_o),
    .b(\exu/lsu/n0_lutinv ),
    .c(addr_ex[2]),
    .o(\biu/cache_ctrl_logic/n185 [3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6328 (
    .a(\exu/lsu/n0_lutinv ),
    .b(addr_ex[2]),
    .o(\biu/cache_ctrl_logic/n172_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u6329 (
    .a(\biu/cache_ctrl_logic/n172_lutinv ),
    .b(_al_u3415_o),
    .c(ex_size[2]),
    .d(ex_size[3]),
    .o(\biu/cache_ctrl_logic/n189 [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6330 (
    .a(addr_ex[0]),
    .b(addr_ex[1]),
    .o(\exu/lsu/n5_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u6331 (
    .a(\biu/cache_ctrl_logic/n189 [6]),
    .b(\biu/cache_ctrl_logic/n176_lutinv ),
    .c(\exu/lsu/n5_lutinv ),
    .d(addr_ex[2]),
    .o(_al_u6331_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u6332 (
    .a(\biu/cache_ctrl_logic/n176_lutinv ),
    .b(\exu/lsu/n8_lutinv ),
    .c(addr_ex[2]),
    .o(\biu/cache_ctrl_logic/n189 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u6333 (
    .a(ex_size[0]),
    .b(ex_size[1]),
    .c(ex_size[2]),
    .d(ex_size[3]),
    .o(\biu/cache_ctrl_logic/n173_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6334 (
    .a(\biu/cache_ctrl_logic/n174_lutinv ),
    .b(\biu/cache_ctrl_logic/n173_lutinv ),
    .o(_al_u6334_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u6335 (
    .a(_al_u6334_o),
    .b(\exu/lsu/n2_lutinv ),
    .c(addr_ex[2]),
    .o(\biu/cache_ctrl_logic/n182 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u6336 (
    .a(\biu/cache_ctrl_logic/n185 [3]),
    .b(_al_u6331_o),
    .c(\biu/cache_ctrl_logic/n189 [2]),
    .d(\biu/cache_ctrl_logic/n182 [4]),
    .o(_al_u6336_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6337 (
    .a(_al_u6323_o),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6336_o),
    .o(\biu/cache/n11 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u6338 (
    .a(_al_u6326_o),
    .b(\exu/lsu/n8_lutinv ),
    .c(addr_ex[2]),
    .o(\biu/cache_ctrl_logic/n185 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6339 (
    .a(\biu/cache_ctrl_logic/n176_lutinv ),
    .b(_al_u6334_o),
    .o(_al_u6339_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*B*~(D)+~(A)*~(B)*D+A*~(B)*D))"),
    .INIT(16'h0308))
    _al_u6340 (
    .a(\biu/cache_ctrl_logic/n176_lutinv ),
    .b(addr_ex[0]),
    .c(addr_ex[1]),
    .d(addr_ex[2]),
    .o(_al_u6340_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*~C))"),
    .INIT(16'h2022))
    _al_u6341 (
    .a(_al_u6331_o),
    .b(\biu/cache_ctrl_logic/n185 [2]),
    .c(_al_u6339_o),
    .d(_al_u6340_o),
    .o(_al_u6341_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6342 (
    .a(_al_u6323_o),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6341_o),
    .o(\biu/cache/n9 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u6343 (
    .a(_al_u6339_o),
    .b(\exu/lsu/n8_lutinv ),
    .c(addr_ex[2]),
    .o(\biu/cache_ctrl_logic/n182 [2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u6344 (
    .a(\biu/cache_ctrl_logic/n176_lutinv ),
    .b(addr_ex[1]),
    .c(addr_ex[2]),
    .o(_al_u6344_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*(D@C))"),
    .INIT(16'h0880))
    _al_u6345 (
    .a(\biu/cache_ctrl_logic/n172_lutinv ),
    .b(_al_u3415_o),
    .c(ex_size[2]),
    .d(ex_size[3]),
    .o(\biu/cache_ctrl_logic/n189 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(C*~B))"),
    .INIT(16'h0045))
    _al_u6346 (
    .a(\biu/cache_ctrl_logic/n182 [2]),
    .b(_al_u6326_o),
    .c(_al_u6344_o),
    .d(\biu/cache_ctrl_logic/n189 [5]),
    .o(_al_u6346_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6347 (
    .a(_al_u6323_o),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6346_o),
    .o(\biu/cache/n7 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*C*~A))"),
    .INIT(16'h3323))
    _al_u6348 (
    .a(_al_u6326_o),
    .b(\biu/cache_ctrl_logic/n189 [5]),
    .c(\exu/lsu/n2_lutinv ),
    .d(addr_ex[2]),
    .o(_al_u6348_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*~B))"),
    .INIT(16'haa8a))
    _al_u6349 (
    .a(_al_u6348_o),
    .b(_al_u6339_o),
    .c(\exu/lsu/n5_lutinv ),
    .d(addr_ex[2]),
    .o(_al_u6349_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6350 (
    .a(_al_u6323_o),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6349_o),
    .o(\biu/cache/n5 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u6351 (
    .a(_al_u6326_o),
    .b(\biu/cache_ctrl_logic/n189 [6]),
    .c(\biu/cache_ctrl_logic/n172_lutinv ),
    .o(_al_u6351_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*~B))"),
    .INIT(16'haa8a))
    _al_u6352 (
    .a(_al_u6351_o),
    .b(_al_u6339_o),
    .c(\exu/lsu/n2_lutinv ),
    .d(addr_ex[2]),
    .o(_al_u6352_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6353 (
    .a(_al_u6323_o),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6352_o),
    .o(\biu/cache/n3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfee9))
    _al_u6354 (
    .a(ex_size[0]),
    .b(ex_size[1]),
    .c(ex_size[2]),
    .d(ex_size[3]),
    .o(_al_u6354_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6355 (
    .a(\biu/cache_ctrl_logic/n172_lutinv ),
    .b(_al_u6354_o),
    .o(\biu/cache_ctrl_logic/ex_bsel [0]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6356 (
    .a(_al_u6323_o),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(\biu/cache_ctrl_logic/ex_bsel [0]),
    .o(\biu/cache/n1 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u6357 (
    .a(\biu/cache_ctrl_logic/n189 [6]),
    .b(\biu/cache_ctrl_logic/n176_lutinv ),
    .c(\exu/lsu/n0_lutinv ),
    .d(addr_ex[2]),
    .o(_al_u6357_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6358 (
    .a(\exu/lsu/n5_lutinv ),
    .b(\biu/cache_ctrl_logic/n174_lutinv ),
    .c(addr_ex[2]),
    .o(\biu/cache_ctrl_logic/n185 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u6359 (
    .a(\biu/cache_ctrl_logic/n185 [5]),
    .b(\exu/lsu/n8_lutinv ),
    .c(\biu/cache_ctrl_logic/n173_lutinv ),
    .d(addr_ex[2]),
    .o(_al_u6359_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6360 (
    .a(_al_u6357_o),
    .b(_al_u6359_o),
    .o(_al_u6360_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6361 (
    .a(_al_u6323_o),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6360_o),
    .o(\biu/cache/n15 ));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*B*~(C)+~(A)*~(B)*C+A*~(B)*C))"),
    .INIT(16'h3800))
    _al_u6362 (
    .a(\biu/cache_ctrl_logic/n174_lutinv ),
    .b(addr_ex[0]),
    .c(addr_ex[1]),
    .d(addr_ex[2]),
    .o(_al_u6362_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*~C))"),
    .INIT(16'h2022))
    _al_u6363 (
    .a(_al_u6357_o),
    .b(\biu/cache_ctrl_logic/n189 [2]),
    .c(_al_u6334_o),
    .d(_al_u6362_o),
    .o(_al_u6363_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6364 (
    .a(_al_u6323_o),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6363_o),
    .o(\biu/cache/n13 ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u6365 (
    .a(\biu/cache_ctrl_logic/l1i_va [48]),
    .b(addr_ex[48]),
    .o(_al_u6365_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6366 (
    .a(\biu/cache_ctrl_logic/l1i_va [38]),
    .b(\biu/cache_ctrl_logic/l1i_va [63]),
    .c(addr_ex[38]),
    .d(addr_ex[63]),
    .o(_al_u6366_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6367 (
    .a(\biu/cache_ctrl_logic/l1i_va [13]),
    .b(\biu/cache_ctrl_logic/l1i_va [25]),
    .c(addr_ex[13]),
    .d(addr_ex[25]),
    .o(_al_u6367_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6368 (
    .a(\biu/cache_ctrl_logic/l1i_va [18]),
    .b(\biu/cache_ctrl_logic/l1i_va [24]),
    .c(addr_ex[18]),
    .d(addr_ex[24]),
    .o(_al_u6368_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6369 (
    .a(_al_u6365_o),
    .b(_al_u6366_o),
    .c(_al_u6367_o),
    .d(_al_u6368_o),
    .o(_al_u6369_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6370 (
    .a(\biu/cache_ctrl_logic/l1i_va [62]),
    .b(\biu/cache_ctrl_logic/l1i_va [63]),
    .c(addr_ex[62]),
    .d(addr_ex[63]),
    .o(_al_u6370_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u6371 (
    .a(_al_u6369_o),
    .b(_al_u6370_o),
    .c(\biu/cache_ctrl_logic/l1i_va [58]),
    .d(addr_ex[58]),
    .o(_al_u6371_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6372 (
    .a(\biu/cache_ctrl_logic/l1i_va [13]),
    .b(\biu/cache_ctrl_logic/l1i_va [15]),
    .c(addr_ex[13]),
    .d(addr_ex[15]),
    .o(_al_u6372_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u6373 (
    .a(_al_u6372_o),
    .b(\biu/cache_ctrl_logic/l1i_va [33]),
    .c(addr_ex[33]),
    .o(_al_u6373_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6374 (
    .a(\biu/cache_ctrl_logic/l1i_va [15]),
    .b(\biu/cache_ctrl_logic/l1i_va [25]),
    .c(addr_ex[15]),
    .d(addr_ex[25]),
    .o(_al_u6374_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u6375 (
    .a(_al_u6374_o),
    .b(\biu/cache_ctrl_logic/l1i_va [47]),
    .c(addr_ex[47]),
    .o(_al_u6375_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6376 (
    .a(\biu/cache_ctrl_logic/l1i_va [23]),
    .b(\biu/cache_ctrl_logic/l1i_va [53]),
    .c(addr_ex[23]),
    .d(addr_ex[53]),
    .o(_al_u6376_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6377 (
    .a(\biu/cache_ctrl_logic/l1i_va [27]),
    .b(\biu/cache_ctrl_logic/l1i_va [35]),
    .c(addr_ex[27]),
    .d(addr_ex[35]),
    .o(_al_u6377_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6378 (
    .a(_al_u6373_o),
    .b(_al_u6375_o),
    .c(_al_u6376_o),
    .d(_al_u6377_o),
    .o(_al_u6378_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6379 (
    .a(\biu/cache_ctrl_logic/l1i_va [42]),
    .b(\biu/cache_ctrl_logic/l1i_va [43]),
    .c(addr_ex[42]),
    .d(addr_ex[43]),
    .o(_al_u6379_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u6380 (
    .a(_al_u6379_o),
    .b(\biu/cache_ctrl_logic/l1i_va [57]),
    .c(addr_ex[57]),
    .o(_al_u6380_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6381 (
    .a(\biu/cache_ctrl_logic/l1i_va [43]),
    .b(\biu/cache_ctrl_logic/l1i_va [45]),
    .c(addr_ex[43]),
    .d(addr_ex[45]),
    .o(_al_u6381_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u6382 (
    .a(_al_u6380_o),
    .b(_al_u6381_o),
    .c(\biu/cache_ctrl_logic/l1i_va [59]),
    .d(addr_ex[59]),
    .o(_al_u6382_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6383 (
    .a(\biu/cache_ctrl_logic/l1i_va [44]),
    .b(\biu/cache_ctrl_logic/l1i_va [46]),
    .c(addr_ex[44]),
    .d(addr_ex[46]),
    .o(_al_u6383_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6384 (
    .a(\biu/cache_ctrl_logic/l1i_va [50]),
    .b(\biu/cache_ctrl_logic/l1i_va [54]),
    .c(addr_ex[50]),
    .d(addr_ex[54]),
    .o(_al_u6384_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6385 (
    .a(\biu/cache_ctrl_logic/l1i_va [45]),
    .b(\biu/cache_ctrl_logic/l1i_va [58]),
    .c(addr_ex[45]),
    .d(addr_ex[58]),
    .o(_al_u6385_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6386 (
    .a(\biu/cache_ctrl_logic/l1i_va [54]),
    .b(\biu/cache_ctrl_logic/l1i_va [56]),
    .c(addr_ex[54]),
    .d(addr_ex[56]),
    .o(_al_u6386_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6387 (
    .a(_al_u6383_o),
    .b(_al_u6384_o),
    .c(_al_u6385_o),
    .d(_al_u6386_o),
    .o(_al_u6387_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6388 (
    .a(_al_u6371_o),
    .b(_al_u6378_o),
    .c(_al_u6382_o),
    .d(_al_u6387_o),
    .o(_al_u6388_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6389 (
    .a(\biu/cache_ctrl_logic/l1i_value ),
    .b(\biu/cache_ctrl_logic/l1i_va [12]),
    .c(addr_ex[12]),
    .o(_al_u6389_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6390 (
    .a(\biu/cache_ctrl_logic/l1i_va [21]),
    .b(\biu/cache_ctrl_logic/l1i_va [39]),
    .c(addr_ex[21]),
    .d(addr_ex[39]),
    .o(_al_u6390_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u6391 (
    .a(_al_u6389_o),
    .b(_al_u6390_o),
    .c(\biu/cache_ctrl_logic/l1i_va [16]),
    .d(addr_ex[16]),
    .o(_al_u6391_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6392 (
    .a(\biu/cache_ctrl_logic/l1i_va [14]),
    .b(\biu/cache_ctrl_logic/l1i_va [22]),
    .c(addr_ex[14]),
    .d(addr_ex[22]),
    .o(_al_u6392_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6393 (
    .a(\biu/cache_ctrl_logic/l1i_va [12]),
    .b(\biu/cache_ctrl_logic/l1i_va [20]),
    .c(addr_ex[12]),
    .d(addr_ex[20]),
    .o(_al_u6393_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6394 (
    .a(\biu/cache_ctrl_logic/l1i_va [20]),
    .b(\biu/cache_ctrl_logic/l1i_va [52]),
    .c(addr_ex[20]),
    .d(addr_ex[52]),
    .o(_al_u6394_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6395 (
    .a(_al_u6391_o),
    .b(_al_u6392_o),
    .c(_al_u6393_o),
    .d(_al_u6394_o),
    .o(_al_u6395_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6396 (
    .a(\biu/cache_ctrl_logic/l1i_va [37]),
    .b(\biu/cache_ctrl_logic/l1i_va [61]),
    .c(addr_ex[37]),
    .d(addr_ex[61]),
    .o(_al_u6396_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u6397 (
    .a(_al_u6396_o),
    .b(\biu/cache_ctrl_logic/l1i_va [60]),
    .c(addr_ex[60]),
    .o(_al_u6397_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6398 (
    .a(\biu/cache_ctrl_logic/l1i_va [31]),
    .b(\biu/cache_ctrl_logic/l1i_va [55]),
    .c(addr_ex[31]),
    .d(addr_ex[55]),
    .o(_al_u6398_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u6399 (
    .a(\biu/cache_ctrl_logic/l1i_va [19]),
    .b(\biu/cache_ctrl_logic/l1i_va [41]),
    .c(addr_ex[19]),
    .d(addr_ex[41]),
    .o(_al_u6399_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6400 (
    .a(_al_u6395_o),
    .b(_al_u6397_o),
    .c(_al_u6398_o),
    .d(_al_u6399_o),
    .o(_al_u6400_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6401 (
    .a(\biu/cache_ctrl_logic/l1i_va [29]),
    .b(\biu/cache_ctrl_logic/l1i_va [56]),
    .c(addr_ex[29]),
    .d(addr_ex[56]),
    .o(_al_u6401_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u6402 (
    .a(_al_u6401_o),
    .b(\biu/cache_ctrl_logic/l1i_va [51]),
    .c(addr_ex[51]),
    .o(_al_u6402_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6403 (
    .a(\biu/cache_ctrl_logic/l1i_va [44]),
    .b(\biu/cache_ctrl_logic/l1i_va [52]),
    .c(addr_ex[44]),
    .d(addr_ex[52]),
    .o(_al_u6403_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u6404 (
    .a(_al_u6402_o),
    .b(_al_u6403_o),
    .c(\biu/cache_ctrl_logic/l1i_va [49]),
    .d(addr_ex[49]),
    .o(_al_u6404_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6405 (
    .a(\biu/cache_ctrl_logic/l1i_va [30]),
    .b(\biu/cache_ctrl_logic/l1i_va [34]),
    .c(addr_ex[30]),
    .d(addr_ex[34]),
    .o(_al_u6405_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6406 (
    .a(\biu/cache_ctrl_logic/l1i_va [36]),
    .b(\biu/cache_ctrl_logic/l1i_va [40]),
    .c(addr_ex[36]),
    .d(addr_ex[40]),
    .o(_al_u6406_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6407 (
    .a(\biu/cache_ctrl_logic/l1i_va [18]),
    .b(\biu/cache_ctrl_logic/l1i_va [32]),
    .c(addr_ex[18]),
    .d(addr_ex[32]),
    .o(_al_u6407_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6408 (
    .a(\biu/cache_ctrl_logic/l1i_va [46]),
    .b(\biu/cache_ctrl_logic/l1i_va [62]),
    .c(addr_ex[46]),
    .d(addr_ex[62]),
    .o(_al_u6408_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6409 (
    .a(_al_u6405_o),
    .b(_al_u6406_o),
    .c(_al_u6407_o),
    .d(_al_u6408_o),
    .o(_al_u6409_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6410 (
    .a(\biu/cache_ctrl_logic/l1i_va [26]),
    .b(\biu/cache_ctrl_logic/l1i_va [32]),
    .c(addr_ex[26]),
    .d(addr_ex[32]),
    .o(_al_u6410_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u6411 (
    .a(_al_u6410_o),
    .b(\biu/cache_ctrl_logic/l1i_va [28]),
    .c(addr_ex[28]),
    .o(_al_u6411_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6412 (
    .a(\biu/cache_ctrl_logic/l1i_va [30]),
    .b(\biu/cache_ctrl_logic/l1i_va [42]),
    .c(addr_ex[30]),
    .d(addr_ex[42]),
    .o(_al_u6412_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u6413 (
    .a(\biu/cache_ctrl_logic/l1i_va [26]),
    .b(\biu/cache_ctrl_logic/l1i_va [36]),
    .c(addr_ex[26]),
    .d(addr_ex[36]),
    .o(_al_u6413_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6414 (
    .a(_al_u6409_o),
    .b(_al_u6411_o),
    .c(_al_u6412_o),
    .d(_al_u6413_o),
    .o(_al_u6414_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u6415 (
    .a(\biu/cache_ctrl_logic/l1i_va [17]),
    .b(\biu/cache_ctrl_logic/l1i_va [34]),
    .c(addr_ex[17]),
    .d(addr_ex[34]),
    .o(_al_u6415_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6416 (
    .a(\biu/cache_ctrl_logic/l1i_va [29]),
    .b(\biu/cache_ctrl_logic/l1i_va [38]),
    .c(addr_ex[29]),
    .d(addr_ex[38]),
    .o(_al_u6416_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u6417 (
    .a(\biu/cache_ctrl_logic/l1i_va [40]),
    .b(\biu/cache_ctrl_logic/l1i_va [50]),
    .c(addr_ex[40]),
    .d(addr_ex[50]),
    .o(_al_u6417_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u6418 (
    .a(\biu/cache_ctrl_logic/l1i_va [17]),
    .b(\biu/cache_ctrl_logic/l1i_va [24]),
    .c(addr_ex[17]),
    .d(addr_ex[24]),
    .o(_al_u6418_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6419 (
    .a(_al_u6415_o),
    .b(_al_u6416_o),
    .c(_al_u6417_o),
    .d(_al_u6418_o),
    .o(_al_u6419_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6420 (
    .a(_al_u6404_o),
    .b(_al_u6414_o),
    .c(_al_u6419_o),
    .o(_al_u6420_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u6421 (
    .a(_al_u6388_o),
    .b(_al_u6400_o),
    .c(_al_u6420_o),
    .d(_al_u6257_o),
    .o(\biu/cache_ctrl_logic/ex_l1i_hit ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(D*C)))"),
    .INIT(16'ha888))
    _al_u6422 (
    .a(read),
    .b(\biu/cache_ctrl_logic/l1i_pte [1]),
    .c(\biu/cache_ctrl_logic/l1i_pte [3]),
    .d(mxr),
    .o(\biu/cache_ctrl_logic/n17 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h1353))
    _al_u6423 (
    .a(\biu/bus_unit/mmu/n7_lutinv ),
    .b(\biu/bus_unit/mmu/n8_lutinv ),
    .c(\biu/cache_ctrl_logic/l1i_pte [4]),
    .d(sum),
    .o(_al_u6423_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~A*~(D*C)))"),
    .INIT(16'h3222))
    _al_u6424 (
    .a(\biu/cache_ctrl_logic/n17 ),
    .b(_al_u6423_o),
    .c(write),
    .d(\biu/cache_ctrl_logic/l1i_pte [2]),
    .o(\biu/cache_ctrl_logic/n26_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6425 (
    .a(\biu/cache_ctrl_logic/n26_lutinv ),
    .b(_al_u6319_o),
    .o(_al_u6425_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6426 (
    .a(\biu/cache_ctrl_logic/ex_l1i_hit ),
    .b(_al_u6425_o),
    .c(write),
    .o(_al_u6426_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u6427 (
    .a(_al_u6426_o),
    .b(_al_u2886_o),
    .c(\biu/cache_write_lutinv ),
    .o(\biu/l1i_write_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6428 (
    .a(\biu/l1i_write_lutinv ),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6360_o),
    .o(\biu/cache/n31 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6429 (
    .a(\biu/l1i_write_lutinv ),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6363_o),
    .o(\biu/cache/n29 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6430 (
    .a(\biu/l1i_write_lutinv ),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6336_o),
    .o(\biu/cache/n27 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6431 (
    .a(\biu/l1i_write_lutinv ),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6341_o),
    .o(\biu/cache/n25 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6432 (
    .a(\biu/l1i_write_lutinv ),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6346_o),
    .o(\biu/cache/n23 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6433 (
    .a(\biu/l1i_write_lutinv ),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6349_o),
    .o(\biu/cache/n21 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6434 (
    .a(\biu/l1i_write_lutinv ),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(_al_u6352_o),
    .o(\biu/cache/n19 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u6435 (
    .a(\biu/l1i_write_lutinv ),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(\biu/cache_ctrl_logic/ex_bsel [0]),
    .o(\biu/cache/n17 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*~B)))"),
    .INIT(16'haa20))
    _al_u6436 (
    .a(_al_u4122_o),
    .b(_al_u4107_o),
    .c(_al_u4127_o),
    .d(_al_u4128_o),
    .o(_al_u6436_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u6437 (
    .a(\cu_ru/mideleg_int_ctrl/sei_ack_m ),
    .b(\cu_ru/m_s_status/n5 [1]),
    .c(_al_u3244_o),
    .d(\cu_ru/mstatus [1]),
    .o(\cu_ru/mideleg_int_ctrl/n33_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~(~C*B)))"),
    .INIT(16'h5504))
    _al_u6438 (
    .a(_al_u4138_o),
    .b(\cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ),
    .c(\cu_ru/mideleg_int_ctrl/n33_neg_lutinv ),
    .d(_al_u4139_o),
    .o(_al_u6438_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(B*~(~D*~A)))"),
    .INIT(16'hfcf8))
    _al_u6439 (
    .a(_al_u6436_o),
    .b(_al_u4142_o),
    .c(_al_u6438_o),
    .d(_al_u4143_o),
    .o(\cu_ru/trap_cause [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6440 (
    .a(_al_u5992_o),
    .b(_al_u3204_o),
    .o(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6441 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [9]),
    .d(data_csr[9]),
    .o(_al_u6441_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6442 (
    .a(_al_u6441_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [9]),
    .o(\cu_ru/m_s_tval/n11 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6443 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [8]),
    .d(data_csr[8]),
    .o(_al_u6443_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6444 (
    .a(_al_u6443_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [8]),
    .o(\cu_ru/m_s_tval/n11 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6445 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [7]),
    .d(data_csr[7]),
    .o(_al_u6445_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6446 (
    .a(_al_u6445_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [7]),
    .o(\cu_ru/m_s_tval/n11 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6447 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [6]),
    .d(data_csr[6]),
    .o(_al_u6447_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6448 (
    .a(_al_u6447_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [6]),
    .o(\cu_ru/m_s_tval/n11 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6449 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [63]),
    .d(data_csr[63]),
    .o(_al_u6449_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6450 (
    .a(_al_u6449_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [63]),
    .o(\cu_ru/m_s_tval/n11 [63]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6451 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [62]),
    .d(data_csr[62]),
    .o(_al_u6451_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6452 (
    .a(_al_u6451_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [62]),
    .o(\cu_ru/m_s_tval/n11 [62]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6453 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [61]),
    .d(data_csr[61]),
    .o(_al_u6453_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6454 (
    .a(_al_u6453_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [61]),
    .o(\cu_ru/m_s_tval/n11 [61]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6455 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [60]),
    .d(data_csr[60]),
    .o(_al_u6455_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6456 (
    .a(_al_u6455_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [60]),
    .o(\cu_ru/m_s_tval/n11 [60]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6457 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [5]),
    .d(data_csr[5]),
    .o(_al_u6457_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6458 (
    .a(_al_u6457_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [5]),
    .o(\cu_ru/m_s_tval/n11 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6459 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [59]),
    .d(data_csr[59]),
    .o(_al_u6459_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6460 (
    .a(_al_u6459_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [59]),
    .o(\cu_ru/m_s_tval/n11 [59]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6461 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [58]),
    .d(data_csr[58]),
    .o(_al_u6461_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6462 (
    .a(_al_u6461_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [58]),
    .o(\cu_ru/m_s_tval/n11 [58]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6463 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [57]),
    .d(data_csr[57]),
    .o(_al_u6463_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6464 (
    .a(_al_u6463_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [57]),
    .o(\cu_ru/m_s_tval/n11 [57]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6465 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [56]),
    .d(data_csr[56]),
    .o(_al_u6465_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6466 (
    .a(_al_u6465_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [56]),
    .o(\cu_ru/m_s_tval/n11 [56]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6467 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [55]),
    .d(data_csr[55]),
    .o(_al_u6467_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6468 (
    .a(_al_u6467_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [55]),
    .o(\cu_ru/m_s_tval/n11 [55]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6469 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [54]),
    .d(data_csr[54]),
    .o(_al_u6469_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6470 (
    .a(_al_u6469_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [54]),
    .o(\cu_ru/m_s_tval/n11 [54]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6471 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [53]),
    .d(data_csr[53]),
    .o(_al_u6471_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6472 (
    .a(_al_u6471_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [53]),
    .o(\cu_ru/m_s_tval/n11 [53]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6473 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [52]),
    .d(data_csr[52]),
    .o(_al_u6473_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6474 (
    .a(_al_u6473_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [52]),
    .o(\cu_ru/m_s_tval/n11 [52]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6475 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [51]),
    .d(data_csr[51]),
    .o(_al_u6475_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6476 (
    .a(_al_u6475_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [51]),
    .o(\cu_ru/m_s_tval/n11 [51]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6477 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [50]),
    .d(data_csr[50]),
    .o(_al_u6477_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6478 (
    .a(_al_u6477_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [50]),
    .o(\cu_ru/m_s_tval/n11 [50]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6479 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [4]),
    .d(data_csr[4]),
    .o(_al_u6479_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6480 (
    .a(_al_u6479_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [4]),
    .o(\cu_ru/m_s_tval/n11 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6481 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [49]),
    .d(data_csr[49]),
    .o(_al_u6481_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6482 (
    .a(_al_u6481_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [49]),
    .o(\cu_ru/m_s_tval/n11 [49]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6483 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [48]),
    .d(data_csr[48]),
    .o(_al_u6483_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6484 (
    .a(_al_u6483_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [48]),
    .o(\cu_ru/m_s_tval/n11 [48]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6485 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [47]),
    .d(data_csr[47]),
    .o(_al_u6485_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6486 (
    .a(_al_u6485_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [47]),
    .o(\cu_ru/m_s_tval/n11 [47]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6487 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [46]),
    .d(data_csr[46]),
    .o(_al_u6487_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6488 (
    .a(_al_u6487_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [46]),
    .o(\cu_ru/m_s_tval/n11 [46]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6489 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [45]),
    .d(data_csr[45]),
    .o(_al_u6489_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6490 (
    .a(_al_u6489_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [45]),
    .o(\cu_ru/m_s_tval/n11 [45]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6491 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [44]),
    .d(data_csr[44]),
    .o(_al_u6491_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6492 (
    .a(_al_u6491_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [44]),
    .o(\cu_ru/m_s_tval/n11 [44]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6493 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [43]),
    .d(data_csr[43]),
    .o(_al_u6493_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6494 (
    .a(_al_u6493_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [43]),
    .o(\cu_ru/m_s_tval/n11 [43]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6495 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [42]),
    .d(data_csr[42]),
    .o(_al_u6495_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6496 (
    .a(_al_u6495_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [42]),
    .o(\cu_ru/m_s_tval/n11 [42]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6497 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [41]),
    .d(data_csr[41]),
    .o(_al_u6497_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6498 (
    .a(_al_u6497_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [41]),
    .o(\cu_ru/m_s_tval/n11 [41]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6499 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [40]),
    .d(data_csr[40]),
    .o(_al_u6499_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6500 (
    .a(_al_u6499_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [40]),
    .o(\cu_ru/m_s_tval/n11 [40]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6501 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [3]),
    .d(data_csr[3]),
    .o(_al_u6501_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6502 (
    .a(_al_u6501_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [3]),
    .o(\cu_ru/m_s_tval/n11 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6503 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [39]),
    .d(data_csr[39]),
    .o(_al_u6503_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6504 (
    .a(_al_u6503_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [39]),
    .o(\cu_ru/m_s_tval/n11 [39]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6505 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [38]),
    .d(data_csr[38]),
    .o(_al_u6505_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6506 (
    .a(_al_u6505_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [38]),
    .o(\cu_ru/m_s_tval/n11 [38]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6507 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [37]),
    .d(data_csr[37]),
    .o(_al_u6507_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6508 (
    .a(_al_u6507_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [37]),
    .o(\cu_ru/m_s_tval/n11 [37]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6509 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [36]),
    .d(data_csr[36]),
    .o(_al_u6509_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6510 (
    .a(_al_u6509_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [36]),
    .o(\cu_ru/m_s_tval/n11 [36]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6511 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [35]),
    .d(data_csr[35]),
    .o(_al_u6511_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6512 (
    .a(_al_u6511_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [35]),
    .o(\cu_ru/m_s_tval/n11 [35]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6513 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [34]),
    .d(data_csr[34]),
    .o(_al_u6513_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6514 (
    .a(_al_u6513_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [34]),
    .o(\cu_ru/m_s_tval/n11 [34]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6515 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [33]),
    .d(data_csr[33]),
    .o(_al_u6515_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6516 (
    .a(_al_u6515_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [33]),
    .o(\cu_ru/m_s_tval/n11 [33]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6517 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [32]),
    .d(data_csr[32]),
    .o(_al_u6517_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6518 (
    .a(_al_u6517_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [32]),
    .o(\cu_ru/m_s_tval/n11 [32]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6519 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [31]),
    .d(data_csr[31]),
    .o(_al_u6519_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6520 (
    .a(_al_u6519_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [31]),
    .o(\cu_ru/m_s_tval/n11 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6521 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [30]),
    .d(data_csr[30]),
    .o(_al_u6521_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6522 (
    .a(_al_u6521_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [30]),
    .o(\cu_ru/m_s_tval/n11 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6523 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [2]),
    .d(data_csr[2]),
    .o(_al_u6523_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6524 (
    .a(_al_u6523_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [2]),
    .o(\cu_ru/m_s_tval/n11 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6525 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [29]),
    .d(data_csr[29]),
    .o(_al_u6525_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6526 (
    .a(_al_u6525_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [29]),
    .o(\cu_ru/m_s_tval/n11 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6527 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [28]),
    .d(data_csr[28]),
    .o(_al_u6527_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6528 (
    .a(_al_u6527_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [28]),
    .o(\cu_ru/m_s_tval/n11 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6529 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [27]),
    .d(data_csr[27]),
    .o(_al_u6529_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6530 (
    .a(_al_u6529_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [27]),
    .o(\cu_ru/m_s_tval/n11 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6531 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [26]),
    .d(data_csr[26]),
    .o(_al_u6531_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6532 (
    .a(_al_u6531_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [26]),
    .o(\cu_ru/m_s_tval/n11 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6533 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [25]),
    .d(data_csr[25]),
    .o(_al_u6533_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6534 (
    .a(_al_u6533_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [25]),
    .o(\cu_ru/m_s_tval/n11 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6535 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [24]),
    .d(data_csr[24]),
    .o(_al_u6535_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6536 (
    .a(_al_u6535_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [24]),
    .o(\cu_ru/m_s_tval/n11 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6537 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [23]),
    .d(data_csr[23]),
    .o(_al_u6537_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6538 (
    .a(_al_u6537_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [23]),
    .o(\cu_ru/m_s_tval/n11 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6539 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [22]),
    .d(data_csr[22]),
    .o(_al_u6539_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6540 (
    .a(_al_u6539_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [22]),
    .o(\cu_ru/m_s_tval/n11 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6541 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [21]),
    .d(data_csr[21]),
    .o(_al_u6541_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6542 (
    .a(_al_u6541_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [21]),
    .o(\cu_ru/m_s_tval/n11 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6543 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [20]),
    .d(data_csr[20]),
    .o(_al_u6543_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6544 (
    .a(_al_u6543_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [20]),
    .o(\cu_ru/m_s_tval/n11 [20]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6545 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [1]),
    .d(data_csr[1]),
    .o(_al_u6545_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6546 (
    .a(_al_u6545_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [1]),
    .o(\cu_ru/m_s_tval/n11 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6547 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [19]),
    .d(data_csr[19]),
    .o(_al_u6547_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6548 (
    .a(_al_u6547_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [19]),
    .o(\cu_ru/m_s_tval/n11 [19]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6549 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [18]),
    .d(data_csr[18]),
    .o(_al_u6549_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6550 (
    .a(_al_u6549_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [18]),
    .o(\cu_ru/m_s_tval/n11 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6551 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [17]),
    .d(data_csr[17]),
    .o(_al_u6551_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6552 (
    .a(_al_u6551_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [17]),
    .o(\cu_ru/m_s_tval/n11 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6553 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [16]),
    .d(data_csr[16]),
    .o(_al_u6553_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6554 (
    .a(_al_u6553_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [16]),
    .o(\cu_ru/m_s_tval/n11 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6555 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [15]),
    .d(data_csr[15]),
    .o(_al_u6555_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6556 (
    .a(_al_u6555_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [15]),
    .o(\cu_ru/m_s_tval/n11 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6557 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [14]),
    .d(data_csr[14]),
    .o(_al_u6557_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6558 (
    .a(_al_u6557_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [14]),
    .o(\cu_ru/m_s_tval/n11 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6559 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [13]),
    .d(data_csr[13]),
    .o(_al_u6559_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6560 (
    .a(_al_u6559_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [13]),
    .o(\cu_ru/m_s_tval/n11 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6561 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [12]),
    .d(data_csr[12]),
    .o(_al_u6561_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6562 (
    .a(_al_u6561_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [12]),
    .o(\cu_ru/m_s_tval/n11 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6563 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [11]),
    .d(data_csr[11]),
    .o(_al_u6563_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6564 (
    .a(_al_u6563_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [11]),
    .o(\cu_ru/m_s_tval/n11 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6565 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [10]),
    .d(data_csr[10]),
    .o(_al_u6565_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6566 (
    .a(_al_u6565_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [10]),
    .o(\cu_ru/m_s_tval/n11 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6567 (
    .a(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mtval [0]),
    .d(data_csr[0]),
    .o(_al_u6567_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6568 (
    .a(_al_u6567_o),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/m_s_tval/n3 [0]),
    .o(\cu_ru/m_s_tval/n11 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u6569 (
    .a(_al_u5992_o),
    .b(_al_u3200_o),
    .c(csr_index[1]),
    .d(csr_index[2]),
    .o(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6570 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [9]),
    .d(data_csr[9]),
    .o(_al_u6570_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6571 (
    .a(_al_u6570_o),
    .b(\cu_ru/m_s_epc/n2 [9]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6572 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [8]),
    .d(data_csr[8]),
    .o(_al_u6572_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6573 (
    .a(_al_u6572_o),
    .b(\cu_ru/m_s_epc/n2 [8]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6574 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [7]),
    .d(data_csr[7]),
    .o(_al_u6574_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6575 (
    .a(_al_u6574_o),
    .b(\cu_ru/m_s_epc/n2 [7]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6576 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [6]),
    .d(data_csr[6]),
    .o(_al_u6576_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6577 (
    .a(_al_u6576_o),
    .b(\cu_ru/m_s_epc/n2 [6]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6578 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [63]),
    .d(data_csr[63]),
    .o(_al_u6578_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6579 (
    .a(_al_u6578_o),
    .b(\cu_ru/m_s_epc/n2 [63]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [63]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6580 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [62]),
    .d(data_csr[62]),
    .o(_al_u6580_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6581 (
    .a(_al_u6580_o),
    .b(\cu_ru/m_s_epc/n2 [62]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [62]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6582 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [61]),
    .d(data_csr[61]),
    .o(_al_u6582_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6583 (
    .a(_al_u6582_o),
    .b(\cu_ru/m_s_epc/n2 [61]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [61]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6584 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [60]),
    .d(data_csr[60]),
    .o(_al_u6584_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6585 (
    .a(_al_u6584_o),
    .b(\cu_ru/m_s_epc/n2 [60]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [60]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6586 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [5]),
    .d(data_csr[5]),
    .o(_al_u6586_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6587 (
    .a(_al_u6586_o),
    .b(\cu_ru/m_s_epc/n2 [5]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6588 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [59]),
    .d(data_csr[59]),
    .o(_al_u6588_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6589 (
    .a(_al_u6588_o),
    .b(\cu_ru/m_s_epc/n2 [59]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [59]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6590 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [58]),
    .d(data_csr[58]),
    .o(_al_u6590_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6591 (
    .a(_al_u6590_o),
    .b(\cu_ru/m_s_epc/n2 [58]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [58]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6592 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [57]),
    .d(data_csr[57]),
    .o(_al_u6592_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6593 (
    .a(_al_u6592_o),
    .b(\cu_ru/m_s_epc/n2 [57]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [57]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6594 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [56]),
    .d(data_csr[56]),
    .o(_al_u6594_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6595 (
    .a(_al_u6594_o),
    .b(\cu_ru/m_s_epc/n2 [56]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [56]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6596 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [55]),
    .d(data_csr[55]),
    .o(_al_u6596_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6597 (
    .a(_al_u6596_o),
    .b(\cu_ru/m_s_epc/n2 [55]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [55]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6598 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [54]),
    .d(data_csr[54]),
    .o(_al_u6598_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6599 (
    .a(_al_u6598_o),
    .b(\cu_ru/m_s_epc/n2 [54]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [54]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6600 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [53]),
    .d(data_csr[53]),
    .o(_al_u6600_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6601 (
    .a(_al_u6600_o),
    .b(\cu_ru/m_s_epc/n2 [53]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [53]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6602 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [52]),
    .d(data_csr[52]),
    .o(_al_u6602_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6603 (
    .a(_al_u6602_o),
    .b(\cu_ru/m_s_epc/n2 [52]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [52]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6604 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [51]),
    .d(data_csr[51]),
    .o(_al_u6604_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6605 (
    .a(_al_u6604_o),
    .b(\cu_ru/m_s_epc/n2 [51]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [51]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6606 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [50]),
    .d(data_csr[50]),
    .o(_al_u6606_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6607 (
    .a(_al_u6606_o),
    .b(\cu_ru/m_s_epc/n2 [50]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [50]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6608 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [4]),
    .d(data_csr[4]),
    .o(_al_u6608_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6609 (
    .a(_al_u6608_o),
    .b(\cu_ru/m_s_epc/n2 [4]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6610 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [49]),
    .d(data_csr[49]),
    .o(_al_u6610_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6611 (
    .a(_al_u6610_o),
    .b(\cu_ru/m_s_epc/n2 [49]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [49]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6612 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [48]),
    .d(data_csr[48]),
    .o(_al_u6612_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6613 (
    .a(_al_u6612_o),
    .b(\cu_ru/m_s_epc/n2 [48]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [48]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6614 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [47]),
    .d(data_csr[47]),
    .o(_al_u6614_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6615 (
    .a(_al_u6614_o),
    .b(\cu_ru/m_s_epc/n2 [47]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [47]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6616 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [46]),
    .d(data_csr[46]),
    .o(_al_u6616_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6617 (
    .a(_al_u6616_o),
    .b(\cu_ru/m_s_epc/n2 [46]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [46]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6618 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [45]),
    .d(data_csr[45]),
    .o(_al_u6618_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6619 (
    .a(_al_u6618_o),
    .b(\cu_ru/m_s_epc/n2 [45]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [45]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6620 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [44]),
    .d(data_csr[44]),
    .o(_al_u6620_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6621 (
    .a(_al_u6620_o),
    .b(\cu_ru/m_s_epc/n2 [44]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [44]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6622 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [43]),
    .d(data_csr[43]),
    .o(_al_u6622_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6623 (
    .a(_al_u6622_o),
    .b(\cu_ru/m_s_epc/n2 [43]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [43]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6624 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [42]),
    .d(data_csr[42]),
    .o(_al_u6624_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6625 (
    .a(_al_u6624_o),
    .b(\cu_ru/m_s_epc/n2 [42]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [42]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6626 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [41]),
    .d(data_csr[41]),
    .o(_al_u6626_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6627 (
    .a(_al_u6626_o),
    .b(\cu_ru/m_s_epc/n2 [41]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [41]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6628 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [40]),
    .d(data_csr[40]),
    .o(_al_u6628_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6629 (
    .a(_al_u6628_o),
    .b(\cu_ru/m_s_epc/n2 [40]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [40]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6630 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [3]),
    .d(data_csr[3]),
    .o(_al_u6630_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6631 (
    .a(_al_u6630_o),
    .b(\cu_ru/m_s_epc/n2 [3]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6632 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [39]),
    .d(data_csr[39]),
    .o(_al_u6632_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6633 (
    .a(_al_u6632_o),
    .b(\cu_ru/m_s_epc/n2 [39]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [39]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6634 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [38]),
    .d(data_csr[38]),
    .o(_al_u6634_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6635 (
    .a(_al_u6634_o),
    .b(\cu_ru/m_s_epc/n2 [38]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [38]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6636 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [37]),
    .d(data_csr[37]),
    .o(_al_u6636_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6637 (
    .a(_al_u6636_o),
    .b(\cu_ru/m_s_epc/n2 [37]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [37]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6638 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [36]),
    .d(data_csr[36]),
    .o(_al_u6638_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6639 (
    .a(_al_u6638_o),
    .b(\cu_ru/m_s_epc/n2 [36]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [36]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6640 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [35]),
    .d(data_csr[35]),
    .o(_al_u6640_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6641 (
    .a(_al_u6640_o),
    .b(\cu_ru/m_s_epc/n2 [35]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [35]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6642 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [34]),
    .d(data_csr[34]),
    .o(_al_u6642_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6643 (
    .a(_al_u6642_o),
    .b(\cu_ru/m_s_epc/n2 [34]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [34]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6644 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [33]),
    .d(data_csr[33]),
    .o(_al_u6644_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6645 (
    .a(_al_u6644_o),
    .b(\cu_ru/m_s_epc/n2 [33]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [33]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6646 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [32]),
    .d(data_csr[32]),
    .o(_al_u6646_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6647 (
    .a(_al_u6646_o),
    .b(\cu_ru/m_s_epc/n2 [32]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [32]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6648 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [31]),
    .d(data_csr[31]),
    .o(_al_u6648_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6649 (
    .a(_al_u6648_o),
    .b(\cu_ru/m_s_epc/n2 [31]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6650 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [30]),
    .d(data_csr[30]),
    .o(_al_u6650_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6651 (
    .a(_al_u6650_o),
    .b(\cu_ru/m_s_epc/n2 [30]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6652 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [2]),
    .d(data_csr[2]),
    .o(_al_u6652_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6653 (
    .a(_al_u6652_o),
    .b(\cu_ru/m_s_epc/n2 [2]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6654 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [29]),
    .d(data_csr[29]),
    .o(_al_u6654_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6655 (
    .a(_al_u6654_o),
    .b(\cu_ru/m_s_epc/n2 [29]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6656 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [28]),
    .d(data_csr[28]),
    .o(_al_u6656_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6657 (
    .a(_al_u6656_o),
    .b(\cu_ru/m_s_epc/n2 [28]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6658 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [27]),
    .d(data_csr[27]),
    .o(_al_u6658_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6659 (
    .a(_al_u6658_o),
    .b(\cu_ru/m_s_epc/n2 [27]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6660 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [26]),
    .d(data_csr[26]),
    .o(_al_u6660_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6661 (
    .a(_al_u6660_o),
    .b(\cu_ru/m_s_epc/n2 [26]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6662 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [25]),
    .d(data_csr[25]),
    .o(_al_u6662_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6663 (
    .a(_al_u6662_o),
    .b(\cu_ru/m_s_epc/n2 [25]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6664 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [24]),
    .d(data_csr[24]),
    .o(_al_u6664_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6665 (
    .a(_al_u6664_o),
    .b(\cu_ru/m_s_epc/n2 [24]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6666 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [23]),
    .d(data_csr[23]),
    .o(_al_u6666_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6667 (
    .a(_al_u6666_o),
    .b(\cu_ru/m_s_epc/n2 [23]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6668 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [22]),
    .d(data_csr[22]),
    .o(_al_u6668_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6669 (
    .a(_al_u6668_o),
    .b(\cu_ru/m_s_epc/n2 [22]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6670 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [21]),
    .d(data_csr[21]),
    .o(_al_u6670_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6671 (
    .a(_al_u6670_o),
    .b(\cu_ru/m_s_epc/n2 [21]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6672 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [20]),
    .d(data_csr[20]),
    .o(_al_u6672_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6673 (
    .a(_al_u6672_o),
    .b(\cu_ru/m_s_epc/n2 [20]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [20]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6674 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [1]),
    .d(data_csr[1]),
    .o(_al_u6674_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6675 (
    .a(_al_u6674_o),
    .b(\cu_ru/m_s_epc/n2 [1]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6676 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [19]),
    .d(data_csr[19]),
    .o(_al_u6676_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6677 (
    .a(_al_u6676_o),
    .b(\cu_ru/m_s_epc/n2 [19]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [19]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6678 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [18]),
    .d(data_csr[18]),
    .o(_al_u6678_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6679 (
    .a(_al_u6678_o),
    .b(\cu_ru/m_s_epc/n2 [18]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6680 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [17]),
    .d(data_csr[17]),
    .o(_al_u6680_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6681 (
    .a(_al_u6680_o),
    .b(\cu_ru/m_s_epc/n2 [17]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6682 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [16]),
    .d(data_csr[16]),
    .o(_al_u6682_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6683 (
    .a(_al_u6682_o),
    .b(\cu_ru/m_s_epc/n2 [16]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6684 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [15]),
    .d(data_csr[15]),
    .o(_al_u6684_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6685 (
    .a(_al_u6684_o),
    .b(\cu_ru/m_s_epc/n2 [15]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6686 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [14]),
    .d(data_csr[14]),
    .o(_al_u6686_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6687 (
    .a(_al_u6686_o),
    .b(\cu_ru/m_s_epc/n2 [14]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6688 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [13]),
    .d(data_csr[13]),
    .o(_al_u6688_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6689 (
    .a(_al_u6688_o),
    .b(\cu_ru/m_s_epc/n2 [13]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6690 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [12]),
    .d(data_csr[12]),
    .o(_al_u6690_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6691 (
    .a(_al_u6690_o),
    .b(\cu_ru/m_s_epc/n2 [12]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6692 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [11]),
    .d(data_csr[11]),
    .o(_al_u6692_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6693 (
    .a(_al_u6692_o),
    .b(\cu_ru/m_s_epc/n2 [11]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6694 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mepc [10]),
    .d(data_csr[10]),
    .o(_al_u6694_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u6695 (
    .a(_al_u6694_o),
    .b(\cu_ru/m_s_epc/n2 [10]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [10]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u6696 (
    .a(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .b(\cu_ru/mepc [0]),
    .c(data_csr[0]),
    .o(_al_u6696_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u6697 (
    .a(_al_u6696_o),
    .b(\cu_ru/m_s_epc/n2 [0]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6698 (
    .a(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mcause [63]),
    .d(data_csr[63]),
    .o(_al_u6698_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u6699 (
    .a(_al_u6698_o),
    .b(\cu_ru/trap_target_m ),
    .c(_al_u4234_o),
    .o(\cu_ru/m_s_cause/n7 [63]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u6700 (
    .a(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/mcause [2]),
    .c(data_csr[2]),
    .o(_al_u6700_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u6701 (
    .a(_al_u6700_o),
    .b(\cu_ru/trap_cause [2]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_cause/n7 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u6702 (
    .a(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/mcause [0]),
    .d(data_csr[0]),
    .o(_al_u6702_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u6703 (
    .a(\cu_ru/trap_cause [0]),
    .b(_al_u6702_o),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_cause/n7 [0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6704 (
    .a(\biu/cache_ctrl_logic/ex_l1i_hit ),
    .b(_al_u6425_o),
    .o(_al_u6704_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u6705 (
    .a(_al_u6321_o),
    .b(_al_u6704_o),
    .o(\biu/ex_data_sel [0]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u6706 (
    .a(\biu/ex_data_sel [0]),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(addr_ex[11]),
    .d(addr_if[11]),
    .o(_al_u6706_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    _al_u6707 (
    .a(_al_u6706_o),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(_al_u2891_o),
    .o(\biu/l1i_addr [8]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u6708 (
    .a(\biu/ex_data_sel [0]),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(addr_ex[10]),
    .d(addr_if[10]),
    .o(_al_u6708_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    _al_u6709 (
    .a(_al_u6708_o),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(_al_u2893_o),
    .o(\biu/l1i_addr [7]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u6710 (
    .a(\biu/ex_data_sel [0]),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(addr_ex[9]),
    .d(addr_if[9]),
    .o(_al_u6710_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    _al_u6711 (
    .a(_al_u6710_o),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(_al_u2895_o),
    .o(\biu/l1i_addr [6]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6712 (
    .a(\biu/ex_data_sel [0]),
    .b(addr_ex[8]),
    .c(addr_if[8]),
    .o(_al_u6712_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u6713 (
    .a(_al_u6712_o),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(_al_u2897_o),
    .o(\biu/l1i_addr [5]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6714 (
    .a(\biu/ex_data_sel [0]),
    .b(addr_ex[7]),
    .c(addr_if[7]),
    .o(_al_u6714_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u6715 (
    .a(_al_u6714_o),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(_al_u2899_o),
    .o(\biu/l1i_addr [4]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6716 (
    .a(\biu/ex_data_sel [0]),
    .b(addr_ex[6]),
    .c(addr_if[6]),
    .o(_al_u6716_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u6717 (
    .a(_al_u6716_o),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(_al_u2901_o),
    .o(\biu/l1i_addr [3]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6718 (
    .a(\biu/ex_data_sel [0]),
    .b(addr_ex[5]),
    .c(addr_if[5]),
    .o(_al_u6718_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u6719 (
    .a(_al_u6718_o),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(_al_u2903_o),
    .o(\biu/l1i_addr [2]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6720 (
    .a(\biu/ex_data_sel [0]),
    .b(addr_ex[4]),
    .c(addr_if[4]),
    .o(_al_u6720_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u6721 (
    .a(_al_u6720_o),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(_al_u2905_o),
    .o(\biu/l1i_addr [1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u6722 (
    .a(\biu/ex_data_sel [0]),
    .b(addr_ex[3]),
    .c(addr_if[3]),
    .o(_al_u6722_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u6723 (
    .a(_al_u6722_o),
    .b(\biu/bus_unit/mux1_b1_sel_is_0_o ),
    .c(_al_u2907_o),
    .o(\biu/l1i_addr [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u6724 (
    .a(_al_u6309_o),
    .b(_al_u6320_o),
    .c(\biu/cache_ctrl_logic/ex_l1i_hit ),
    .d(_al_u6425_o),
    .o(_al_u6724_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6725 (
    .a(_al_u2835_o),
    .b(_al_u2837_o),
    .o(_al_u6725_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u6726 (
    .a(_al_u6724_o),
    .b(_al_u6725_o),
    .o(load_page_fault));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u6727 (
    .a(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/mcause [3]),
    .c(data_csr[3]),
    .o(_al_u6727_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u6728 (
    .a(_al_u6727_o),
    .b(\cu_ru/trap_cause [3]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_cause/n7 [3]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u6729 (
    .a(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .b(\cu_ru/scause [3]),
    .c(data_csr[3]),
    .o(_al_u6729_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u6730 (
    .a(\cu_ru/trap_cause [3]),
    .b(_al_u5157_o),
    .c(_al_u6729_o),
    .o(\cu_ru/m_s_cause/n5 [3]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6731 (
    .a(\cu_ru/trap_target_m ),
    .b(_al_u2844_o),
    .c(\cu_ru/mtvec [3]),
    .o(_al_u6731_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6732 (
    .a(_al_u6055_o),
    .b(_al_u6731_o),
    .c(new_pc[1]),
    .o(_al_u6732_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6733 (
    .a(_al_u6732_o),
    .b(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .c(\cu_ru/stvec [3]),
    .o(_al_u6733_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6734 (
    .a(_al_u2844_o),
    .b(\cu_ru/sepc [1]),
    .o(_al_u6734_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u6735 (
    .a(_al_u6733_o),
    .b(_al_u6734_o),
    .c(\cu_ru/m_s_status/n2 ),
    .d(\cu_ru/mepc [1]),
    .o(flush_pc[1]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u6736 (
    .a(\cu_ru/trap_target_m ),
    .b(_al_u2844_o),
    .c(\cu_ru/mtvec [2]),
    .o(_al_u6736_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u6737 (
    .a(_al_u6055_o),
    .b(_al_u6736_o),
    .c(new_pc[0]),
    .o(_al_u6737_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6738 (
    .a(_al_u6737_o),
    .b(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .c(\cu_ru/stvec [2]),
    .o(_al_u6738_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6739 (
    .a(_al_u2844_o),
    .b(\cu_ru/sepc [0]),
    .o(_al_u6739_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u6740 (
    .a(_al_u6738_o),
    .b(_al_u6739_o),
    .c(\cu_ru/m_s_status/n2 ),
    .d(\cu_ru/mepc [0]),
    .o(flush_pc[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6741 (
    .a(\cu_ru/trap_target_m ),
    .b(wb_s_ret),
    .o(\cu_ru/m_s_status/mux3_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6742 (
    .a(_al_u3427_o),
    .b(\cu_ru/m_s_status/n2 ),
    .c(\cu_ru/mstatus [7]),
    .o(_al_u6742_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u6743 (
    .a(\cu_ru/m_s_status/mux3_b0_sel_is_2_o ),
    .b(_al_u6742_o),
    .c(\cu_ru/m_s_status/n2 ),
    .d(\cu_ru/mie ),
    .o(_al_u6743_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6744 (
    .a(_al_u3427_o),
    .b(\cu_ru/mie ),
    .o(_al_u6744_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u6745 (
    .a(_al_u6743_o),
    .b(_al_u6744_o),
    .c(\cu_ru/m_s_status/n0 ),
    .d(data_csr[3]),
    .o(\cu_ru/m_s_status/n37 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6746 (
    .a(_al_u3427_o),
    .b(\cu_ru/m_s_status/n2 ),
    .o(_al_u6746_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u6747 (
    .a(\cu_ru/m_s_status/mux3_b0_sel_is_2_o ),
    .b(_al_u6746_o),
    .c(\cu_ru/mie ),
    .d(\cu_ru/mstatus [7]),
    .o(_al_u6747_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6748 (
    .a(_al_u3427_o),
    .b(\cu_ru/mstatus [7]),
    .o(_al_u6748_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6749 (
    .a(_al_u6747_o),
    .b(_al_u6748_o),
    .c(\cu_ru/m_s_status/n0 ),
    .d(data_csr[7]),
    .o(\cu_ru/m_s_status/n45 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6750 (
    .a(\cu_ru/m_s_status/n5 [1]),
    .b(priv[3]),
    .o(_al_u6750_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))"),
    .INIT(16'h4c08))
    _al_u6751 (
    .a(\cu_ru/m_s_status/mux3_b0_sel_is_2_o ),
    .b(_al_u6746_o),
    .c(_al_u6750_o),
    .d(\cu_ru/mstatus [12]),
    .o(_al_u6751_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6752 (
    .a(_al_u3427_o),
    .b(\cu_ru/mstatus [12]),
    .o(_al_u6752_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6753 (
    .a(_al_u6751_o),
    .b(_al_u6752_o),
    .c(\cu_ru/m_s_status/n0 ),
    .d(data_csr[12]),
    .o(\cu_ru/m_s_status/n47 [1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))"),
    .INIT(16'h4c08))
    _al_u6754 (
    .a(\cu_ru/m_s_status/mux3_b0_sel_is_2_o ),
    .b(_al_u6746_o),
    .c(_al_u6313_o),
    .d(\cu_ru/mstatus [11]),
    .o(_al_u6754_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6755 (
    .a(_al_u3427_o),
    .b(\cu_ru/mstatus [11]),
    .o(_al_u6755_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u6756 (
    .a(_al_u6754_o),
    .b(_al_u6755_o),
    .c(\cu_ru/m_s_status/n0 ),
    .d(data_csr[11]),
    .o(\cu_ru/m_s_status/n47 [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u6757 (
    .a(_al_u3400_o),
    .b(id_ins[31]),
    .c(id_ins[30]),
    .d(id_ins[29]),
    .o(_al_u6757_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u6758 (
    .a(_al_u3393_o),
    .b(id_ins[22]),
    .c(id_ins[21]),
    .d(id_ins[20]),
    .o(_al_u6758_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6759 (
    .a(_al_u6757_o),
    .b(_al_u6758_o),
    .o(\cu_ru/read_minstret_sel_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6760 (
    .a(id_ins[31]),
    .b(id_ins[30]),
    .o(_al_u6760_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6761 (
    .a(\ins_dec/n80_lutinv ),
    .b(_al_u6760_o),
    .c(_al_u3387_o),
    .o(_al_u6761_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6762 (
    .a(_al_u6761_o),
    .b(_al_u6758_o),
    .o(\cu_ru/read_instret_sel_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6763 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_instret_sel_lutinv ),
    .o(_al_u6763_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u6764 (
    .a(_al_u3393_o),
    .b(id_ins[22]),
    .c(id_ins[21]),
    .d(id_ins[20]),
    .o(_al_u6764_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u6765 (
    .a(id_ins[28]),
    .b(id_ins[27]),
    .c(id_ins[26]),
    .o(_al_u6765_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6766 (
    .a(_al_u6765_o),
    .b(id_ins[29]),
    .c(_al_u3388_o),
    .o(_al_u6766_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6767 (
    .a(_al_u6764_o),
    .b(_al_u6766_o),
    .o(\cu_ru/read_mtval_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6768 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/minstret [59]),
    .d(\cu_ru/mtval [59]),
    .o(_al_u6768_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6769 (
    .a(_al_u3399_o),
    .b(_al_u6765_o),
    .o(_al_u6769_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6770 (
    .a(_al_u6769_o),
    .b(_al_u3397_o),
    .o(\cu_ru/read_sscratch_sel_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6771 (
    .a(_al_u6758_o),
    .b(_al_u6766_o),
    .o(\cu_ru/read_mcause_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6772 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [59]),
    .d(\cu_ru/sscratch [59]),
    .o(_al_u6772_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6773 (
    .a(_al_u6769_o),
    .b(_al_u6758_o),
    .o(\cu_ru/read_scause_sel_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6774 (
    .a(_al_u6766_o),
    .b(_al_u3397_o),
    .o(\cu_ru/read_mscratch_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6775 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [59]),
    .d(\cu_ru/mscratch [59]),
    .o(_al_u6775_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6776 (
    .a(_al_u3395_o),
    .b(_al_u6766_o),
    .o(\cu_ru/read_mepc_sel_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6777 (
    .a(_al_u3399_o),
    .b(_al_u3400_o),
    .o(_al_u6777_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u6778 (
    .a(_al_u3393_o),
    .b(id_ins[22]),
    .c(id_ins[21]),
    .d(id_ins[20]),
    .o(_al_u6778_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6779 (
    .a(_al_u6777_o),
    .b(_al_u6778_o),
    .o(\cu_ru/read_stvec_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6780 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [59]),
    .d(\cu_ru/stvec [59]),
    .o(_al_u6780_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6781 (
    .a(_al_u6772_o),
    .b(_al_u6775_o),
    .c(_al_u6780_o),
    .o(_al_u6781_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6782 (
    .a(_al_u3395_o),
    .b(_al_u6761_o),
    .o(\cu_ru/read_time_sel_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6783 (
    .a(_al_u3395_o),
    .b(_al_u6769_o),
    .o(\cu_ru/read_sepc_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6784 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(mtime_pad[59]),
    .d(\cu_ru/sepc [59]),
    .o(_al_u6784_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6785 (
    .a(_al_u6768_o),
    .b(_al_u6781_o),
    .c(_al_u6784_o),
    .o(_al_u6785_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6786 (
    .a(_al_u6757_o),
    .b(_al_u3397_o),
    .o(\cu_ru/read_mcycle_sel_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6787 (
    .a(_al_u6761_o),
    .b(_al_u3397_o),
    .o(\cu_ru/read_cycle_sel_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u6788 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_cycle_sel_lutinv ),
    .o(_al_u6788_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6789 (
    .a(_al_u6764_o),
    .b(_al_u6769_o),
    .o(\cu_ru/read_stval_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6790 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/mcycle [59]),
    .d(\cu_ru/stval [59]),
    .o(_al_u6790_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u6791 (
    .a(id_ins[29]),
    .b(id_ins[28]),
    .c(_al_u3387_o),
    .d(_al_u3388_o),
    .o(_al_u6791_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6792 (
    .a(_al_u6778_o),
    .b(_al_u6791_o),
    .o(\cu_ru/read_mtvec_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u6793 (
    .a(_al_u6785_o),
    .b(_al_u6790_o),
    .c(\cu_ru/read_mtvec_sel_lutinv ),
    .d(\cu_ru/mtvec [59]),
    .o(csr_data[59]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6794 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [58]),
    .d(\cu_ru/stval [58]),
    .o(_al_u6794_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6795 (
    .a(_al_u6763_o),
    .b(_al_u6794_o),
    .c(\cu_ru/minstret [58]),
    .o(_al_u6795_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6796 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [58]),
    .d(\cu_ru/stvec [58]),
    .o(_al_u6796_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6797 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [58]),
    .d(\cu_ru/mcause [58]),
    .o(_al_u6797_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6798 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mscratch [58]),
    .d(\cu_ru/sscratch [58]),
    .o(_al_u6798_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6799 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [58]),
    .d(\cu_ru/mtval [58]),
    .o(_al_u6799_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6800 (
    .a(_al_u6797_o),
    .b(_al_u6798_o),
    .c(_al_u6799_o),
    .o(_al_u6800_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6801 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[58]),
    .d(\cu_ru/mtvec [58]),
    .o(_al_u6801_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6802 (
    .a(_al_u6795_o),
    .b(_al_u6796_o),
    .c(_al_u6800_o),
    .d(_al_u6801_o),
    .o(csr_data[58]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6803 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [57]),
    .d(\cu_ru/stvec [57]),
    .o(_al_u6803_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6804 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [57]),
    .d(\cu_ru/sscratch [57]),
    .o(_al_u6804_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6805 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [57]),
    .d(\cu_ru/mscratch [57]),
    .o(_al_u6805_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6806 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [57]),
    .d(\cu_ru/mtval [57]),
    .o(_al_u6806_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6807 (
    .a(_al_u6804_o),
    .b(_al_u6805_o),
    .c(_al_u6806_o),
    .o(_al_u6807_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6808 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[57]),
    .d(\cu_ru/mtvec [57]),
    .o(_al_u6808_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6809 (
    .a(_al_u6803_o),
    .b(_al_u6807_o),
    .c(_al_u6808_o),
    .o(_al_u6809_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6810 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/minstret [57]),
    .d(\cu_ru/stval [57]),
    .o(_al_u6810_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u6811 (
    .a(_al_u6809_o),
    .b(_al_u6810_o),
    .c(\cu_ru/read_sepc_sel_lutinv ),
    .d(\cu_ru/sepc [57]),
    .o(csr_data[57]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6812 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/minstret [56]),
    .d(\cu_ru/stval [56]),
    .o(_al_u6812_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6813 (
    .a(_al_u6812_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [56]),
    .o(_al_u6813_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6814 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/mcycle [56]),
    .d(\cu_ru/scause [56]),
    .o(_al_u6814_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6815 (
    .a(_al_u6814_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mtval [56]),
    .o(_al_u6815_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6816 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcause [56]),
    .d(\cu_ru/mscratch [56]),
    .o(_al_u6816_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6817 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [56]),
    .d(\cu_ru/sscratch [56]),
    .o(_al_u6817_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6818 (
    .a(_al_u6815_o),
    .b(_al_u6816_o),
    .c(_al_u6817_o),
    .o(_al_u6818_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6819 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stvec [56]),
    .d(\cu_ru/mtvec [56]),
    .o(_al_u6819_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6820 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(mtime_pad[56]),
    .d(\cu_ru/mepc [56]),
    .o(_al_u6820_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6821 (
    .a(_al_u6813_o),
    .b(_al_u6818_o),
    .c(_al_u6819_o),
    .d(_al_u6820_o),
    .o(csr_data[56]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6822 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mcycle [55]),
    .d(\cu_ru/mtval [55]),
    .o(_al_u6822_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6823 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mscratch [55]),
    .d(\cu_ru/sscratch [55]),
    .o(_al_u6823_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6824 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [55]),
    .d(\cu_ru/mcause [55]),
    .o(_al_u6824_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6825 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [55]),
    .d(\cu_ru/stvec [55]),
    .o(_al_u6825_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6826 (
    .a(_al_u6823_o),
    .b(_al_u6824_o),
    .c(_al_u6825_o),
    .o(_al_u6826_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6827 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(mtime_pad[55]),
    .d(\cu_ru/sepc [55]),
    .o(_al_u6827_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6828 (
    .a(_al_u6822_o),
    .b(_al_u6826_o),
    .c(_al_u6827_o),
    .o(_al_u6828_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6829 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/minstret [55]),
    .d(\cu_ru/stval [55]),
    .o(_al_u6829_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u6830 (
    .a(_al_u6828_o),
    .b(_al_u6829_o),
    .c(\cu_ru/read_mtvec_sel_lutinv ),
    .d(\cu_ru/mtvec [55]),
    .o(csr_data[55]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6831 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/mcycle [54]),
    .d(\cu_ru/scause [54]),
    .o(_al_u6831_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6832 (
    .a(_al_u6831_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mtval [54]),
    .o(_al_u6832_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6833 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcause [54]),
    .d(\cu_ru/mscratch [54]),
    .o(_al_u6833_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6834 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [54]),
    .d(\cu_ru/sscratch [54]),
    .o(_al_u6834_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6835 (
    .a(_al_u6832_o),
    .b(_al_u6833_o),
    .c(_al_u6834_o),
    .o(_al_u6835_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6836 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[54]),
    .d(\cu_ru/stval [54]),
    .o(_al_u6836_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6837 (
    .a(_al_u6836_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [54]),
    .o(_al_u6837_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6838 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/minstret [54]),
    .d(\cu_ru/stvec [54]),
    .o(_al_u6838_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6839 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [54]),
    .d(\cu_ru/mtvec [54]),
    .o(_al_u6839_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6840 (
    .a(_al_u6835_o),
    .b(_al_u6837_o),
    .c(_al_u6838_o),
    .d(_al_u6839_o),
    .o(csr_data[54]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6841 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/minstret [53]),
    .d(\cu_ru/stvec [53]),
    .o(_al_u6841_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6842 (
    .a(_al_u6841_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [53]),
    .o(_al_u6842_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6843 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [53]),
    .d(\cu_ru/sscratch [53]),
    .o(_al_u6843_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u6844 (
    .a(_al_u6843_o),
    .b(\cu_ru/read_mcycle_sel_lutinv ),
    .c(\cu_ru/read_cycle_sel_lutinv ),
    .d(\cu_ru/mcycle [53]),
    .o(_al_u6844_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6845 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [53]),
    .d(\cu_ru/mscratch [53]),
    .o(_al_u6845_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6846 (
    .a(_al_u6844_o),
    .b(_al_u6845_o),
    .c(\cu_ru/read_mtvec_sel_lutinv ),
    .d(\cu_ru/mtvec [53]),
    .o(_al_u6846_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6847 (
    .a(\cu_ru/read_sepc_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/sepc [53]),
    .d(\cu_ru/mepc [53]),
    .o(_al_u6847_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6848 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[53]),
    .d(\cu_ru/mtval [53]),
    .o(_al_u6848_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6849 (
    .a(_al_u6842_o),
    .b(_al_u6846_o),
    .c(_al_u6847_o),
    .d(_al_u6848_o),
    .o(csr_data[53]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6850 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [52]),
    .d(\cu_ru/sscratch [52]),
    .o(_al_u6850_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6851 (
    .a(_al_u6850_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mtval [52]),
    .o(_al_u6851_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6852 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [52]),
    .d(\cu_ru/mscratch [52]),
    .o(_al_u6852_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6853 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcycle [52]),
    .d(\cu_ru/mcause [52]),
    .o(_al_u6853_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6854 (
    .a(_al_u6851_o),
    .b(_al_u6852_o),
    .c(_al_u6853_o),
    .o(_al_u6854_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6855 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(mtime_pad[52]),
    .d(\cu_ru/sepc [52]),
    .o(_al_u6855_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6856 (
    .a(_al_u6855_o),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [52]),
    .o(_al_u6856_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6857 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/minstret [52]),
    .d(\cu_ru/stvec [52]),
    .o(_al_u6857_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6858 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [52]),
    .d(\cu_ru/mtvec [52]),
    .o(_al_u6858_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6859 (
    .a(_al_u6854_o),
    .b(_al_u6856_o),
    .c(_al_u6857_o),
    .d(_al_u6858_o),
    .o(csr_data[52]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6860 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [51]),
    .d(\cu_ru/sscratch [51]),
    .o(_al_u6860_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6861 (
    .a(_al_u6860_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mtval [51]),
    .o(_al_u6861_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6862 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [51]),
    .d(\cu_ru/mscratch [51]),
    .o(_al_u6862_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6863 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcycle [51]),
    .d(\cu_ru/mcause [51]),
    .o(_al_u6863_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6864 (
    .a(_al_u6861_o),
    .b(_al_u6862_o),
    .c(_al_u6863_o),
    .o(_al_u6864_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6865 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(mtime_pad[51]),
    .d(\cu_ru/sepc [51]),
    .o(_al_u6865_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6866 (
    .a(_al_u6865_o),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [51]),
    .o(_al_u6866_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6867 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/minstret [51]),
    .d(\cu_ru/stvec [51]),
    .o(_al_u6867_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6868 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [51]),
    .d(\cu_ru/mtvec [51]),
    .o(_al_u6868_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6869 (
    .a(_al_u6864_o),
    .b(_al_u6866_o),
    .c(_al_u6867_o),
    .d(_al_u6868_o),
    .o(csr_data[51]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6870 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/minstret [50]),
    .d(\cu_ru/stval [50]),
    .o(_al_u6870_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6871 (
    .a(_al_u6870_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[50]),
    .o(_al_u6871_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6872 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [50]),
    .d(\cu_ru/mscratch [50]),
    .o(_al_u6872_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6873 (
    .a(_al_u6872_o),
    .b(\cu_ru/read_mtvec_sel_lutinv ),
    .c(\cu_ru/mtvec [50]),
    .o(_al_u6873_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6874 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcycle [50]),
    .d(\cu_ru/mcause [50]),
    .o(_al_u6874_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6875 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [50]),
    .d(\cu_ru/sscratch [50]),
    .o(_al_u6875_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6876 (
    .a(_al_u6873_o),
    .b(_al_u6874_o),
    .c(_al_u6875_o),
    .o(_al_u6876_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6877 (
    .a(\cu_ru/read_sepc_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/sepc [50]),
    .d(\cu_ru/mepc [50]),
    .o(_al_u6877_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6878 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mtval [50]),
    .d(\cu_ru/stvec [50]),
    .o(_al_u6878_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6879 (
    .a(_al_u6871_o),
    .b(_al_u6876_o),
    .c(_al_u6877_o),
    .d(_al_u6878_o),
    .o(csr_data[50]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6880 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/minstret [49]),
    .d(\cu_ru/sepc [49]),
    .o(_al_u6880_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6881 (
    .a(_al_u6880_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[49]),
    .o(_al_u6881_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6882 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [49]),
    .d(\cu_ru/mscratch [49]),
    .o(_al_u6882_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6883 (
    .a(_al_u6882_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [49]),
    .o(_al_u6883_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6884 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcycle [49]),
    .d(\cu_ru/mcause [49]),
    .o(_al_u6884_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6885 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [49]),
    .d(\cu_ru/sscratch [49]),
    .o(_al_u6885_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6886 (
    .a(_al_u6883_o),
    .b(_al_u6884_o),
    .c(_al_u6885_o),
    .o(_al_u6886_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6887 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [49]),
    .d(\cu_ru/stvec [49]),
    .o(_al_u6887_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6888 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mtval [49]),
    .d(\cu_ru/mtvec [49]),
    .o(_al_u6888_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6889 (
    .a(_al_u6881_o),
    .b(_al_u6886_o),
    .c(_al_u6887_o),
    .d(_al_u6888_o),
    .o(csr_data[49]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6890 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [48]),
    .d(\cu_ru/stvec [48]),
    .o(_al_u6890_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6891 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [48]),
    .d(\cu_ru/sscratch [48]),
    .o(_al_u6891_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6892 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [48]),
    .d(\cu_ru/mscratch [48]),
    .o(_al_u6892_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6893 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [48]),
    .d(\cu_ru/mtval [48]),
    .o(_al_u6893_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6894 (
    .a(_al_u6891_o),
    .b(_al_u6892_o),
    .c(_al_u6893_o),
    .o(_al_u6894_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6895 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(mtime_pad[48]),
    .d(\cu_ru/sepc [48]),
    .o(_al_u6895_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6896 (
    .a(_al_u6890_o),
    .b(_al_u6894_o),
    .c(_al_u6895_o),
    .o(_al_u6896_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6897 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/minstret [48]),
    .d(\cu_ru/stval [48]),
    .o(_al_u6897_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u6898 (
    .a(_al_u6896_o),
    .b(_al_u6897_o),
    .c(\cu_ru/read_mtvec_sel_lutinv ),
    .d(\cu_ru/mtvec [48]),
    .o(csr_data[48]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6899 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/minstret [47]),
    .d(\cu_ru/mtval [47]),
    .o(_al_u6899_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6900 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [47]),
    .d(\cu_ru/sscratch [47]),
    .o(_al_u6900_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6901 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [47]),
    .d(\cu_ru/mscratch [47]),
    .o(_al_u6901_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6902 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [47]),
    .d(\cu_ru/stvec [47]),
    .o(_al_u6902_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6903 (
    .a(_al_u6900_o),
    .b(_al_u6901_o),
    .c(_al_u6902_o),
    .o(_al_u6903_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6904 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[47]),
    .d(\cu_ru/mtvec [47]),
    .o(_al_u6904_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6905 (
    .a(_al_u6899_o),
    .b(_al_u6903_o),
    .c(_al_u6904_o),
    .o(_al_u6905_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6906 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/mcycle [47]),
    .d(\cu_ru/stval [47]),
    .o(_al_u6906_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u6907 (
    .a(_al_u6905_o),
    .b(_al_u6906_o),
    .c(\cu_ru/read_sepc_sel_lutinv ),
    .d(\cu_ru/sepc [47]),
    .o(csr_data[47]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6908 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [46]),
    .d(\cu_ru/stval [46]),
    .o(_al_u6908_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6909 (
    .a(_al_u6788_o),
    .b(_al_u6908_o),
    .c(\cu_ru/mcycle [46]),
    .o(_al_u6909_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6910 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/minstret [46]),
    .d(\cu_ru/stvec [46]),
    .o(_al_u6910_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6911 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [46]),
    .d(\cu_ru/mscratch [46]),
    .o(_al_u6911_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6912 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [46]),
    .d(\cu_ru/sscratch [46]),
    .o(_al_u6912_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6913 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [46]),
    .d(\cu_ru/mtval [46]),
    .o(_al_u6913_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6914 (
    .a(_al_u6911_o),
    .b(_al_u6912_o),
    .c(_al_u6913_o),
    .o(_al_u6914_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6915 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[46]),
    .d(\cu_ru/mtvec [46]),
    .o(_al_u6915_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6916 (
    .a(_al_u6909_o),
    .b(_al_u6910_o),
    .c(_al_u6914_o),
    .d(_al_u6915_o),
    .o(csr_data[46]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6917 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [45]),
    .d(\cu_ru/stval [45]),
    .o(_al_u6917_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6918 (
    .a(_al_u6788_o),
    .b(_al_u6917_o),
    .c(\cu_ru/mcycle [45]),
    .o(_al_u6918_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6919 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/minstret [45]),
    .d(\cu_ru/mtval [45]),
    .o(_al_u6919_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6920 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [45]),
    .d(\cu_ru/mcause [45]),
    .o(_al_u6920_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6921 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mscratch [45]),
    .d(\cu_ru/sscratch [45]),
    .o(_al_u6921_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6922 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [45]),
    .d(\cu_ru/stvec [45]),
    .o(_al_u6922_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6923 (
    .a(_al_u6920_o),
    .b(_al_u6921_o),
    .c(_al_u6922_o),
    .o(_al_u6923_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6924 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[45]),
    .d(\cu_ru/mtvec [45]),
    .o(_al_u6924_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6925 (
    .a(_al_u6918_o),
    .b(_al_u6919_o),
    .c(_al_u6923_o),
    .d(_al_u6924_o),
    .o(csr_data[45]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6926 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [44]),
    .d(\cu_ru/stval [44]),
    .o(_al_u6926_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6927 (
    .a(_al_u6763_o),
    .b(_al_u6926_o),
    .c(\cu_ru/minstret [44]),
    .o(_al_u6927_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6928 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [44]),
    .d(\cu_ru/stvec [44]),
    .o(_al_u6928_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6929 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [44]),
    .d(\cu_ru/mscratch [44]),
    .o(_al_u6929_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6930 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [44]),
    .d(\cu_ru/sscratch [44]),
    .o(_al_u6930_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6931 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [44]),
    .d(\cu_ru/mtval [44]),
    .o(_al_u6931_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6932 (
    .a(_al_u6929_o),
    .b(_al_u6930_o),
    .c(_al_u6931_o),
    .o(_al_u6932_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6933 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[44]),
    .d(\cu_ru/mtvec [44]),
    .o(_al_u6933_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u6934 (
    .a(_al_u6927_o),
    .b(_al_u6928_o),
    .c(_al_u6932_o),
    .d(_al_u6933_o),
    .o(csr_data[44]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h3120))
    _al_u6935 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(_al_u2842_o),
    .c(priv[1]),
    .d(\cu_ru/mstatus [8]),
    .o(_al_u6935_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6936 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mstatus [8]),
    .o(_al_u6936_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((~C*~A))*~(B)+~D*(~C*~A)*~(B)+~(~D)*(~C*~A)*B+~D*(~C*~A)*B)"),
    .INIT(16'hfbc8))
    _al_u6937 (
    .a(_al_u6935_o),
    .b(\cu_ru/m_s_status/u34_sel_is_0_o ),
    .c(_al_u6936_o),
    .d(data_csr[8]),
    .o(\cu_ru/m_s_status/n46 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u6938 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/mstatus [5]),
    .o(_al_u6938_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u6939 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(_al_u6938_o),
    .c(_al_u2844_o),
    .d(\cu_ru/mstatus [1]),
    .o(_al_u6939_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u6940 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mstatus [1]),
    .o(_al_u6940_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B)"),
    .INIT(16'h3704))
    _al_u6941 (
    .a(_al_u6939_o),
    .b(\cu_ru/m_s_status/u34_sel_is_0_o ),
    .c(_al_u6940_o),
    .d(data_csr[1]),
    .o(\cu_ru/m_s_status/n36 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h3120))
    _al_u6942 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(_al_u2842_o),
    .c(\cu_ru/mstatus [1]),
    .d(\cu_ru/mstatus [5]),
    .o(_al_u6942_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u6943 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mstatus [5]),
    .o(_al_u6943_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((~C*~A))*~(B)+~D*(~C*~A)*~(B)+~(~D)*(~C*~A)*B+~D*(~C*~A)*B)"),
    .INIT(16'hfbc8))
    _al_u6944 (
    .a(_al_u6942_o),
    .b(\cu_ru/m_s_status/u34_sel_is_0_o ),
    .c(_al_u6943_o),
    .d(data_csr[5]),
    .o(\cu_ru/m_s_status/n44 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u6945 (
    .a(id_ins[28]),
    .b(id_ins[27]),
    .c(id_ins[26]),
    .o(_al_u6945_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6946 (
    .a(_al_u3397_o),
    .b(_al_u3399_o),
    .c(_al_u6945_o),
    .o(\cu_ru/read_satp_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6947 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[63]),
    .d(\cu_ru/sscratch [63]),
    .o(_al_u6947_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6948 (
    .a(_al_u6947_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [63]),
    .o(_al_u6948_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6949 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [63]),
    .d(\cu_ru/mcause [63]),
    .o(_al_u6949_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6950 (
    .a(_al_u6948_o),
    .b(_al_u6949_o),
    .c(\cu_ru/read_mscratch_sel_lutinv ),
    .d(\cu_ru/mscratch [63]),
    .o(_al_u6950_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6951 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[63]),
    .d(\cu_ru/mtvec [63]),
    .o(_al_u6951_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6952 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [63]),
    .d(\cu_ru/mtval [63]),
    .o(_al_u6952_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6953 (
    .a(_al_u6950_o),
    .b(_al_u6951_o),
    .c(_al_u6952_o),
    .o(_al_u6953_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6954 (
    .a(_al_u6788_o),
    .b(_al_u6763_o),
    .c(\cu_ru/minstret [63]),
    .d(\cu_ru/mcycle [63]),
    .o(_al_u6954_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6955 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [63]),
    .d(\cu_ru/stvec [63]),
    .o(_al_u6955_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u6956 (
    .a(_al_u6953_o),
    .b(_al_u6954_o),
    .c(_al_u6955_o),
    .o(csr_data[63]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6957 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[62]),
    .d(\cu_ru/sscratch [62]),
    .o(_al_u6957_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6958 (
    .a(_al_u6763_o),
    .b(_al_u6957_o),
    .c(\cu_ru/minstret [62]),
    .o(_al_u6958_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6959 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [62]),
    .d(\cu_ru/mscratch [62]),
    .o(_al_u6959_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6960 (
    .a(_al_u6958_o),
    .b(_al_u6959_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [62]),
    .o(_al_u6960_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6961 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [62]),
    .d(\cu_ru/stvec [62]),
    .o(_al_u6961_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6962 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[62]),
    .d(\cu_ru/mtval [62]),
    .o(_al_u6962_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6963 (
    .a(_al_u6960_o),
    .b(_al_u6961_o),
    .c(_al_u6962_o),
    .o(_al_u6963_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6964 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [62]),
    .d(\cu_ru/stval [62]),
    .o(_al_u6964_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6965 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [62]),
    .d(\cu_ru/mtvec [62]),
    .o(_al_u6965_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u6966 (
    .a(_al_u6963_o),
    .b(_al_u6964_o),
    .c(_al_u6965_o),
    .o(csr_data[62]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6967 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[61]),
    .d(\cu_ru/sscratch [61]),
    .o(_al_u6967_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6968 (
    .a(_al_u6967_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [61]),
    .o(_al_u6968_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6969 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [61]),
    .d(\cu_ru/mscratch [61]),
    .o(_al_u6969_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6970 (
    .a(_al_u6968_o),
    .b(_al_u6969_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [61]),
    .o(_al_u6970_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6971 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[61]),
    .d(\cu_ru/mtvec [61]),
    .o(_al_u6971_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6972 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [61]),
    .d(\cu_ru/mtval [61]),
    .o(_al_u6972_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6973 (
    .a(_al_u6970_o),
    .b(_al_u6971_o),
    .c(_al_u6972_o),
    .o(_al_u6973_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6974 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/minstret [61]),
    .d(\cu_ru/stvec [61]),
    .o(_al_u6974_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6975 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/mcycle [61]),
    .d(\cu_ru/sepc [61]),
    .o(_al_u6975_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u6976 (
    .a(_al_u6973_o),
    .b(_al_u6974_o),
    .c(_al_u6975_o),
    .o(csr_data[61]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6977 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[60]),
    .d(\cu_ru/sscratch [60]),
    .o(_al_u6977_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u6978 (
    .a(_al_u6763_o),
    .b(_al_u6977_o),
    .c(\cu_ru/minstret [60]),
    .o(_al_u6978_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6979 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [60]),
    .d(\cu_ru/mscratch [60]),
    .o(_al_u6979_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6980 (
    .a(_al_u6978_o),
    .b(_al_u6979_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [60]),
    .o(_al_u6980_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u6981 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [60]),
    .d(\cu_ru/stvec [60]),
    .o(_al_u6981_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6982 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[60]),
    .d(\cu_ru/mtval [60]),
    .o(_al_u6982_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6983 (
    .a(_al_u6980_o),
    .b(_al_u6981_o),
    .c(_al_u6982_o),
    .o(_al_u6983_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6984 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [60]),
    .d(\cu_ru/stval [60]),
    .o(_al_u6984_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6985 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [60]),
    .d(\cu_ru/mtvec [60]),
    .o(_al_u6985_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u6986 (
    .a(_al_u6983_o),
    .b(_al_u6984_o),
    .c(_al_u6985_o),
    .o(csr_data[60]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6987 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [43]),
    .d(\cu_ru/mscratch [43]),
    .o(_al_u6987_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6988 (
    .a(_al_u6987_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [43]),
    .o(_al_u6988_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6989 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[43]),
    .d(\cu_ru/sscratch [43]),
    .o(_al_u6989_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u6990 (
    .a(_al_u6988_o),
    .b(_al_u6989_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [43]),
    .o(_al_u6990_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6991 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stvec [43]),
    .d(\cu_ru/mtvec [43]),
    .o(_al_u6991_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6992 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/stval [43]),
    .d(\cu_ru/mtval [43]),
    .o(_al_u6992_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u6993 (
    .a(_al_u6990_o),
    .b(_al_u6991_o),
    .c(_al_u6992_o),
    .o(_al_u6993_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u6994 (
    .a(_al_u6788_o),
    .b(_al_u6763_o),
    .c(\cu_ru/minstret [43]),
    .d(\cu_ru/mcycle [43]),
    .o(_al_u6994_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6995 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(mtime_pad[43]),
    .d(\cu_ru/mepc [43]),
    .o(_al_u6995_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u6996 (
    .a(_al_u6993_o),
    .b(_al_u6994_o),
    .c(_al_u6995_o),
    .o(csr_data[43]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u6997 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [42]),
    .d(\cu_ru/mcause [42]),
    .o(_al_u6997_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u6998 (
    .a(_al_u6997_o),
    .b(\cu_ru/read_instret_sel_lutinv ),
    .c(\cu_ru/minstret [42]),
    .o(_al_u6998_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u6999 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/minstret [42]),
    .d(\cu_ru/sscratch [42]),
    .o(_al_u6999_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7000 (
    .a(\cu_ru/read_mscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[42]),
    .d(\cu_ru/mscratch [42]),
    .o(_al_u7000_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7001 (
    .a(_al_u6998_o),
    .b(_al_u6999_o),
    .c(_al_u7000_o),
    .o(_al_u7001_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7002 (
    .a(\cu_ru/read_sepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/sepc [42]),
    .d(\cu_ru/stvec [42]),
    .o(_al_u7002_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7003 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/stval [42]),
    .d(\cu_ru/mtval [42]),
    .o(_al_u7003_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7004 (
    .a(_al_u7001_o),
    .b(_al_u7002_o),
    .c(_al_u7003_o),
    .o(_al_u7004_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7005 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mcycle [42]),
    .d(\cu_ru/mepc [42]),
    .o(_al_u7005_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7006 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[42]),
    .d(\cu_ru/mtvec [42]),
    .o(_al_u7006_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7007 (
    .a(_al_u7004_o),
    .b(_al_u7005_o),
    .c(_al_u7006_o),
    .o(csr_data[42]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7008 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[41]),
    .d(\cu_ru/sscratch [41]),
    .o(_al_u7008_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7009 (
    .a(_al_u6763_o),
    .b(_al_u7008_o),
    .c(\cu_ru/minstret [41]),
    .o(_al_u7009_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7010 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [41]),
    .d(\cu_ru/mscratch [41]),
    .o(_al_u7010_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7011 (
    .a(_al_u7009_o),
    .b(_al_u7010_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [41]),
    .o(_al_u7011_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7012 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [41]),
    .d(\cu_ru/stvec [41]),
    .o(_al_u7012_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7013 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[41]),
    .d(\cu_ru/mtval [41]),
    .o(_al_u7013_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7014 (
    .a(_al_u7011_o),
    .b(_al_u7012_o),
    .c(_al_u7013_o),
    .o(_al_u7014_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7015 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [41]),
    .d(\cu_ru/stval [41]),
    .o(_al_u7015_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7016 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [41]),
    .d(\cu_ru/mtvec [41]),
    .o(_al_u7016_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7017 (
    .a(_al_u7014_o),
    .b(_al_u7015_o),
    .c(_al_u7016_o),
    .o(csr_data[41]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7018 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[40]),
    .d(\cu_ru/sscratch [40]),
    .o(_al_u7018_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7019 (
    .a(_al_u6763_o),
    .b(_al_u7018_o),
    .c(\cu_ru/minstret [40]),
    .o(_al_u7019_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7020 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [40]),
    .d(\cu_ru/mscratch [40]),
    .o(_al_u7020_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7021 (
    .a(_al_u7019_o),
    .b(_al_u7020_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [40]),
    .o(_al_u7021_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7022 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [40]),
    .d(\cu_ru/stvec [40]),
    .o(_al_u7022_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7023 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[40]),
    .d(\cu_ru/mtval [40]),
    .o(_al_u7023_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7024 (
    .a(_al_u7021_o),
    .b(_al_u7022_o),
    .c(_al_u7023_o),
    .o(_al_u7024_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7025 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [40]),
    .d(\cu_ru/stval [40]),
    .o(_al_u7025_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7026 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [40]),
    .d(\cu_ru/mtvec [40]),
    .o(_al_u7026_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7027 (
    .a(_al_u7024_o),
    .b(_al_u7025_o),
    .c(_al_u7026_o),
    .o(csr_data[40]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7028 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[39]),
    .d(\cu_ru/sscratch [39]),
    .o(_al_u7028_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7029 (
    .a(_al_u6763_o),
    .b(_al_u7028_o),
    .c(\cu_ru/minstret [39]),
    .o(_al_u7029_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7030 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [39]),
    .d(\cu_ru/mscratch [39]),
    .o(_al_u7030_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7031 (
    .a(_al_u7029_o),
    .b(_al_u7030_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [39]),
    .o(_al_u7031_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u7032 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[39]),
    .d(\cu_ru/mcycle [39]),
    .o(_al_u7032_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7033 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stvec [39]),
    .d(\cu_ru/mtvec [39]),
    .o(_al_u7033_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7034 (
    .a(_al_u7031_o),
    .b(_al_u7032_o),
    .c(_al_u7033_o),
    .o(_al_u7034_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7035 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [39]),
    .d(\cu_ru/mtval [39]),
    .o(_al_u7035_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7036 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [39]),
    .d(\cu_ru/stval [39]),
    .o(_al_u7036_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7037 (
    .a(_al_u7034_o),
    .b(_al_u7035_o),
    .c(_al_u7036_o),
    .o(csr_data[39]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7038 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mscratch [38]),
    .d(\cu_ru/sscratch [38]),
    .o(_al_u7038_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7039 (
    .a(_al_u6763_o),
    .b(_al_u7038_o),
    .c(\cu_ru/minstret [38]),
    .o(_al_u7039_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7040 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[38]),
    .d(\cu_ru/scause [38]),
    .o(_al_u7040_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7041 (
    .a(_al_u7039_o),
    .b(_al_u7040_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [38]),
    .o(_al_u7041_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7042 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mtval [38]),
    .d(\cu_ru/stvec [38]),
    .o(_al_u7042_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7043 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[38]),
    .d(\cu_ru/stval [38]),
    .o(_al_u7043_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7044 (
    .a(_al_u7041_o),
    .b(_al_u7042_o),
    .c(_al_u7043_o),
    .o(_al_u7044_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7045 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/mcycle [38]),
    .d(\cu_ru/sepc [38]),
    .o(_al_u7045_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7046 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [38]),
    .d(\cu_ru/mtvec [38]),
    .o(_al_u7046_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7047 (
    .a(_al_u7044_o),
    .b(_al_u7045_o),
    .c(_al_u7046_o),
    .o(csr_data[38]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7048 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[37]),
    .d(\cu_ru/sscratch [37]),
    .o(_al_u7048_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7049 (
    .a(_al_u6763_o),
    .b(_al_u7048_o),
    .c(\cu_ru/minstret [37]),
    .o(_al_u7049_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7050 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [37]),
    .d(\cu_ru/mcause [37]),
    .o(_al_u7050_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7051 (
    .a(_al_u7049_o),
    .b(_al_u7050_o),
    .c(\cu_ru/read_mscratch_sel_lutinv ),
    .d(\cu_ru/mscratch [37]),
    .o(_al_u7051_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7052 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [37]),
    .d(\cu_ru/stvec [37]),
    .o(_al_u7052_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7053 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[37]),
    .d(\cu_ru/mtval [37]),
    .o(_al_u7053_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7054 (
    .a(_al_u7051_o),
    .b(_al_u7052_o),
    .c(_al_u7053_o),
    .o(_al_u7054_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7055 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [37]),
    .d(\cu_ru/stval [37]),
    .o(_al_u7055_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7056 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [37]),
    .d(\cu_ru/mtvec [37]),
    .o(_al_u7056_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7057 (
    .a(_al_u7054_o),
    .b(_al_u7055_o),
    .c(_al_u7056_o),
    .o(csr_data[37]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7058 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[36]),
    .d(\cu_ru/scause [36]),
    .o(_al_u7058_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7059 (
    .a(_al_u7058_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [36]),
    .o(_al_u7059_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7060 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [36]),
    .d(\cu_ru/sscratch [36]),
    .o(_al_u7060_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7061 (
    .a(_al_u7059_o),
    .b(_al_u7060_o),
    .c(\cu_ru/read_mscratch_sel_lutinv ),
    .d(\cu_ru/mscratch [36]),
    .o(_al_u7061_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7062 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_mtvec_sel_lutinv ),
    .c(\cu_ru/mcycle [36]),
    .d(\cu_ru/mtvec [36]),
    .o(_al_u7062_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7063 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[36]),
    .d(\cu_ru/stval [36]),
    .o(_al_u7063_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7064 (
    .a(_al_u7061_o),
    .b(_al_u7062_o),
    .c(_al_u7063_o),
    .o(_al_u7064_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7065 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/minstret [36]),
    .d(\cu_ru/stvec [36]),
    .o(_al_u7065_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7066 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [36]),
    .d(\cu_ru/mtval [36]),
    .o(_al_u7066_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7067 (
    .a(_al_u7064_o),
    .b(_al_u7065_o),
    .c(_al_u7066_o),
    .o(csr_data[36]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7068 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[31]),
    .d(\cu_ru/sscratch [31]),
    .o(_al_u7068_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7069 (
    .a(_al_u6763_o),
    .b(_al_u7068_o),
    .c(\cu_ru/minstret [31]),
    .o(_al_u7069_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7070 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [31]),
    .d(\cu_ru/mscratch [31]),
    .o(_al_u7070_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7071 (
    .a(_al_u7069_o),
    .b(_al_u7070_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [31]),
    .o(_al_u7071_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7072 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_mtvec_sel_lutinv ),
    .c(\cu_ru/mcycle [31]),
    .d(\cu_ru/mtvec [31]),
    .o(_al_u7072_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7073 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(mtime_pad[31]),
    .d(\cu_ru/stvec [31]),
    .o(_al_u7073_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7074 (
    .a(_al_u7071_o),
    .b(_al_u7072_o),
    .c(_al_u7073_o),
    .o(_al_u7074_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7075 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [31]),
    .d(\cu_ru/mtval [31]),
    .o(_al_u7075_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7076 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [31]),
    .d(\cu_ru/stval [31]),
    .o(_al_u7076_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7077 (
    .a(_al_u7074_o),
    .b(_al_u7075_o),
    .c(_al_u7076_o),
    .o(csr_data[31]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7078 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[29]),
    .d(\cu_ru/sscratch [29]),
    .o(_al_u7078_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7079 (
    .a(_al_u6763_o),
    .b(_al_u7078_o),
    .c(\cu_ru/minstret [29]),
    .o(_al_u7079_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7080 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [29]),
    .d(\cu_ru/mscratch [29]),
    .o(_al_u7080_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7081 (
    .a(_al_u7079_o),
    .b(_al_u7080_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [29]),
    .o(_al_u7081_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7082 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [29]),
    .d(\cu_ru/stvec [29]),
    .o(_al_u7082_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7083 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[29]),
    .d(\cu_ru/mtval [29]),
    .o(_al_u7083_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7084 (
    .a(_al_u7081_o),
    .b(_al_u7082_o),
    .c(_al_u7083_o),
    .o(_al_u7084_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7085 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [29]),
    .d(\cu_ru/stval [29]),
    .o(_al_u7085_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7086 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [29]),
    .d(\cu_ru/mtvec [29]),
    .o(_al_u7086_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7087 (
    .a(_al_u7084_o),
    .b(_al_u7085_o),
    .c(_al_u7086_o),
    .o(csr_data[29]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7088 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[27]),
    .d(\cu_ru/sscratch [27]),
    .o(_al_u7088_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7089 (
    .a(_al_u6763_o),
    .b(_al_u7088_o),
    .c(\cu_ru/minstret [27]),
    .o(_al_u7089_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7090 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [27]),
    .d(\cu_ru/mscratch [27]),
    .o(_al_u7090_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7091 (
    .a(_al_u7089_o),
    .b(_al_u7090_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [27]),
    .o(_al_u7091_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7092 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_mtvec_sel_lutinv ),
    .c(\cu_ru/mcycle [27]),
    .d(\cu_ru/mtvec [27]),
    .o(_al_u7092_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7093 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(mtime_pad[27]),
    .d(\cu_ru/stvec [27]),
    .o(_al_u7093_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7094 (
    .a(_al_u7091_o),
    .b(_al_u7092_o),
    .c(_al_u7093_o),
    .o(_al_u7094_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7095 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [27]),
    .d(\cu_ru/mtval [27]),
    .o(_al_u7095_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7096 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [27]),
    .d(\cu_ru/stval [27]),
    .o(_al_u7096_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7097 (
    .a(_al_u7094_o),
    .b(_al_u7095_o),
    .c(_al_u7096_o),
    .o(csr_data[27]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7098 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [26]),
    .d(\cu_ru/sscratch [26]),
    .o(_al_u7098_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7099 (
    .a(_al_u7098_o),
    .b(\cu_ru/read_instret_sel_lutinv ),
    .c(\cu_ru/minstret [26]),
    .o(_al_u7099_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7100 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/minstret [26]),
    .d(\cu_ru/scause [26]),
    .o(_al_u7100_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7101 (
    .a(\cu_ru/read_mscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[26]),
    .d(\cu_ru/mscratch [26]),
    .o(_al_u7101_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7102 (
    .a(_al_u7099_o),
    .b(_al_u7100_o),
    .c(_al_u7101_o),
    .o(_al_u7102_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7103 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [26]),
    .d(\cu_ru/mtvec [26]),
    .o(_al_u7103_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7104 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stval [26]),
    .d(\cu_ru/stvec [26]),
    .o(_al_u7104_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7105 (
    .a(_al_u7102_o),
    .b(_al_u7103_o),
    .c(_al_u7104_o),
    .o(_al_u7105_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7106 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mcycle [26]),
    .d(\cu_ru/mepc [26]),
    .o(_al_u7106_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7107 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[26]),
    .d(\cu_ru/mtval [26]),
    .o(_al_u7107_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7108 (
    .a(_al_u7105_o),
    .b(_al_u7106_o),
    .c(_al_u7107_o),
    .o(csr_data[26]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7109 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[24]),
    .d(\cu_ru/sscratch [24]),
    .o(_al_u7109_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7110 (
    .a(_al_u7109_o),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [24]),
    .o(_al_u7110_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7111 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/minstret [24]),
    .d(\cu_ru/scause [24]),
    .o(_al_u7111_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7112 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/minstret [24]),
    .d(\cu_ru/mscratch [24]),
    .o(_al_u7112_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7113 (
    .a(_al_u7110_o),
    .b(_al_u7111_o),
    .c(_al_u7112_o),
    .o(_al_u7113_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7114 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [24]),
    .d(\cu_ru/mtvec [24]),
    .o(_al_u7114_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7115 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stval [24]),
    .d(\cu_ru/stvec [24]),
    .o(_al_u7115_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7116 (
    .a(_al_u7113_o),
    .b(_al_u7114_o),
    .c(_al_u7115_o),
    .o(_al_u7116_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u7117 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[24]),
    .d(\cu_ru/mcycle [24]),
    .o(_al_u7117_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7118 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [24]),
    .d(\cu_ru/mtval [24]),
    .o(_al_u7118_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7119 (
    .a(_al_u7116_o),
    .b(_al_u7117_o),
    .c(_al_u7118_o),
    .o(csr_data[24]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7120 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[23]),
    .d(\cu_ru/sscratch [23]),
    .o(_al_u7120_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7121 (
    .a(_al_u7120_o),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [23]),
    .o(_al_u7121_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7122 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/minstret [23]),
    .d(\cu_ru/scause [23]),
    .o(_al_u7122_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7123 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/minstret [23]),
    .d(\cu_ru/mscratch [23]),
    .o(_al_u7123_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7124 (
    .a(_al_u7121_o),
    .b(_al_u7122_o),
    .c(_al_u7123_o),
    .o(_al_u7124_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7125 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [23]),
    .d(\cu_ru/mtvec [23]),
    .o(_al_u7125_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7126 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stval [23]),
    .d(\cu_ru/stvec [23]),
    .o(_al_u7126_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7127 (
    .a(_al_u7124_o),
    .b(_al_u7125_o),
    .c(_al_u7126_o),
    .o(_al_u7127_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u7128 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[23]),
    .d(\cu_ru/mcycle [23]),
    .o(_al_u7128_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7129 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [23]),
    .d(\cu_ru/mtval [23]),
    .o(_al_u7129_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7130 (
    .a(_al_u7127_o),
    .b(_al_u7128_o),
    .c(_al_u7129_o),
    .o(csr_data[23]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7131 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[16]),
    .d(\cu_ru/sscratch [16]),
    .o(_al_u7131_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7132 (
    .a(_al_u6763_o),
    .b(_al_u7131_o),
    .c(\cu_ru/minstret [16]),
    .o(_al_u7132_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7133 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [16]),
    .d(\cu_ru/mcause [16]),
    .o(_al_u7133_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7134 (
    .a(_al_u7132_o),
    .b(_al_u7133_o),
    .c(\cu_ru/read_mscratch_sel_lutinv ),
    .d(\cu_ru/mscratch [16]),
    .o(_al_u7134_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7135 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mcycle [16]),
    .d(\cu_ru/stvec [16]),
    .o(_al_u7135_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7136 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[16]),
    .d(\cu_ru/mtval [16]),
    .o(_al_u7136_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7137 (
    .a(_al_u7134_o),
    .b(_al_u7135_o),
    .c(_al_u7136_o),
    .o(_al_u7137_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7138 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [16]),
    .d(\cu_ru/stval [16]),
    .o(_al_u7138_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7139 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [16]),
    .d(\cu_ru/mtvec [16]),
    .o(_al_u7139_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7140 (
    .a(_al_u7137_o),
    .b(_al_u7138_o),
    .c(_al_u7139_o),
    .o(csr_data[16]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u7141 (
    .a(_al_u3927_o),
    .b(_al_u3925_o),
    .c(_al_u4064_o),
    .o(_al_u7141_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u7142 (
    .a(\ins_dec/op_load ),
    .b(id_system),
    .o(_al_u7142_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7143 (
    .a(_al_u3956_o),
    .b(_al_u4161_o),
    .c(_al_u7141_o),
    .d(_al_u7142_o),
    .o(\ins_dec/dec_ins_dec_fault_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u7144 (
    .a(_al_u3399_o),
    .b(_al_u3400_o),
    .c(id_ins[25]),
    .o(\ins_dec/funct7_8_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfcc7))
    _al_u7145 (
    .a(\ins_dec/n80_lutinv ),
    .b(priv[0]),
    .c(priv[1]),
    .d(priv[3]),
    .o(_al_u7145_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7146 (
    .a(id_system),
    .b(tw),
    .o(_al_u7146_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(~C*A))"),
    .INIT(16'h31f5))
    _al_u7147 (
    .a(\ins_dec/n239 ),
    .b(\ins_dec/funct7_8_lutinv ),
    .c(_al_u7145_o),
    .d(_al_u7146_o),
    .o(_al_u7147_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~A*~(D*C))"),
    .INIT(16'hfbbb))
    _al_u7148 (
    .a(\ins_dec/dec_ins_dec_fault_lutinv ),
    .b(_al_u7147_o),
    .c(tvm),
    .d(\ins_dec/ins_sfencevma ),
    .o(id_ill_ins));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*A))"),
    .INIT(16'h1333))
    _al_u7149 (
    .a(_al_u2705_o),
    .b(_al_u3407_o),
    .c(_al_u4195_o),
    .d(\biu/bus_unit/mmu/statu [0]),
    .o(_al_u7149_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u7150 (
    .a(_al_u3944_o),
    .b(\biu/cache_ctrl_logic/statu [0]),
    .c(\biu/cache_ctrl_logic/statu [1]),
    .o(_al_u7150_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hceea))
    _al_u7151 (
    .a(_al_u2835_o),
    .b(_al_u2838_o),
    .c(\biu/cache_ctrl_logic/statu [0]),
    .d(\biu/cache_ctrl_logic/statu [1]),
    .o(_al_u7151_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*~(D*~C)))"),
    .INIT(16'h4544))
    _al_u7152 (
    .a(\biu/cache_ctrl_logic/n97_lutinv ),
    .b(_al_u7150_o),
    .c(_al_u7151_o),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(_al_u7152_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*C*B))"),
    .INIT(16'h5515))
    _al_u7153 (
    .a(_al_u3224_o),
    .b(_al_u2847_o),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .d(\biu/cache_ctrl_logic/statu [4]),
    .o(\biu/cache_ctrl_logic/mux31_b4_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(D*A)))"),
    .INIT(16'hb030))
    _al_u7154 (
    .a(_al_u7149_o),
    .b(_al_u7152_o),
    .c(\biu/cache_ctrl_logic/mux31_b4_sel_is_2_o ),
    .d(_al_u7150_o),
    .o(_al_u7154_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7155 (
    .a(_al_u7149_o),
    .b(\biu/cache_ctrl_logic/mux31_b4_sel_is_2_o ),
    .o(_al_u7155_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D*A)))"),
    .INIT(16'h0b03))
    _al_u7156 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u7154_o),
    .c(_al_u7155_o),
    .d(\biu/cache_ctrl_logic/n97_lutinv ),
    .o(_al_u7156_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u7157 (
    .a(_al_u2705_o),
    .b(_al_u4195_o),
    .c(\biu/bus_unit/mmu/statu [0]),
    .o(_al_u7157_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(~D*~C)))"),
    .INIT(16'h444c))
    _al_u7158 (
    .a(_al_u7157_o),
    .b(\biu/cache_ctrl_logic/n75_lutinv ),
    .c(read),
    .d(write),
    .o(_al_u7158_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u7159 (
    .a(_al_u7149_o),
    .b(_al_u6257_o),
    .c(\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ),
    .d(\biu/cache_ctrl_logic/n75_lutinv ),
    .o(_al_u7159_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7160 (
    .a(_al_u7149_o),
    .b(_al_u2885_o),
    .c(\biu/cache_ctrl_logic/statu [1]),
    .o(_al_u7160_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(C*~A)))"),
    .INIT(16'h00dc))
    _al_u7161 (
    .a(_al_u7156_o),
    .b(_al_u7158_o),
    .c(_al_u7159_o),
    .d(_al_u7160_o),
    .o(_al_u7161_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7162 (
    .a(_al_u6426_o),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .o(_al_u7162_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7163 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u7149_o),
    .o(_al_u7163_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7164 (
    .a(cacheability_block_pad[21]),
    .b(cacheability_block_pad[1]),
    .c(\biu/paddress [33]),
    .d(\biu/paddress [53]),
    .o(_al_u7164_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u7165 (
    .a(cacheability_block_pad[22]),
    .b(cacheability_block_pad[12]),
    .c(\biu/paddress [44]),
    .d(\biu/paddress [54]),
    .o(_al_u7165_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u7166 (
    .a(_al_u7164_o),
    .b(_al_u7165_o),
    .c(cacheability_block_pad[10]),
    .d(\biu/paddress [42]),
    .o(_al_u7166_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7167 (
    .a(cacheability_block_pad[26]),
    .b(cacheability_block_pad[18]),
    .c(\biu/paddress [50]),
    .d(\biu/paddress [58]),
    .o(_al_u7167_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7168 (
    .a(cacheability_block_pad[2]),
    .b(cacheability_block_pad[0]),
    .c(\biu/paddress [32]),
    .d(\biu/paddress [34]),
    .o(_al_u7168_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7169 (
    .a(_al_u7166_o),
    .b(_al_u7167_o),
    .c(_al_u7168_o),
    .o(_al_u7169_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7170 (
    .a(cacheability_block_pad[30]),
    .b(cacheability_block_pad[28]),
    .c(\biu/paddress [60]),
    .d(\biu/paddress [62]),
    .o(_al_u7170_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u7171 (
    .a(_al_u3411_o),
    .b(_al_u7170_o),
    .c(cacheability_block_pad[29]),
    .d(\biu/paddress [61]),
    .o(_al_u7171_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7172 (
    .a(cacheability_block_pad[24]),
    .b(cacheability_block_pad[20]),
    .c(\biu/paddress [52]),
    .d(\biu/paddress [56]),
    .o(_al_u7172_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u7173 (
    .a(cacheability_block_pad[22]),
    .b(cacheability_block_pad[12]),
    .c(\biu/paddress [44]),
    .d(\biu/paddress [54]),
    .o(_al_u7173_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u7174 (
    .a(_al_u7172_o),
    .b(_al_u7173_o),
    .c(cacheability_block_pad[13]),
    .d(\biu/paddress [45]),
    .o(_al_u7174_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7175 (
    .a(_al_u7169_o),
    .b(_al_u7171_o),
    .c(_al_u7174_o),
    .o(_al_u7175_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7176 (
    .a(cacheability_block_pad[27]),
    .b(cacheability_block_pad[23]),
    .c(\biu/paddress [55]),
    .d(\biu/paddress [59]),
    .o(_al_u7176_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7177 (
    .a(cacheability_block_pad[19]),
    .b(cacheability_block_pad[8]),
    .c(\biu/paddress [40]),
    .d(\biu/paddress [51]),
    .o(_al_u7177_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7178 (
    .a(cacheability_block_pad[25]),
    .b(cacheability_block_pad[3]),
    .c(\biu/paddress [35]),
    .d(\biu/paddress [57]),
    .o(_al_u7178_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7179 (
    .a(cacheability_block_pad[7]),
    .b(cacheability_block_pad[4]),
    .c(\biu/paddress [36]),
    .d(\biu/paddress [39]),
    .o(_al_u7179_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7180 (
    .a(_al_u7176_o),
    .b(_al_u7177_o),
    .c(_al_u7178_o),
    .d(_al_u7179_o),
    .o(_al_u7180_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7181 (
    .a(cacheability_block_pad[15]),
    .b(cacheability_block_pad[9]),
    .c(\biu/paddress [41]),
    .d(\biu/paddress [47]),
    .o(_al_u7181_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u7182 (
    .a(_al_u7180_o),
    .b(_al_u7181_o),
    .c(cacheability_block_pad[6]),
    .d(\biu/paddress [38]),
    .o(_al_u7182_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(~D*A))"),
    .INIT(16'hcf45))
    _al_u7183 (
    .a(cacheability_block_pad[31]),
    .b(cacheability_block_pad[17]),
    .c(\biu/paddress [49]),
    .d(\biu/paddress [63]),
    .o(_al_u7183_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(~D*A))"),
    .INIT(16'hcf45))
    _al_u7184 (
    .a(cacheability_block_pad[17]),
    .b(cacheability_block_pad[16]),
    .c(\biu/paddress [48]),
    .d(\biu/paddress [49]),
    .o(_al_u7184_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u7185 (
    .a(cacheability_block_pad[16]),
    .b(cacheability_block_pad[11]),
    .c(\biu/paddress [43]),
    .d(\biu/paddress [48]),
    .o(_al_u7185_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u7186 (
    .a(cacheability_block_pad[31]),
    .b(cacheability_block_pad[11]),
    .c(\biu/paddress [43]),
    .d(\biu/paddress [63]),
    .o(_al_u7186_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7187 (
    .a(_al_u7183_o),
    .b(_al_u7184_o),
    .c(_al_u7185_o),
    .d(_al_u7186_o),
    .o(_al_u7187_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u7188 (
    .a(cacheability_block_pad[14]),
    .b(cacheability_block_pad[5]),
    .c(\biu/paddress [37]),
    .d(\biu/paddress [46]),
    .o(_al_u7188_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7189 (
    .a(_al_u7175_o),
    .b(_al_u7182_o),
    .c(_al_u7187_o),
    .d(_al_u7188_o),
    .o(\biu/cacheable ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7190 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(\biu/cacheable ),
    .o(_al_u7190_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7191 (
    .a(_al_u7157_o),
    .b(\biu/bus_unit/mmu/n19_lutinv ),
    .o(_al_u7191_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*~(~C*~B)))"),
    .INIT(16'h0155))
    _al_u7192 (
    .a(_al_u7162_o),
    .b(_al_u7163_o),
    .c(_al_u7190_o),
    .d(_al_u7191_o),
    .o(_al_u7192_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7193 (
    .a(_al_u6321_o),
    .b(\biu/cache_ctrl_logic/n55_lutinv ),
    .c(write),
    .o(_al_u7193_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7194 (
    .a(_al_u7161_o),
    .b(_al_u7192_o),
    .c(_al_u7193_o),
    .o(\biu/cache_ctrl_logic/n127[4]_d ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7195 (
    .a(_al_u2835_o),
    .b(_al_u3209_o),
    .o(_al_u7195_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*A*~(C*B))"),
    .INIT(16'hffd5))
    _al_u7196 (
    .a(_al_u6724_o),
    .b(_al_u2910_o),
    .c(_al_u6725_o),
    .d(_al_u7195_o),
    .o(\exu/n92 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7197 (
    .a(\biu/cache_ctrl_logic/n75_lutinv ),
    .b(write),
    .o(\biu/bus_unit/mmu/n12_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*~(D*C)))"),
    .INIT(16'h5444))
    _al_u7198 (
    .a(\biu/bus_unit/mmu/n19_lutinv ),
    .b(\biu/bus_unit/mmu_hwdata [1]),
    .c(\biu/bus_unit/mmu_hwdata [3]),
    .d(mxr),
    .o(_al_u7198_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u7199 (
    .a(\biu/bus_unit/mmu/n19_lutinv ),
    .b(\biu/bus_unit/mmu_hwdata [3]),
    .c(priv[3]),
    .o(_al_u7199_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h10b0))
    _al_u7200 (
    .a(\biu/bus_unit/mmu/n12_lutinv ),
    .b(_al_u7198_o),
    .c(_al_u7199_o),
    .d(\biu/bus_unit/mmu_hwdata [2]),
    .o(_al_u7200_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfcc7))
    _al_u7201 (
    .a(\biu/bus_unit/mmu_hwdata [4]),
    .b(priv[0]),
    .c(priv[1]),
    .d(priv[3]),
    .o(_al_u7201_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u7202 (
    .a(_al_u7200_o),
    .b(_al_u2915_o),
    .c(_al_u7201_o),
    .o(_al_u7202_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u7203 (
    .a(_al_u7202_o),
    .b(\biu/bus_unit/mmu/n37_lutinv ),
    .o(_al_u7203_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u7204 (
    .a(\biu/bus_unit/mmu/statu [0]),
    .b(\biu/bus_unit/mmu/statu [1]),
    .c(\biu/bus_unit/mmu/statu [2]),
    .d(\biu/bus_unit/mmu/statu [3]),
    .o(\biu/bus_unit/mmu/n45_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u7205 (
    .a(_al_u4195_o),
    .b(\biu/bus_unit/mmu/n45_lutinv ),
    .c(hresp_pad),
    .d(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u7205_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u7206 (
    .a(_al_u7203_o),
    .b(_al_u7205_o),
    .c(_al_u2915_o),
    .o(_al_u7206_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u7207 (
    .a(\biu/bus_unit/mmu/n39 [0]),
    .b(\biu/bus_unit/mmu/i [0]),
    .c(\biu/bus_unit/mmu/i [1]),
    .d(\biu/bus_unit/mmu_hwdata [2]),
    .o(\biu/bus_unit/mmu/n2 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7208 (
    .a(\biu/bus_unit/mmu/n2 ),
    .b(\biu/bus_unit/mmu/n37_lutinv ),
    .c(\biu/bus_unit/mmu_hwdata [6]),
    .o(_al_u7208_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7209 (
    .a(_al_u7206_o),
    .b(_al_u7208_o),
    .c(_al_u2964_o),
    .d(hresp_pad),
    .o(\biu/bus_unit/mmu/n54 [3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(~D*~C)))"),
    .INIT(16'h444c))
    _al_u7210 (
    .a(\cu_ru/medeleg_exc_ctrl/n85_neg_lutinv ),
    .b(\cu_ru/medeleg_exc_ctrl/n84_neg_lutinv ),
    .c(_al_u4106_o),
    .d(\cu_ru/medeleg_exc_ctrl/n87_neg_lutinv ),
    .o(_al_u7210_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(~C*~A))"),
    .INIT(16'h00c8))
    _al_u7211 (
    .a(_al_u7210_o),
    .b(\cu_ru/medeleg_exc_ctrl/n80_neg_lutinv ),
    .c(_al_u4126_o),
    .d(_al_u4128_o),
    .o(_al_u7211_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(~B*~A))"),
    .INIT(16'h00e0))
    _al_u7212 (
    .a(_al_u7211_o),
    .b(_al_u4117_o),
    .c(_al_u5099_o),
    .d(_al_u5154_o),
    .o(_al_u7212_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((~D*~A))*~(B)+C*(~D*~A)*~(B)+~(C)*(~D*~A)*B+C*(~D*~A)*B)"),
    .INIT(16'hcf8b))
    _al_u7213 (
    .a(_al_u7212_o),
    .b(_al_u4138_o),
    .c(_al_u4233_o),
    .d(_al_u4141_o),
    .o(\cu_ru/trap_cause [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u7214 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[35]),
    .d(\cu_ru/mcycle [35]),
    .o(_al_u7214_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7215 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [35]),
    .d(\cu_ru/mscratch [35]),
    .o(_al_u7215_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7216 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [35]),
    .d(\cu_ru/sscratch [35]),
    .o(_al_u7216_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7217 (
    .a(_al_u3397_o),
    .b(_al_u6791_o),
    .o(\cu_ru/n90 [32]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u7218 (
    .a(\cu_ru/read_satp_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(satp[35]),
    .o(_al_u7218_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7219 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(_al_u7218_o),
    .c(\cu_ru/stval [35]),
    .o(_al_u7219_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7220 (
    .a(_al_u7215_o),
    .b(_al_u7216_o),
    .c(_al_u7219_o),
    .o(_al_u7220_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7221 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [35]),
    .d(\cu_ru/mtvec [35]),
    .o(_al_u7221_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7222 (
    .a(_al_u7214_o),
    .b(_al_u7220_o),
    .c(_al_u7221_o),
    .o(_al_u7222_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7223 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/minstret [35]),
    .d(\cu_ru/stvec [35]),
    .o(_al_u7223_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7224 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [35]),
    .d(\cu_ru/mtval [35]),
    .o(_al_u7224_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7225 (
    .a(_al_u7222_o),
    .b(_al_u7223_o),
    .c(_al_u7224_o),
    .o(csr_data[35]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u7226 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/scause [34]),
    .o(_al_u7226_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7227 (
    .a(_al_u7226_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mtval [34]),
    .o(_al_u7227_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7228 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mscratch [34]),
    .d(\cu_ru/sscratch [34]),
    .o(_al_u7228_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7229 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[34]),
    .d(\cu_ru/mcause [34]),
    .o(_al_u7229_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7230 (
    .a(_al_u7227_o),
    .b(_al_u7228_o),
    .c(_al_u7229_o),
    .o(_al_u7230_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7231 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mcycle [34]),
    .d(\cu_ru/mepc [34]),
    .o(_al_u7231_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7232 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(mtime_pad[34]),
    .d(\cu_ru/stvec [34]),
    .o(_al_u7232_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7233 (
    .a(_al_u7230_o),
    .b(_al_u7231_o),
    .c(_al_u7232_o),
    .o(_al_u7233_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7234 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/minstret [34]),
    .d(\cu_ru/sepc [34]),
    .o(_al_u7234_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7235 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [34]),
    .d(\cu_ru/mtvec [34]),
    .o(_al_u7235_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7236 (
    .a(_al_u7233_o),
    .b(_al_u7234_o),
    .c(_al_u7235_o),
    .o(csr_data[34]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7237 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [25]),
    .d(\cu_ru/sscratch [25]),
    .o(_al_u7237_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7238 (
    .a(_al_u3400_o),
    .b(id_ins[31]),
    .c(id_ins[30]),
    .d(id_ins[29]),
    .o(_al_u7238_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7239 (
    .a(_al_u7238_o),
    .b(id_ins[20]),
    .o(_al_u7239_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u7240 (
    .a(id_ins[25]),
    .b(id_ins[24]),
    .c(id_ins[23]),
    .o(_al_u7240_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7241 (
    .a(_al_u7239_o),
    .b(_al_u7240_o),
    .c(_al_u3394_o),
    .o(\cu_ru/n82 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u7242 (
    .a(_al_u7237_o),
    .b(\cu_ru/n82 [14]),
    .c(\cu_ru/read_mscratch_sel_lutinv ),
    .d(\cu_ru/mscratch [25]),
    .o(_al_u7242_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7243 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[25]),
    .d(\cu_ru/scause [25]),
    .o(_al_u7243_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7244 (
    .a(_al_u7242_o),
    .b(_al_u7243_o),
    .c(\cu_ru/read_sepc_sel_lutinv ),
    .d(\cu_ru/sepc [25]),
    .o(_al_u7244_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u7245 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[25]),
    .d(\cu_ru/minstret [25]),
    .o(_al_u7245_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7246 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [25]),
    .d(\cu_ru/mtvec [25]),
    .o(_al_u7246_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7247 (
    .a(_al_u7244_o),
    .b(_al_u7245_o),
    .c(_al_u7246_o),
    .o(_al_u7247_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7248 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mcycle [25]),
    .d(\cu_ru/mtval [25]),
    .o(_al_u7248_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7249 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [25]),
    .d(\cu_ru/stvec [25]),
    .o(_al_u7249_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7250 (
    .a(_al_u7247_o),
    .b(_al_u7248_o),
    .c(_al_u7249_o),
    .o(csr_data[25]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7251 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_instret_sel_lutinv ),
    .c(\cu_ru/minstret [21]),
    .d(\cu_ru/mcycle [21]),
    .o(_al_u7251_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7252 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [21]),
    .d(\cu_ru/mtval [21]),
    .o(_al_u7252_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7253 (
    .a(_al_u7251_o),
    .b(_al_u7252_o),
    .c(\cu_ru/read_stval_sel_lutinv ),
    .d(\cu_ru/stval [21]),
    .o(_al_u7253_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7254 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/minstret [21]),
    .d(\cu_ru/mscratch [21]),
    .o(_al_u7254_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7255 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/mcycle [21]),
    .d(tw),
    .o(_al_u7255_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7256 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[21]),
    .d(\cu_ru/sscratch [21]),
    .o(_al_u7256_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7257 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [21]),
    .d(\cu_ru/mcause [21]),
    .o(_al_u7257_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7258 (
    .a(_al_u7254_o),
    .b(_al_u7255_o),
    .c(_al_u7256_o),
    .d(_al_u7257_o),
    .o(_al_u7258_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7259 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [21]),
    .d(\cu_ru/mtvec [21]),
    .o(_al_u7259_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7260 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(mtime_pad[21]),
    .d(\cu_ru/stvec [21]),
    .o(_al_u7260_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7261 (
    .a(_al_u7253_o),
    .b(_al_u7258_o),
    .c(_al_u7259_o),
    .d(_al_u7260_o),
    .o(csr_data[21]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7262 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [15]),
    .d(\cu_ru/mcause [15]),
    .o(_al_u7262_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7263 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[15]),
    .d(\cu_ru/mtval [15]),
    .o(_al_u7263_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7264 (
    .a(_al_u7262_o),
    .b(_al_u7263_o),
    .c(\cu_ru/read_mepc_sel_lutinv ),
    .d(\cu_ru/mepc [15]),
    .o(_al_u7264_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7265 (
    .a(_al_u6758_o),
    .b(_al_u6791_o),
    .o(\cu_ru/read_medeleg_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7266 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_medeleg_sel_lutinv ),
    .c(\cu_ru/mcycle [15]),
    .d(\cu_ru/medeleg [15]),
    .o(_al_u7266_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7267 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/minstret [15]),
    .d(\cu_ru/mscratch [15]),
    .o(_al_u7267_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7268 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[15]),
    .d(\cu_ru/minstret [15]),
    .o(_al_u7268_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7269 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [15]),
    .d(\cu_ru/sscratch [15]),
    .o(_al_u7269_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7270 (
    .a(_al_u7266_o),
    .b(_al_u7267_o),
    .c(_al_u7268_o),
    .d(_al_u7269_o),
    .o(_al_u7270_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7271 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [15]),
    .d(\cu_ru/mtvec [15]),
    .o(_al_u7271_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7272 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stval [15]),
    .d(\cu_ru/stvec [15]),
    .o(_al_u7272_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7273 (
    .a(_al_u7264_o),
    .b(_al_u7270_o),
    .c(_al_u7271_o),
    .d(_al_u7272_o),
    .o(csr_data[15]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7274 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [13]),
    .d(\cu_ru/sscratch [13]),
    .o(_al_u7274_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7275 (
    .a(_al_u6788_o),
    .b(_al_u7274_o),
    .c(\cu_ru/mcycle [13]),
    .o(_al_u7275_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7276 (
    .a(\cu_ru/read_medeleg_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[13]),
    .d(\cu_ru/medeleg [13]),
    .o(_al_u7276_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7277 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcause [13]),
    .d(\cu_ru/mscratch [13]),
    .o(_al_u7277_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7278 (
    .a(_al_u7275_o),
    .b(_al_u7276_o),
    .c(_al_u7277_o),
    .o(_al_u7278_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7279 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/minstret [13]),
    .d(\cu_ru/mepc [13]),
    .o(_al_u7279_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7280 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mtval [13]),
    .d(\cu_ru/stvec [13]),
    .o(_al_u7280_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7281 (
    .a(_al_u7278_o),
    .b(_al_u7279_o),
    .c(_al_u7280_o),
    .o(_al_u7281_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7282 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(mtime_pad[13]),
    .d(\cu_ru/sepc [13]),
    .o(_al_u7282_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7283 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [13]),
    .d(\cu_ru/mtvec [13]),
    .o(_al_u7283_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7284 (
    .a(_al_u7281_o),
    .b(_al_u7282_o),
    .c(_al_u7283_o),
    .o(csr_data[13]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u7285 (
    .a(_al_u7240_o),
    .b(id_ins[22]),
    .c(id_ins[21]),
    .d(id_ins[20]),
    .o(_al_u7285_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7286 (
    .a(_al_u7238_o),
    .b(_al_u7285_o),
    .o(\cu_ru/n84 [10]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u7287 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/n84 [10]),
    .c(\cu_ru/scause [10]),
    .o(_al_u7287_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7288 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[10]),
    .d(\cu_ru/mtvec [10]),
    .o(_al_u7288_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7289 (
    .a(_al_u7287_o),
    .b(_al_u7288_o),
    .c(\cu_ru/read_stvec_sel_lutinv ),
    .d(\cu_ru/stvec [10]),
    .o(_al_u7289_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7290 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/minstret [10]),
    .d(\cu_ru/mscratch [10]),
    .o(_al_u7290_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7291 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcycle [10]),
    .d(\cu_ru/mcause [10]),
    .o(_al_u7291_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7292 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_minstret_sel_lutinv ),
    .c(\cu_ru/minstret [10]),
    .d(\cu_ru/mcycle [10]),
    .o(_al_u7292_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7293 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[10]),
    .d(\cu_ru/sscratch [10]),
    .o(_al_u7293_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7294 (
    .a(_al_u7290_o),
    .b(_al_u7291_o),
    .c(_al_u7292_o),
    .d(_al_u7293_o),
    .o(_al_u7294_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7295 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [10]),
    .d(\cu_ru/mtval [10]),
    .o(_al_u7295_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7296 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [10]),
    .d(\cu_ru/stval [10]),
    .o(_al_u7296_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7297 (
    .a(_al_u7289_o),
    .b(_al_u7294_o),
    .c(_al_u7295_o),
    .d(_al_u7296_o),
    .o(csr_data[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7298 (
    .a(id_ill_ins),
    .b(id_ins[9]),
    .o(\ins_dec/n342 [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7299 (
    .a(id_ill_ins),
    .b(id_ins[8]),
    .o(\ins_dec/n342 [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7300 (
    .a(id_ill_ins),
    .b(id_ins[7]),
    .o(\ins_dec/n342 [7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u7301 (
    .a(id_ill_ins),
    .b(_al_u2940_o),
    .c(_al_u2941_o),
    .o(\ins_dec/n342 [6]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u7302 (
    .a(id_ill_ins),
    .b(_al_u2942_o),
    .c(_al_u2943_o),
    .o(\ins_dec/n342 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7303 (
    .a(id_ill_ins),
    .b(_al_u3924_o),
    .o(\ins_dec/n342 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7304 (
    .a(id_ill_ins),
    .b(id_ins[31]),
    .o(\ins_dec/n342 [31]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7305 (
    .a(id_ill_ins),
    .b(id_ins[30]),
    .o(\ins_dec/n342 [30]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7306 (
    .a(id_ill_ins),
    .b(_al_u3928_o),
    .o(\ins_dec/n342 [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7307 (
    .a(id_ill_ins),
    .b(id_ins[29]),
    .o(\ins_dec/n342 [29]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7308 (
    .a(id_ill_ins),
    .b(id_ins[28]),
    .o(\ins_dec/n342 [28]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7309 (
    .a(id_ill_ins),
    .b(id_ins[27]),
    .o(\ins_dec/n342 [27]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7310 (
    .a(id_ill_ins),
    .b(id_ins[26]),
    .o(\ins_dec/n342 [26]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7311 (
    .a(id_ill_ins),
    .b(id_ins[25]),
    .o(\ins_dec/n342 [25]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7312 (
    .a(id_ill_ins),
    .b(id_ins[24]),
    .o(\ins_dec/n342 [24]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7313 (
    .a(id_ill_ins),
    .b(id_ins[23]),
    .o(\ins_dec/n342 [23]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7314 (
    .a(id_ill_ins),
    .b(id_ins[22]),
    .o(\ins_dec/n342 [22]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7315 (
    .a(id_ill_ins),
    .b(id_ins[21]),
    .o(\ins_dec/n342 [21]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7316 (
    .a(id_ill_ins),
    .b(id_ins[20]),
    .o(\ins_dec/n342 [20]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7317 (
    .a(id_ill_ins),
    .b(_al_u2939_o),
    .o(\ins_dec/n342 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7318 (
    .a(id_ill_ins),
    .b(id_ins[19]),
    .o(\ins_dec/n342 [19]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7319 (
    .a(id_ill_ins),
    .b(id_ins[18]),
    .o(\ins_dec/n342 [18]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7320 (
    .a(id_ill_ins),
    .b(id_ins[17]),
    .o(\ins_dec/n342 [17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7321 (
    .a(id_ill_ins),
    .b(id_ins[16]),
    .o(\ins_dec/n342 [16]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7322 (
    .a(id_ill_ins),
    .b(id_ins[15]),
    .o(\ins_dec/n342 [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7323 (
    .a(id_ill_ins),
    .b(_al_u3216_o),
    .o(\ins_dec/n342 [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7324 (
    .a(id_ill_ins),
    .b(_al_u3217_o),
    .o(\ins_dec/n342 [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7325 (
    .a(id_ill_ins),
    .b(_al_u3384_o),
    .o(\ins_dec/n342 [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7326 (
    .a(id_ill_ins),
    .b(id_ins[11]),
    .o(\ins_dec/n342 [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7327 (
    .a(id_ill_ins),
    .b(id_ins[10]),
    .o(\ins_dec/n342 [10]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u7328 (
    .a(id_ill_ins),
    .b(_al_u2936_o),
    .c(_al_u2937_o),
    .o(\ins_dec/n342 [1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u7329 (
    .a(id_ill_ins),
    .b(_al_u2934_o),
    .c(_al_u2935_o),
    .o(\ins_dec/n342 [0]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u7330 (
    .a(_al_u2707_o),
    .b(\biu/bus_unit/mmu/n45_lutinv ),
    .c(hresp_pad),
    .o(_al_u7330_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7331 (
    .a(_al_u7330_o),
    .b(\biu/bus_unit/mmu/statu [2]),
    .c(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u7331_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7332 (
    .a(\biu/bus_unit/mmu/n39 [0]),
    .b(\biu/bus_unit/mmu_hwdata [6]),
    .o(\biu/bus_unit/mmu/n40 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'ha8ac))
    _al_u7333 (
    .a(_al_u7203_o),
    .b(_al_u7331_o),
    .c(_al_u2915_o),
    .d(\biu/bus_unit/mmu/n40 [2]),
    .o(_al_u7333_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u7334 (
    .a(_al_u7333_o),
    .b(_al_u2963_o),
    .o(\biu/bus_unit/mmu/n56 [2]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u7335 (
    .a(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .b(\cu_ru/mcause [1]),
    .c(data_csr[1]),
    .o(_al_u7335_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u7336 (
    .a(_al_u7335_o),
    .b(\cu_ru/trap_cause [1]),
    .c(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_cause/n7 [1]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u7337 (
    .a(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .b(\cu_ru/scause [1]),
    .c(data_csr[1]),
    .o(_al_u7337_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u7338 (
    .a(\cu_ru/trap_cause [1]),
    .b(_al_u5157_o),
    .c(_al_u7337_o),
    .o(\cu_ru/m_s_cause/n5 [1]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u7339 (
    .a(\cu_ru/n82 [14]),
    .b(\cu_ru/read_cycle_sel_lutinv ),
    .c(\cu_ru/mcycle [6]),
    .o(_al_u7339_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7340 (
    .a(_al_u7339_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [6]),
    .o(_al_u7340_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7341 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_medeleg_sel_lutinv ),
    .c(\cu_ru/sscratch [6]),
    .d(\cu_ru/medeleg [6]),
    .o(_al_u7341_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7342 (
    .a(_al_u7341_o),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mscratch [6]),
    .o(_al_u7342_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7343 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[6]),
    .d(\cu_ru/mcause [6]),
    .o(_al_u7343_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7344 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/mcycle [6]),
    .d(\cu_ru/scause [6]),
    .o(_al_u7344_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7345 (
    .a(_al_u7340_o),
    .b(_al_u7342_o),
    .c(_al_u7343_o),
    .d(_al_u7344_o),
    .o(_al_u7345_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7346 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [6]),
    .d(\cu_ru/mtval [6]),
    .o(_al_u7346_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7347 (
    .a(_al_u7346_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stvec [6]),
    .o(_al_u7347_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7348 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mtvec_sel_lutinv ),
    .c(\cu_ru/minstret [6]),
    .d(\cu_ru/mtvec [6]),
    .o(_al_u7348_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7349 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(mtime_pad[6]),
    .d(\cu_ru/sepc [6]),
    .o(_al_u7349_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7350 (
    .a(_al_u7345_o),
    .b(_al_u7347_o),
    .c(_al_u7348_o),
    .d(_al_u7349_o),
    .o(csr_data[6]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7351 (
    .a(csr_data[59]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[59]),
    .o(_al_u7351_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7352 (
    .a(_al_u7351_o),
    .b(rs1_data[59]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7352_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7353 (
    .a(\ins_dec/op_lui_lutinv ),
    .b(id_ins[31]),
    .o(_al_u7353_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7354 (
    .a(_al_u7352_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [59]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7355 (
    .a(csr_data[58]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[58]),
    .o(_al_u7355_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7356 (
    .a(_al_u7355_o),
    .b(rs1_data[58]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7356_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7357 (
    .a(_al_u7356_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [58]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7358 (
    .a(csr_data[57]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[57]),
    .o(_al_u7358_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7359 (
    .a(_al_u7358_o),
    .b(rs1_data[57]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7359_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7360 (
    .a(_al_u7359_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [57]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7361 (
    .a(csr_data[56]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[56]),
    .o(_al_u7361_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7362 (
    .a(_al_u7361_o),
    .b(rs1_data[56]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7362_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7363 (
    .a(_al_u7362_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [56]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7364 (
    .a(csr_data[55]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[55]),
    .o(_al_u7364_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7365 (
    .a(_al_u7364_o),
    .b(rs1_data[55]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7365_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7366 (
    .a(_al_u7365_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [55]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7367 (
    .a(csr_data[54]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[54]),
    .o(_al_u7367_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7368 (
    .a(_al_u7367_o),
    .b(rs1_data[54]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7368_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7369 (
    .a(_al_u7368_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [54]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7370 (
    .a(csr_data[53]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[53]),
    .o(_al_u7370_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7371 (
    .a(_al_u7370_o),
    .b(rs1_data[53]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7371_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7372 (
    .a(_al_u7371_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [53]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7373 (
    .a(csr_data[52]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[52]),
    .o(_al_u7373_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7374 (
    .a(_al_u7373_o),
    .b(rs1_data[52]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7374_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7375 (
    .a(_al_u7374_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [52]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7376 (
    .a(csr_data[51]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[51]),
    .o(_al_u7376_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7377 (
    .a(_al_u7376_o),
    .b(rs1_data[51]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7377_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7378 (
    .a(_al_u7377_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [51]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7379 (
    .a(csr_data[50]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[50]),
    .o(_al_u7379_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7380 (
    .a(_al_u7379_o),
    .b(rs1_data[50]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7380_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7381 (
    .a(_al_u7380_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [50]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7382 (
    .a(csr_data[49]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[49]),
    .o(_al_u7382_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7383 (
    .a(_al_u7382_o),
    .b(rs1_data[49]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7383_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7384 (
    .a(_al_u7383_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [49]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7385 (
    .a(csr_data[48]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[48]),
    .o(_al_u7385_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7386 (
    .a(_al_u7385_o),
    .b(rs1_data[48]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7386_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7387 (
    .a(_al_u7386_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [48]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7388 (
    .a(csr_data[47]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[47]),
    .o(_al_u7388_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7389 (
    .a(_al_u7388_o),
    .b(rs1_data[47]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7389_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7390 (
    .a(_al_u7389_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [47]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7391 (
    .a(csr_data[46]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[46]),
    .o(_al_u7391_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7392 (
    .a(_al_u7391_o),
    .b(rs1_data[46]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7392_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7393 (
    .a(_al_u7392_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [46]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7394 (
    .a(csr_data[45]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[45]),
    .o(_al_u7394_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7395 (
    .a(_al_u7394_o),
    .b(rs1_data[45]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7395_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7396 (
    .a(_al_u7395_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [45]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7397 (
    .a(csr_data[44]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[44]),
    .o(_al_u7397_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7398 (
    .a(_al_u7397_o),
    .b(rs1_data[44]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7398_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7399 (
    .a(_al_u7398_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [44]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7400 (
    .a(_al_u6777_o),
    .b(_al_u3397_o),
    .o(\cu_ru/n64 [32]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u7401 (
    .a(\cu_ru/n64 [32]),
    .b(\cu_ru/n90 [32]),
    .o(_al_u7401_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7402 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [33]),
    .d(\cu_ru/sscratch [33]),
    .o(_al_u7402_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7403 (
    .a(_al_u7401_o),
    .b(_al_u7402_o),
    .c(\cu_ru/read_scause_sel_lutinv ),
    .d(\cu_ru/scause [33]),
    .o(_al_u7403_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7404 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[33]),
    .d(\cu_ru/mcycle [33]),
    .o(_al_u7404_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7405 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [33]),
    .d(\cu_ru/mscratch [33]),
    .o(_al_u7405_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7406 (
    .a(_al_u7403_o),
    .b(_al_u7404_o),
    .c(_al_u7405_o),
    .o(_al_u7406_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u7407 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[33]),
    .d(\cu_ru/minstret [33]),
    .o(_al_u7407_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7408 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [33]),
    .d(\cu_ru/mtval [33]),
    .o(_al_u7408_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7409 (
    .a(_al_u7406_o),
    .b(_al_u7407_o),
    .c(_al_u7408_o),
    .o(_al_u7409_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7410 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [33]),
    .d(\cu_ru/stval [33]),
    .o(_al_u7410_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7411 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stvec [33]),
    .d(\cu_ru/mtvec [33]),
    .o(_al_u7411_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7412 (
    .a(_al_u7409_o),
    .b(_al_u7410_o),
    .c(_al_u7411_o),
    .o(csr_data[33]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7413 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [32]),
    .d(\cu_ru/sscratch [32]),
    .o(_al_u7413_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7414 (
    .a(_al_u7401_o),
    .b(_al_u7413_o),
    .c(\cu_ru/read_mcycle_sel_lutinv ),
    .d(\cu_ru/mcycle [32]),
    .o(_al_u7414_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7415 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcause [32]),
    .d(\cu_ru/mscratch [32]),
    .o(_al_u7415_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7416 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[32]),
    .d(\cu_ru/mcycle [32]),
    .o(_al_u7416_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7417 (
    .a(_al_u7414_o),
    .b(_al_u7415_o),
    .c(_al_u7416_o),
    .o(_al_u7417_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7418 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/minstret [32]),
    .d(\cu_ru/mtval [32]),
    .o(_al_u7418_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7419 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(mtime_pad[32]),
    .d(\cu_ru/mepc [32]),
    .o(_al_u7419_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7420 (
    .a(_al_u7417_o),
    .b(_al_u7418_o),
    .c(_al_u7419_o),
    .o(_al_u7420_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7421 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [32]),
    .d(\cu_ru/mtvec [32]),
    .o(_al_u7421_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7422 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stval [32]),
    .d(\cu_ru/stvec [32]),
    .o(_al_u7422_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*B*A)"),
    .INIT(8'h7f))
    _al_u7423 (
    .a(_al_u7420_o),
    .b(_al_u7421_o),
    .c(_al_u7422_o),
    .o(csr_data[32]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7424 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[30]),
    .d(\cu_ru/mcycle [30]),
    .o(_al_u7424_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7425 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [30]),
    .d(\cu_ru/sscratch [30]),
    .o(_al_u7425_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7426 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [30]),
    .d(\cu_ru/mtvec [30]),
    .o(_al_u7426_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7427 (
    .a(_al_u7424_o),
    .b(_al_u7425_o),
    .c(_al_u7426_o),
    .o(_al_u7427_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7428 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [30]),
    .d(\cu_ru/mscratch [30]),
    .o(_al_u7428_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7429 (
    .a(_al_u7427_o),
    .b(_al_u7428_o),
    .c(\cu_ru/read_mcause_sel_lutinv ),
    .d(\cu_ru/mcause [30]),
    .o(_al_u7429_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u7430 (
    .a(\cu_ru/n82 [14]),
    .b(\cu_ru/n84 [10]),
    .o(_al_u7430_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7431 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/minstret [30]),
    .d(\cu_ru/mtval [30]),
    .o(_al_u7431_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7432 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(mtime_pad[30]),
    .d(\cu_ru/sepc [30]),
    .o(_al_u7432_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7433 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [30]),
    .d(\cu_ru/stvec [30]),
    .o(_al_u7433_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7434 (
    .a(_al_u7430_o),
    .b(_al_u7431_o),
    .c(_al_u7432_o),
    .d(_al_u7433_o),
    .o(_al_u7434_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7435 (
    .a(_al_u7429_o),
    .b(_al_u7434_o),
    .o(csr_data[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7436 (
    .a(_al_u7430_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [28]),
    .o(_al_u7436_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7437 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [28]),
    .d(\cu_ru/sscratch [28]),
    .o(_al_u7437_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7438 (
    .a(_al_u7437_o),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[28]),
    .o(_al_u7438_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7439 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcycle [28]),
    .d(\cu_ru/mcause [28]),
    .o(_al_u7439_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7440 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [28]),
    .d(\cu_ru/mscratch [28]),
    .o(_al_u7440_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7441 (
    .a(_al_u7436_o),
    .b(_al_u7438_o),
    .c(_al_u7439_o),
    .d(_al_u7440_o),
    .o(_al_u7441_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7442 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [28]),
    .d(\cu_ru/mtvec [28]),
    .o(_al_u7442_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7443 (
    .a(_al_u7442_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stvec [28]),
    .o(_al_u7443_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7444 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/minstret [28]),
    .d(\cu_ru/mtval [28]),
    .o(_al_u7444_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7445 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(mtime_pad[28]),
    .d(\cu_ru/mepc [28]),
    .o(_al_u7445_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7446 (
    .a(_al_u7441_o),
    .b(_al_u7443_o),
    .c(_al_u7444_o),
    .d(_al_u7445_o),
    .o(csr_data[28]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7447 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/mcycle [19]),
    .d(mxr),
    .o(_al_u7447_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7448 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/minstret [19]),
    .d(\cu_ru/mscratch [19]),
    .o(_al_u7448_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7449 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[19]),
    .d(\cu_ru/mcause [19]),
    .o(_al_u7449_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7450 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/mcycle [19]),
    .d(\cu_ru/scause [19]),
    .o(_al_u7450_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7451 (
    .a(_al_u7447_o),
    .b(_al_u7448_o),
    .c(_al_u7449_o),
    .d(_al_u7450_o),
    .o(_al_u7451_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7452 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/n64 [32]),
    .c(\cu_ru/minstret [19]),
    .d(mxr),
    .o(_al_u7452_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7453 (
    .a(_al_u7451_o),
    .b(_al_u7452_o),
    .c(\cu_ru/read_sscratch_sel_lutinv ),
    .d(\cu_ru/sscratch [19]),
    .o(_al_u7453_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7454 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/stval [19]),
    .d(\cu_ru/mtval [19]),
    .o(_al_u7454_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7455 (
    .a(_al_u7454_o),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [19]),
    .o(_al_u7455_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7456 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(mtime_pad[19]),
    .d(\cu_ru/stvec [19]),
    .o(_al_u7456_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7457 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [19]),
    .d(\cu_ru/mtvec [19]),
    .o(_al_u7457_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7458 (
    .a(_al_u7453_o),
    .b(_al_u7455_o),
    .c(_al_u7456_o),
    .d(_al_u7457_o),
    .o(csr_data[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7459 (
    .a(_al_u7430_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mtval [14]),
    .o(_al_u7459_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7460 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[14]),
    .d(\cu_ru/mcycle [14]),
    .o(_al_u7460_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7461 (
    .a(_al_u7460_o),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [14]),
    .o(_al_u7461_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7462 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mscratch [14]),
    .d(\cu_ru/sscratch [14]),
    .o(_al_u7462_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7463 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/mcycle [14]),
    .d(\cu_ru/scause [14]),
    .o(_al_u7463_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7464 (
    .a(_al_u7459_o),
    .b(_al_u7461_o),
    .c(_al_u7462_o),
    .d(_al_u7463_o),
    .o(_al_u7464_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7465 (
    .a(\cu_ru/read_sepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/sepc [14]),
    .d(\cu_ru/stvec [14]),
    .o(_al_u7465_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7466 (
    .a(_al_u7465_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [14]),
    .o(_al_u7466_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7467 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/minstret [14]),
    .d(\cu_ru/mepc [14]),
    .o(_al_u7467_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7468 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[14]),
    .d(\cu_ru/mtvec [14]),
    .o(_al_u7468_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7469 (
    .a(_al_u7464_o),
    .b(_al_u7466_o),
    .c(_al_u7467_o),
    .d(_al_u7468_o),
    .o(csr_data[14]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7470 (
    .a(\cu_ru/read_mscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[11]),
    .d(\cu_ru/mscratch [11]),
    .o(_al_u7470_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7471 (
    .a(_al_u7470_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [11]),
    .o(_al_u7471_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7472 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_minstret_sel_lutinv ),
    .c(\cu_ru/minstret [11]),
    .d(\cu_ru/mcycle [11]),
    .o(_al_u7472_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7473 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [11]),
    .d(\cu_ru/sscratch [11]),
    .o(_al_u7473_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7474 (
    .a(_al_u7471_o),
    .b(_al_u7472_o),
    .c(_al_u7473_o),
    .o(_al_u7474_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7475 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [11]),
    .d(\cu_ru/stvec [11]),
    .o(_al_u7475_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7476 (
    .a(_al_u7475_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mtval [11]),
    .o(_al_u7476_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7477 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [11]),
    .d(\cu_ru/mtvec [11]),
    .o(_al_u7477_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u7478 (
    .a(_al_u3393_o),
    .b(id_ins[22]),
    .c(id_ins[21]),
    .d(id_ins[20]),
    .o(_al_u7478_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7479 (
    .a(_al_u6766_o),
    .b(_al_u7478_o),
    .o(\cu_ru/read_mip_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7480 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_mip_sel_lutinv ),
    .c(mtime_pad[11]),
    .d(\cu_ru/m_sip [11]),
    .o(_al_u7480_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7481 (
    .a(_al_u7476_o),
    .b(_al_u7477_o),
    .c(_al_u7480_o),
    .o(_al_u7481_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7482 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/minstret [11]),
    .d(\cu_ru/scause [11]),
    .o(_al_u7482_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7483 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/mcause [11]),
    .d(\cu_ru/mstatus [11]),
    .o(_al_u7483_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7484 (
    .a(_al_u7474_o),
    .b(_al_u7481_o),
    .c(_al_u7482_o),
    .d(_al_u7483_o),
    .o(csr_data[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7485 (
    .a(_al_u7330_o),
    .b(\biu/bus_unit/mmu/statu [1]),
    .c(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u7485_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'h4e))
    _al_u7486 (
    .a(_al_u7202_o),
    .b(_al_u7485_o),
    .c(\biu/bus_unit/mmu_hwdata [6]),
    .o(_al_u7486_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7487 (
    .a(\biu/bus_unit/mmu/n37_lutinv ),
    .b(\biu/bus_unit/mmu/n39 [0]),
    .c(\biu/bus_unit/mmu_hwdata [6]),
    .o(_al_u7487_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7488 (
    .a(_al_u7486_o),
    .b(_al_u7487_o),
    .c(\biu/bus_unit/mmu_hwdata [2]),
    .o(_al_u7488_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .INIT(16'h3202))
    _al_u7489 (
    .a(_al_u7488_o),
    .b(_al_u2697_o),
    .c(_al_u2964_o),
    .d(hresp_pad),
    .o(_al_u7489_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(~C*~A))"),
    .INIT(8'hcd))
    _al_u7490 (
    .a(_al_u7489_o),
    .b(_al_u2963_o),
    .c(_al_u2698_o),
    .o(\biu/bus_unit/mmu/n56 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*A))"),
    .INIT(16'h51f3))
    _al_u7491 (
    .a(\biu/bus_unit/mmu/mux10_b0_sel_is_2_o ),
    .b(\biu/bus_unit/mmu/n45_lutinv ),
    .c(hresp_pad),
    .d(\biu/bus_unit/mmu/statu [0]),
    .o(_al_u7491_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u7492 (
    .a(_al_u7491_o),
    .b(\biu/bus_unit/mmu/statu [1]),
    .c(\biu/bus_unit/mmu/statu [3]),
    .o(_al_u7492_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u7493 (
    .a(\biu/bus_unit/mmu/n2 ),
    .b(_al_u7487_o),
    .c(_al_u2964_o),
    .o(_al_u7493_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(~B*~A)))"),
    .INIT(16'hf010))
    _al_u7494 (
    .a(_al_u7202_o),
    .b(_al_u7492_o),
    .c(_al_u7493_o),
    .d(\biu/bus_unit/mmu/n37_lutinv ),
    .o(_al_u7494_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u7495 (
    .a(_al_u2964_o),
    .b(hready_pad),
    .c(hresp_pad),
    .o(_al_u7495_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*~B)*~(~D*~A))"),
    .INIT(16'h3075))
    _al_u7496 (
    .a(_al_u7494_o),
    .b(_al_u2914_o),
    .c(_al_u2698_o),
    .d(_al_u7495_o),
    .o(\biu/bus_unit/mmu/n56 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7497 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/mcycle [7]),
    .d(\cu_ru/mstatus [7]),
    .o(_al_u7497_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7498 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mscratch [7]),
    .d(\cu_ru/sscratch [7]),
    .o(_al_u7498_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7499 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/minstret [7]),
    .d(\cu_ru/mcause [7]),
    .o(_al_u7499_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7500 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[7]),
    .d(\cu_ru/mcycle [7]),
    .o(_al_u7500_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7501 (
    .a(_al_u7497_o),
    .b(_al_u7498_o),
    .c(_al_u7499_o),
    .d(_al_u7500_o),
    .o(_al_u7501_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7502 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_medeleg_sel_lutinv ),
    .c(\cu_ru/scause [7]),
    .d(\cu_ru/medeleg [7]),
    .o(_al_u7502_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7503 (
    .a(_al_u7501_o),
    .b(_al_u7502_o),
    .c(\cu_ru/read_instret_sel_lutinv ),
    .d(\cu_ru/minstret [7]),
    .o(_al_u7503_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7504 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(mtime_pad[7]),
    .d(\cu_ru/stvec [7]),
    .o(_al_u7504_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7505 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mtval [7]),
    .d(\cu_ru/mtvec [7]),
    .o(_al_u7505_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7506 (
    .a(\cu_ru/read_sepc_sel_lutinv ),
    .b(\cu_ru/read_mip_sel_lutinv ),
    .c(\cu_ru/sepc [7]),
    .d(\cu_ru/m_sip [7]),
    .o(_al_u7506_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7507 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [7]),
    .d(\cu_ru/stval [7]),
    .o(_al_u7507_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7508 (
    .a(_al_u7504_o),
    .b(_al_u7505_o),
    .c(_al_u7506_o),
    .d(_al_u7507_o),
    .o(_al_u7508_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7509 (
    .a(_al_u7503_o),
    .b(_al_u7508_o),
    .o(csr_data[7]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7510 (
    .a(rs1_data[63]),
    .b(_al_u7141_o),
    .o(_al_u7510_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7511 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[63]),
    .o(_al_u7511_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7512 (
    .a(csr_data[63]),
    .b(_al_u7510_o),
    .c(_al_u7511_o),
    .d(id_system),
    .o(_al_u7512_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7513 (
    .a(_al_u7512_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [63]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7514 (
    .a(rs1_data[62]),
    .b(_al_u7141_o),
    .o(_al_u7514_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7515 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[62]),
    .o(_al_u7515_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7516 (
    .a(csr_data[62]),
    .b(_al_u7514_o),
    .c(_al_u7515_o),
    .d(id_system),
    .o(_al_u7516_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7517 (
    .a(_al_u7516_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [62]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7518 (
    .a(rs1_data[61]),
    .b(_al_u7141_o),
    .o(_al_u7518_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7519 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[61]),
    .o(_al_u7519_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7520 (
    .a(csr_data[61]),
    .b(_al_u7518_o),
    .c(_al_u7519_o),
    .d(id_system),
    .o(_al_u7520_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7521 (
    .a(_al_u7520_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [61]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7522 (
    .a(rs1_data[60]),
    .b(_al_u7141_o),
    .o(_al_u7522_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7523 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[60]),
    .o(_al_u7523_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7524 (
    .a(csr_data[60]),
    .b(_al_u7522_o),
    .c(_al_u7523_o),
    .d(id_system),
    .o(_al_u7524_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7525 (
    .a(_al_u7524_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [60]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7526 (
    .a(rs1_data[43]),
    .b(_al_u7141_o),
    .o(_al_u7526_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7527 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[43]),
    .o(_al_u7527_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7528 (
    .a(csr_data[43]),
    .b(_al_u7526_o),
    .c(_al_u7527_o),
    .d(id_system),
    .o(_al_u7528_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7529 (
    .a(_al_u7528_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [43]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7530 (
    .a(csr_data[42]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[42]),
    .o(_al_u7530_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7531 (
    .a(rs1_data[42]),
    .b(_al_u7141_o),
    .o(_al_u7531_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7532 (
    .a(_al_u7530_o),
    .b(_al_u7531_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[31]),
    .o(\ins_dec/n272 [42]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7533 (
    .a(rs1_data[41]),
    .b(_al_u7141_o),
    .o(_al_u7533_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7534 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[41]),
    .o(_al_u7534_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7535 (
    .a(csr_data[41]),
    .b(_al_u7533_o),
    .c(_al_u7534_o),
    .d(id_system),
    .o(_al_u7535_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7536 (
    .a(_al_u7535_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [41]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7537 (
    .a(rs1_data[40]),
    .b(_al_u7141_o),
    .o(_al_u7537_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7538 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[40]),
    .o(_al_u7538_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7539 (
    .a(csr_data[40]),
    .b(_al_u7537_o),
    .c(_al_u7538_o),
    .d(id_system),
    .o(_al_u7539_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7540 (
    .a(_al_u7539_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [40]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7541 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/minstret [4]),
    .d(\cu_ru/mcause [4]),
    .o(_al_u7541_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7542 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/mcycle [4]),
    .d(\cu_ru/scause [4]),
    .o(_al_u7542_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7543 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[4]),
    .d(\cu_ru/mcycle [4]),
    .o(_al_u7543_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7544 (
    .a(_al_u7430_o),
    .b(_al_u7541_o),
    .c(_al_u7542_o),
    .d(_al_u7543_o),
    .o(_al_u7544_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7545 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [4]),
    .d(\cu_ru/mtvec [4]),
    .o(_al_u7545_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7546 (
    .a(_al_u7545_o),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [4]),
    .o(_al_u7546_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7547 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(mtime_pad[4]),
    .d(\cu_ru/sepc [4]),
    .o(_al_u7547_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7548 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mtval [4]),
    .d(\cu_ru/stvec [4]),
    .o(_al_u7548_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7549 (
    .a(_al_u7546_o),
    .b(_al_u7547_o),
    .c(_al_u7548_o),
    .o(_al_u7549_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7550 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/minstret [4]),
    .d(\cu_ru/mscratch [4]),
    .o(_al_u7550_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7551 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_medeleg_sel_lutinv ),
    .c(\cu_ru/sscratch [4]),
    .d(\cu_ru/medeleg [4]),
    .o(_al_u7551_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7552 (
    .a(_al_u7544_o),
    .b(_al_u7549_o),
    .c(_al_u7550_o),
    .d(_al_u7551_o),
    .o(csr_data[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7553 (
    .a(rs1_data[39]),
    .b(_al_u7141_o),
    .o(_al_u7553_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7554 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[39]),
    .o(_al_u7554_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7555 (
    .a(csr_data[39]),
    .b(_al_u7553_o),
    .c(_al_u7554_o),
    .d(id_system),
    .o(_al_u7555_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7556 (
    .a(_al_u7555_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [39]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7557 (
    .a(rs1_data[38]),
    .b(_al_u7141_o),
    .o(_al_u7557_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7558 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[38]),
    .o(_al_u7558_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7559 (
    .a(csr_data[38]),
    .b(_al_u7557_o),
    .c(_al_u7558_o),
    .d(id_system),
    .o(_al_u7559_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7560 (
    .a(_al_u7559_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [38]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7561 (
    .a(rs1_data[37]),
    .b(_al_u7141_o),
    .o(_al_u7561_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7562 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[37]),
    .o(_al_u7562_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7563 (
    .a(csr_data[37]),
    .b(_al_u7561_o),
    .c(_al_u7562_o),
    .d(id_system),
    .o(_al_u7563_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7564 (
    .a(_al_u7563_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [37]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7565 (
    .a(rs1_data[36]),
    .b(_al_u7141_o),
    .o(_al_u7565_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7566 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[36]),
    .o(_al_u7566_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7567 (
    .a(csr_data[36]),
    .b(_al_u7565_o),
    .c(_al_u7566_o),
    .d(id_system),
    .o(_al_u7567_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7568 (
    .a(_al_u7567_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [36]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7569 (
    .a(rs1_data[31]),
    .b(_al_u7141_o),
    .o(_al_u7569_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7570 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[31]),
    .o(_al_u7570_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7571 (
    .a(csr_data[31]),
    .b(_al_u7569_o),
    .c(_al_u7570_o),
    .d(id_system),
    .o(_al_u7571_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7572 (
    .a(_al_u7571_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7573 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/scause [3]),
    .d(\cu_ru/mie ),
    .o(_al_u7573_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7574 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[3]),
    .d(\cu_ru/sscratch [3]),
    .o(_al_u7574_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7575 (
    .a(\cu_ru/read_sepc_sel_lutinv ),
    .b(\cu_ru/read_mip_sel_lutinv ),
    .c(\cu_ru/sepc [3]),
    .d(\cu_ru/m_sip [3]),
    .o(_al_u7575_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7576 (
    .a(_al_u7573_o),
    .b(_al_u7574_o),
    .c(_al_u7575_o),
    .o(_al_u7576_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7577 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcause [3]),
    .d(\cu_ru/mscratch [3]),
    .o(_al_u7577_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7578 (
    .a(_al_u7576_o),
    .b(_al_u7577_o),
    .c(\cu_ru/read_medeleg_sel_lutinv ),
    .d(\cu_ru/medeleg [3]),
    .o(_al_u7578_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u7579 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[3]),
    .d(\cu_ru/minstret [3]),
    .o(_al_u7579_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7580 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mcycle [3]),
    .d(\cu_ru/mtval [3]),
    .o(_al_u7580_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7581 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [3]),
    .d(\cu_ru/stvec [3]),
    .o(_al_u7581_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7582 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [3]),
    .d(\cu_ru/mtvec [3]),
    .o(_al_u7582_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7583 (
    .a(_al_u7579_o),
    .b(_al_u7580_o),
    .c(_al_u7581_o),
    .d(_al_u7582_o),
    .o(_al_u7583_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7584 (
    .a(_al_u7578_o),
    .b(_al_u7583_o),
    .o(csr_data[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7585 (
    .a(csr_data[29]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[29]),
    .o(_al_u7585_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7586 (
    .a(rs1_data[29]),
    .b(_al_u7141_o),
    .o(_al_u7586_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7587 (
    .a(_al_u7585_o),
    .b(_al_u7586_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[29]),
    .o(\ins_dec/n272 [29]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7588 (
    .a(csr_data[27]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[27]),
    .o(_al_u7588_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7589 (
    .a(rs1_data[27]),
    .b(_al_u7141_o),
    .o(_al_u7589_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7590 (
    .a(_al_u7588_o),
    .b(_al_u7589_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[27]),
    .o(\ins_dec/n272 [27]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7591 (
    .a(csr_data[26]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[26]),
    .o(_al_u7591_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7592 (
    .a(rs1_data[26]),
    .b(_al_u7141_o),
    .o(_al_u7592_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7593 (
    .a(_al_u7591_o),
    .b(_al_u7592_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[26]),
    .o(\ins_dec/n272 [26]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7594 (
    .a(csr_data[24]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[24]),
    .o(_al_u7594_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7595 (
    .a(rs1_data[24]),
    .b(_al_u7141_o),
    .o(_al_u7595_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7596 (
    .a(_al_u7594_o),
    .b(_al_u7595_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[24]),
    .o(\ins_dec/n272 [24]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7597 (
    .a(csr_data[23]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[23]),
    .o(_al_u7597_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7598 (
    .a(rs1_data[23]),
    .b(_al_u7141_o),
    .o(_al_u7598_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7599 (
    .a(_al_u7597_o),
    .b(_al_u7598_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[23]),
    .o(\ins_dec/n272 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7600 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcycle [22]),
    .d(\cu_ru/mcause [22]),
    .o(_al_u7600_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7601 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[22]),
    .d(\cu_ru/scause [22]),
    .o(_al_u7601_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7602 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/minstret [22]),
    .d(tsr),
    .o(_al_u7602_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7603 (
    .a(_al_u7430_o),
    .b(_al_u7600_o),
    .c(_al_u7601_o),
    .d(_al_u7602_o),
    .o(_al_u7603_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7604 (
    .a(\cu_ru/read_mepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mepc [22]),
    .d(\cu_ru/stvec [22]),
    .o(_al_u7604_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7605 (
    .a(_al_u7604_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[22]),
    .o(_al_u7605_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7606 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/stval [22]),
    .d(\cu_ru/mtval [22]),
    .o(_al_u7606_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7607 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [22]),
    .d(\cu_ru/mtvec [22]),
    .o(_al_u7607_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7608 (
    .a(_al_u7605_o),
    .b(_al_u7606_o),
    .c(_al_u7607_o),
    .o(_al_u7608_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7609 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/minstret [22]),
    .d(\cu_ru/mscratch [22]),
    .o(_al_u7609_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7610 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [22]),
    .d(\cu_ru/sscratch [22]),
    .o(_al_u7610_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7611 (
    .a(_al_u7603_o),
    .b(_al_u7608_o),
    .c(_al_u7609_o),
    .d(_al_u7610_o),
    .o(csr_data[22]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7612 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[20]),
    .d(\cu_ru/mcause [20]),
    .o(_al_u7612_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7613 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/minstret [20]),
    .d(\cu_ru/sscratch [20]),
    .o(_al_u7613_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7614 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/mcycle [20]),
    .d(\cu_ru/scause [20]),
    .o(_al_u7614_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7615 (
    .a(_al_u7430_o),
    .b(_al_u7612_o),
    .c(_al_u7613_o),
    .d(_al_u7614_o),
    .o(_al_u7615_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7616 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(mtime_pad[20]),
    .d(\cu_ru/stvec [20]),
    .o(_al_u7616_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7617 (
    .a(_al_u7616_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [20]),
    .o(_al_u7617_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7618 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [20]),
    .d(\cu_ru/mtvec [20]),
    .o(_al_u7618_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7619 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/stval [20]),
    .d(\cu_ru/mtval [20]),
    .o(_al_u7619_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7620 (
    .a(_al_u7617_o),
    .b(_al_u7618_o),
    .c(_al_u7619_o),
    .o(_al_u7620_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7621 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/minstret [20]),
    .d(tvm),
    .o(_al_u7621_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7622 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [20]),
    .d(\cu_ru/mscratch [20]),
    .o(_al_u7622_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7623 (
    .a(_al_u7615_o),
    .b(_al_u7620_o),
    .c(_al_u7621_o),
    .d(_al_u7622_o),
    .o(csr_data[20]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u7624 (
    .a(\cu_ru/n82 [14]),
    .b(\cu_ru/n64 [32]),
    .c(sum),
    .o(_al_u7624_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7625 (
    .a(_al_u7624_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stvec [18]),
    .o(_al_u7625_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7626 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcycle [18]),
    .d(\cu_ru/mcause [18]),
    .o(_al_u7626_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7627 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [18]),
    .d(\cu_ru/mscratch [18]),
    .o(_al_u7627_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7628 (
    .a(_al_u7625_o),
    .b(_al_u7626_o),
    .c(_al_u7627_o),
    .o(_al_u7628_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7629 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[18]),
    .d(\cu_ru/stval [18]),
    .o(_al_u7629_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7630 (
    .a(_al_u7629_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mtval [18]),
    .o(_al_u7630_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7631 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/minstret [18]),
    .d(\cu_ru/sepc [18]),
    .o(_al_u7631_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7632 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [18]),
    .d(\cu_ru/mtvec [18]),
    .o(_al_u7632_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7633 (
    .a(_al_u7630_o),
    .b(_al_u7631_o),
    .c(_al_u7632_o),
    .o(_al_u7633_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7634 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/sscratch [18]),
    .d(sum),
    .o(_al_u7634_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7635 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[18]),
    .d(\cu_ru/scause [18]),
    .o(_al_u7635_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7636 (
    .a(_al_u7628_o),
    .b(_al_u7633_o),
    .c(_al_u7634_o),
    .d(_al_u7635_o),
    .o(csr_data[18]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7637 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/minstret [17]),
    .d(mprv),
    .o(_al_u7637_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7638 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcause [17]),
    .d(\cu_ru/mscratch [17]),
    .o(_al_u7638_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7639 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_minstret_sel_lutinv ),
    .c(\cu_ru/minstret [17]),
    .d(\cu_ru/mcycle [17]),
    .o(_al_u7639_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7640 (
    .a(_al_u7430_o),
    .b(_al_u7637_o),
    .c(_al_u7638_o),
    .d(_al_u7639_o),
    .o(_al_u7640_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7641 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/stval [17]),
    .d(\cu_ru/mtval [17]),
    .o(_al_u7641_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7642 (
    .a(_al_u7641_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[17]),
    .o(_al_u7642_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7643 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [17]),
    .d(\cu_ru/mtvec [17]),
    .o(_al_u7643_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7644 (
    .a(\cu_ru/read_sepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/sepc [17]),
    .d(\cu_ru/stvec [17]),
    .o(_al_u7644_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7645 (
    .a(_al_u7642_o),
    .b(_al_u7643_o),
    .c(_al_u7644_o),
    .o(_al_u7645_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7646 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [17]),
    .d(\cu_ru/sscratch [17]),
    .o(_al_u7646_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7647 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[17]),
    .d(\cu_ru/scause [17]),
    .o(_al_u7647_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7648 (
    .a(_al_u7640_o),
    .b(_al_u7645_o),
    .c(_al_u7646_o),
    .d(_al_u7647_o),
    .o(csr_data[17]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7649 (
    .a(csr_data[16]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[16]),
    .o(_al_u7649_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7650 (
    .a(rs1_data[16]),
    .b(_al_u7141_o),
    .o(_al_u7650_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7651 (
    .a(_al_u7649_o),
    .b(_al_u7650_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[16]),
    .o(\ins_dec/n272 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7652 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/n90 [32]),
    .c(\cu_ru/sscratch [12]),
    .d(\cu_ru/mstatus [12]),
    .o(_al_u7652_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u7653 (
    .a(_al_u7652_o),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/n84 [10]),
    .d(\cu_ru/mcause [12]),
    .o(_al_u7653_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7654 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[12]),
    .d(\cu_ru/mcycle [12]),
    .o(_al_u7654_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7655 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/mcycle [12]),
    .d(\cu_ru/scause [12]),
    .o(_al_u7655_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7656 (
    .a(_al_u7653_o),
    .b(_al_u7654_o),
    .c(_al_u7655_o),
    .o(_al_u7656_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7657 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mtval [12]),
    .d(\cu_ru/stvec [12]),
    .o(_al_u7657_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7658 (
    .a(_al_u7657_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/stval [12]),
    .o(_al_u7658_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7659 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [12]),
    .d(\cu_ru/mtvec [12]),
    .o(_al_u7659_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7660 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(mtime_pad[12]),
    .d(\cu_ru/sepc [12]),
    .o(_al_u7660_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7661 (
    .a(_al_u7658_o),
    .b(_al_u7659_o),
    .c(_al_u7660_o),
    .o(_al_u7661_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7662 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/read_medeleg_sel_lutinv ),
    .c(\cu_ru/minstret [12]),
    .d(\cu_ru/medeleg [12]),
    .o(_al_u7662_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7663 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/minstret [12]),
    .d(\cu_ru/mscratch [12]),
    .o(_al_u7663_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7664 (
    .a(_al_u7656_o),
    .b(_al_u7661_o),
    .c(_al_u7662_o),
    .d(_al_u7663_o),
    .o(csr_data[12]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u7665 (
    .a(\cu_ru/n82 [14]),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/sscratch [8]),
    .o(_al_u7665_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7666 (
    .a(_al_u7665_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [8]),
    .o(_al_u7666_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7667 (
    .a(\cu_ru/read_scause_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/scause [8]),
    .d(\cu_ru/mscratch [8]),
    .o(_al_u7667_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7668 (
    .a(_al_u7667_o),
    .b(\cu_ru/read_instret_sel_lutinv ),
    .c(\cu_ru/minstret [8]),
    .o(_al_u7668_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7669 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[8]),
    .d(\cu_ru/minstret [8]),
    .o(_al_u7669_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7670 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_medeleg_sel_lutinv ),
    .c(\cu_ru/mcause [8]),
    .d(\cu_ru/medeleg [8]),
    .o(_al_u7670_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7671 (
    .a(_al_u7666_o),
    .b(_al_u7668_o),
    .c(_al_u7669_o),
    .d(_al_u7670_o),
    .o(_al_u7671_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7672 (
    .a(_al_u7401_o),
    .b(\cu_ru/read_mtval_sel_lutinv ),
    .c(\cu_ru/mstatus [8]),
    .d(\cu_ru/mtval [8]),
    .o(_al_u7672_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7673 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/mcycle [8]),
    .d(\cu_ru/stval [8]),
    .o(_al_u7673_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7674 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(mtime_pad[8]),
    .d(\cu_ru/stvec [8]),
    .o(_al_u7674_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7675 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [8]),
    .d(\cu_ru/mtvec [8]),
    .o(_al_u7675_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7676 (
    .a(_al_u7672_o),
    .b(_al_u7673_o),
    .c(_al_u7674_o),
    .d(_al_u7675_o),
    .o(_al_u7676_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7677 (
    .a(_al_u7671_o),
    .b(_al_u7676_o),
    .o(csr_data[8]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7678 (
    .a(csr_data[35]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[35]),
    .o(_al_u7678_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    _al_u7679 (
    .a(_al_u7678_o),
    .b(rs1_data[35]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7679_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u7680 (
    .a(_al_u7679_o),
    .b(_al_u7353_o),
    .o(\ins_dec/n272 [35]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7681 (
    .a(rs1_data[34]),
    .b(_al_u7141_o),
    .o(_al_u7681_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7682 (
    .a(_al_u7141_o),
    .b(id_system),
    .c(id_ins_pc[34]),
    .o(_al_u7682_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*~A)))"),
    .INIT(16'h1303))
    _al_u7683 (
    .a(csr_data[34]),
    .b(_al_u7681_o),
    .c(_al_u7682_o),
    .d(id_system),
    .o(_al_u7683_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u7684 (
    .a(_al_u7683_o),
    .b(\ins_dec/op_lui_lutinv ),
    .c(id_ins[31]),
    .o(\ins_dec/n272 [34]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7685 (
    .a(csr_data[25]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[25]),
    .o(_al_u7685_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7686 (
    .a(rs1_data[25]),
    .b(_al_u7141_o),
    .o(_al_u7686_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7687 (
    .a(_al_u7685_o),
    .b(_al_u7686_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[25]),
    .o(\ins_dec/n272 [25]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7688 (
    .a(rs1_data[21]),
    .b(_al_u7141_o),
    .o(_al_u7688_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7689 (
    .a(csr_data[21]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[21]),
    .o(_al_u7689_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7690 (
    .a(_al_u7688_o),
    .b(_al_u7689_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[21]),
    .o(\ins_dec/n272 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7691 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_sscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [2]),
    .d(\cu_ru/sscratch [2]),
    .o(_al_u7691_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7692 (
    .a(_al_u7691_o),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[2]),
    .o(_al_u7692_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7693 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [2]),
    .d(\cu_ru/mscratch [2]),
    .o(_al_u7693_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u7694 (
    .a(_al_u7239_o),
    .b(_al_u7240_o),
    .c(id_ins[22]),
    .o(_al_u7694_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u7695 (
    .a(_al_u7693_o),
    .b(_al_u7694_o),
    .c(\cu_ru/read_medeleg_sel_lutinv ),
    .d(\cu_ru/medeleg [2]),
    .o(_al_u7695_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7696 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/scause [2]),
    .d(\cu_ru/mcause [2]),
    .o(_al_u7696_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7697 (
    .a(_al_u7430_o),
    .b(_al_u7692_o),
    .c(_al_u7695_o),
    .d(_al_u7696_o),
    .o(_al_u7697_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u7698 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[2]),
    .d(\cu_ru/minstret [2]),
    .o(_al_u7698_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7699 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [2]),
    .d(\cu_ru/mtval [2]),
    .o(_al_u7699_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7700 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stvec [2]),
    .d(\cu_ru/mtvec [2]),
    .o(_al_u7700_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7701 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [2]),
    .d(\cu_ru/stval [2]),
    .o(_al_u7701_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7702 (
    .a(_al_u7698_o),
    .b(_al_u7699_o),
    .c(_al_u7700_o),
    .d(_al_u7701_o),
    .o(_al_u7702_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u7703 (
    .a(_al_u7697_o),
    .b(_al_u7702_o),
    .o(csr_data[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7704 (
    .a(rs1_data[15]),
    .b(_al_u7141_o),
    .o(_al_u7704_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7705 (
    .a(csr_data[15]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[15]),
    .o(_al_u7705_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7706 (
    .a(_al_u7704_o),
    .b(_al_u7705_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[15]),
    .o(\ins_dec/n272 [15]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7707 (
    .a(csr_data[13]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[13]),
    .o(_al_u7707_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7708 (
    .a(rs1_data[13]),
    .b(_al_u7141_o),
    .o(_al_u7708_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7709 (
    .a(_al_u7707_o),
    .b(_al_u7708_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(_al_u3217_o),
    .o(\ins_dec/n272 [13]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7710 (
    .a(csr_data[10]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[10]),
    .o(_al_u7710_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7711 (
    .a(_al_u7710_o),
    .b(rs1_data[10]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7712 (
    .a(\cu_ru/read_instret_sel_lutinv ),
    .b(\cu_ru/read_medeleg_sel_lutinv ),
    .c(\cu_ru/minstret [0]),
    .d(\cu_ru/medeleg [0]),
    .o(_al_u7712_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7713 (
    .a(_al_u7712_o),
    .b(\cu_ru/read_mtvec_sel_lutinv ),
    .c(\cu_ru/mtvec [0]),
    .o(_al_u7713_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7714 (
    .a(_al_u6777_o),
    .b(_al_u7478_o),
    .c(\cu_ru/mstatus [1]),
    .o(\cu_ru/n66_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u7715 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/n66_lutinv ),
    .c(\cu_ru/sscratch [0]),
    .o(_al_u7715_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u7716 (
    .a(id_ins[25]),
    .b(_al_u3392_o),
    .c(\cu_ru/mcountinhibit ),
    .o(_al_u7716_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u7717 (
    .a(_al_u7716_o),
    .b(id_ins[20]),
    .c(_al_u3394_o),
    .o(_al_u7717_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(D*A)))"),
    .INIT(16'he0c0))
    _al_u7718 (
    .a(_al_u7478_o),
    .b(_al_u7717_o),
    .c(_al_u6791_o),
    .d(\cu_ru/mie ),
    .o(_al_u7718_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u7719 (
    .a(_al_u7715_o),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(_al_u7718_o),
    .d(\cu_ru/mcause [0]),
    .o(_al_u7719_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7720 (
    .a(\cu_ru/read_minstret_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/minstret [0]),
    .d(\cu_ru/scause [0]),
    .o(_al_u7720_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7721 (
    .a(\cu_ru/read_mscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[0]),
    .d(\cu_ru/mscratch [0]),
    .o(_al_u7721_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7722 (
    .a(_al_u7713_o),
    .b(_al_u7719_o),
    .c(_al_u7720_o),
    .d(_al_u7721_o),
    .o(_al_u7722_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7723 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mcycle [0]),
    .d(\cu_ru/mepc [0]),
    .o(_al_u7723_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7724 (
    .a(_al_u7723_o),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/stvec [0]),
    .o(_al_u7724_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7725 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [0]),
    .d(\cu_ru/stval [0]),
    .o(_al_u7725_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7726 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[0]),
    .d(\cu_ru/mtval [0]),
    .o(_al_u7726_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7727 (
    .a(_al_u7722_o),
    .b(_al_u7724_o),
    .c(_al_u7725_o),
    .d(_al_u7726_o),
    .o(csr_data[0]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf55c))
    _al_u7728 (
    .a(_al_u3399_o),
    .b(_al_u6760_o),
    .c(id_ins[28]),
    .d(id_ins[27]),
    .o(_al_u7728_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(~D*B))"),
    .INIT(16'h0501))
    _al_u7729 (
    .a(\ins_dec/n71 ),
    .b(_al_u3938_o),
    .c(\ins_dec/n141_lutinv ),
    .d(_al_u7728_o),
    .o(_al_u7729_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u7730 (
    .a(_al_u7729_o),
    .b(\ins_dec/n149_lutinv ),
    .c(_al_u6059_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(_al_u7730_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7731 (
    .a(\ins_dec/n235 ),
    .b(_al_u7730_o),
    .o(_al_u7731_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~A*~(D*C))"),
    .INIT(16'hfbbb))
    _al_u7732 (
    .a(\ins_dec/n232 ),
    .b(_al_u7731_o),
    .c(_al_u3384_o),
    .d(_al_u3939_o),
    .o(\ins_dec/n126 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u7733 (
    .a(load_acc_fault),
    .b(_al_u2838_o),
    .c(_al_u2847_o),
    .o(_al_u7733_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u7734 (
    .a(\exu/load_addr_mis ),
    .b(\exu/store_addr_mis ),
    .c(_al_u7733_o),
    .o(_al_u7734_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u7735 (
    .a(_al_u6724_o),
    .b(_al_u7734_o),
    .c(_al_u6725_o),
    .d(_al_u7195_o),
    .o(ex_more_exception_neg_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7736 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[9]),
    .c(ex_exc_code[9]),
    .o(\exu/n71 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7737 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[8]),
    .c(ex_exc_code[8]),
    .o(\exu/n71 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7738 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[7]),
    .c(ex_exc_code[7]),
    .o(\exu/n71 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7739 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[63]),
    .o(\exu/n71 [63]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7740 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[62]),
    .o(\exu/n71 [62]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7741 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[61]),
    .o(\exu/n71 [61]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7742 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[60]),
    .o(\exu/n71 [60]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7743 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[6]),
    .c(ex_exc_code[6]),
    .o(\exu/n71 [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7744 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[59]),
    .o(\exu/n71 [59]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7745 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[58]),
    .o(\exu/n71 [58]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7746 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[57]),
    .o(\exu/n71 [57]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7747 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[56]),
    .o(\exu/n71 [56]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7748 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[55]),
    .o(\exu/n71 [55]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7749 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[54]),
    .o(\exu/n71 [54]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7750 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[53]),
    .o(\exu/n71 [53]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7751 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[52]),
    .o(\exu/n71 [52]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7752 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[51]),
    .o(\exu/n71 [51]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7753 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[50]),
    .o(\exu/n71 [50]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7754 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[5]),
    .c(ex_exc_code[5]),
    .o(\exu/n71 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7755 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[49]),
    .o(\exu/n71 [49]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7756 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[48]),
    .o(\exu/n71 [48]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7757 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[47]),
    .o(\exu/n71 [47]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7758 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[46]),
    .o(\exu/n71 [46]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7759 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[45]),
    .o(\exu/n71 [45]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7760 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[44]),
    .o(\exu/n71 [44]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7761 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[43]),
    .o(\exu/n71 [43]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7762 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[42]),
    .o(\exu/n71 [42]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7763 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[41]),
    .o(\exu/n71 [41]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7764 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[40]),
    .o(\exu/n71 [40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7765 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[4]),
    .c(ex_exc_code[4]),
    .o(\exu/n71 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7766 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[39]),
    .o(\exu/n71 [39]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7767 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[38]),
    .o(\exu/n71 [38]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7768 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[37]),
    .o(\exu/n71 [37]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7769 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[36]),
    .o(\exu/n71 [36]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7770 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[35]),
    .o(\exu/n71 [35]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7771 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[34]),
    .o(\exu/n71 [34]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7772 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[33]),
    .o(\exu/n71 [33]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7773 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[32]),
    .o(\exu/n71 [32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7774 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[31]),
    .c(ex_exc_code[31]),
    .o(\exu/n71 [31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7775 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[30]),
    .c(ex_exc_code[30]),
    .o(\exu/n71 [30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7776 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[3]),
    .c(ex_exc_code[3]),
    .o(\exu/n71 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7777 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[29]),
    .c(ex_exc_code[29]),
    .o(\exu/n71 [29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7778 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[28]),
    .c(ex_exc_code[28]),
    .o(\exu/n71 [28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7779 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[27]),
    .c(ex_exc_code[27]),
    .o(\exu/n71 [27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7780 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[26]),
    .c(ex_exc_code[26]),
    .o(\exu/n71 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7781 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[25]),
    .c(ex_exc_code[25]),
    .o(\exu/n71 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7782 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[24]),
    .c(ex_exc_code[24]),
    .o(\exu/n71 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7783 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[23]),
    .c(ex_exc_code[23]),
    .o(\exu/n71 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7784 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[22]),
    .c(ex_exc_code[22]),
    .o(\exu/n71 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7785 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[21]),
    .c(ex_exc_code[21]),
    .o(\exu/n71 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7786 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[20]),
    .c(ex_exc_code[20]),
    .o(\exu/n71 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7787 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[2]),
    .c(ex_exc_code[2]),
    .o(\exu/n71 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7788 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[19]),
    .c(ex_exc_code[19]),
    .o(\exu/n71 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7789 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[18]),
    .c(ex_exc_code[18]),
    .o(\exu/n71 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7790 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[17]),
    .c(ex_exc_code[17]),
    .o(\exu/n71 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7791 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[16]),
    .c(ex_exc_code[16]),
    .o(\exu/n71 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7792 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[15]),
    .c(ex_exc_code[15]),
    .o(\exu/n71 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7793 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[14]),
    .c(ex_exc_code[14]),
    .o(\exu/n71 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7794 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[13]),
    .c(ex_exc_code[13]),
    .o(\exu/n71 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7795 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[12]),
    .c(ex_exc_code[12]),
    .o(\exu/n71 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7796 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[11]),
    .c(ex_exc_code[11]),
    .o(\exu/n71 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7797 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[10]),
    .c(ex_exc_code[10]),
    .o(\exu/n71 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7798 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[1]),
    .c(ex_exc_code[1]),
    .o(\exu/n71 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u7799 (
    .a(ex_more_exception_neg_lutinv),
    .b(addr_ex[0]),
    .c(ex_exc_code[0]),
    .o(\exu/n71 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7800 (
    .a(_al_u6788_o),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/mcycle [9]),
    .d(\cu_ru/sepc [9]),
    .o(_al_u7800_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7801 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [9]),
    .d(\cu_ru/stval [9]),
    .o(_al_u7801_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7802 (
    .a(_al_u6764_o),
    .b(_al_u6791_o),
    .o(\cu_ru/read_mideleg_sel_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7803 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_mideleg_sel_lutinv ),
    .c(mtime_pad[9]),
    .d(\cu_ru/mideleg [9]),
    .o(_al_u7803_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7804 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/mtval [9]),
    .d(\cu_ru/stvec [9]),
    .o(_al_u7804_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7805 (
    .a(_al_u7800_o),
    .b(_al_u7801_o),
    .c(_al_u7803_o),
    .d(_al_u7804_o),
    .o(_al_u7805_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7806 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mscratch [9]),
    .d(\cu_ru/sscratch [9]),
    .o(_al_u7806_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7807 (
    .a(_al_u6765_o),
    .b(_al_u3388_o),
    .o(_al_u7807_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*~C))"),
    .INIT(16'h8880))
    _al_u7808 (
    .a(_al_u7478_o),
    .b(_al_u7807_o),
    .c(s_ext_int_pad),
    .d(\cu_ru/m_s_ip/seip ),
    .o(_al_u7808_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u7809 (
    .a(_al_u7806_o),
    .b(_al_u7808_o),
    .c(\cu_ru/read_satp_sel_lutinv ),
    .d(satp[9]),
    .o(_al_u7809_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7810 (
    .a(\cu_ru/read_mcause_sel_lutinv ),
    .b(\cu_ru/read_medeleg_sel_lutinv ),
    .c(\cu_ru/mcause [9]),
    .d(\cu_ru/medeleg [9]),
    .o(_al_u7810_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u7811 (
    .a(_al_u7810_o),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/n84 [10]),
    .d(\cu_ru/scause [9]),
    .o(_al_u7811_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7812 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mtvec_sel_lutinv ),
    .c(\cu_ru/minstret [9]),
    .d(\cu_ru/mtvec [9]),
    .o(_al_u7812_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7813 (
    .a(_al_u7805_o),
    .b(_al_u7809_o),
    .c(_al_u7811_o),
    .d(_al_u7812_o),
    .o(csr_data[9]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7814 (
    .a(csr_data[6]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[6]),
    .o(_al_u7814_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7815 (
    .a(_al_u7814_o),
    .b(rs1_data[6]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [6]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7816 (
    .a(csr_data[33]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[33]),
    .o(_al_u7816_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7817 (
    .a(rs1_data[33]),
    .b(_al_u7141_o),
    .o(_al_u7817_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7818 (
    .a(_al_u7816_o),
    .b(_al_u7817_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[31]),
    .o(\ins_dec/n272 [33]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7819 (
    .a(csr_data[32]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[32]),
    .o(_al_u7819_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7820 (
    .a(rs1_data[32]),
    .b(_al_u7141_o),
    .o(_al_u7820_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7821 (
    .a(_al_u7819_o),
    .b(_al_u7820_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[31]),
    .o(\ins_dec/n272 [32]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7822 (
    .a(csr_data[30]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[30]),
    .o(_al_u7822_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7823 (
    .a(rs1_data[30]),
    .b(_al_u7141_o),
    .o(_al_u7823_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7824 (
    .a(_al_u7822_o),
    .b(_al_u7823_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[30]),
    .o(\ins_dec/n272 [30]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7825 (
    .a(csr_data[28]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[28]),
    .o(_al_u7825_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7826 (
    .a(rs1_data[28]),
    .b(_al_u7141_o),
    .o(_al_u7826_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7827 (
    .a(_al_u7825_o),
    .b(_al_u7826_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[28]),
    .o(\ins_dec/n272 [28]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7828 (
    .a(csr_data[19]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[19]),
    .o(_al_u7828_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7829 (
    .a(rs1_data[19]),
    .b(_al_u7141_o),
    .o(_al_u7829_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7830 (
    .a(_al_u7828_o),
    .b(_al_u7829_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[19]),
    .o(\ins_dec/n272 [19]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7831 (
    .a(csr_data[14]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[14]),
    .o(_al_u7831_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7832 (
    .a(rs1_data[14]),
    .b(_al_u7141_o),
    .o(_al_u7832_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7833 (
    .a(_al_u7831_o),
    .b(_al_u7832_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(_al_u3216_o),
    .o(\ins_dec/n272 [14]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7834 (
    .a(csr_data[11]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[11]),
    .o(_al_u7834_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7835 (
    .a(_al_u7834_o),
    .b(rs1_data[11]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [11]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7836 (
    .a(csr_data[7]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[7]),
    .o(_al_u7836_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7837 (
    .a(_al_u7836_o),
    .b(rs1_data[7]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [7]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7838 (
    .a(csr_data[4]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[4]),
    .o(_al_u7838_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7839 (
    .a(_al_u7838_o),
    .b(rs1_data[4]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [4]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7840 (
    .a(csr_data[3]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[3]),
    .o(_al_u7840_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7841 (
    .a(_al_u7840_o),
    .b(rs1_data[3]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [3]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7842 (
    .a(csr_data[22]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[22]),
    .o(_al_u7842_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7843 (
    .a(rs1_data[22]),
    .b(_al_u7141_o),
    .o(_al_u7843_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7844 (
    .a(_al_u7842_o),
    .b(_al_u7843_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[22]),
    .o(\ins_dec/n272 [22]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7845 (
    .a(csr_data[20]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[20]),
    .o(_al_u7845_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7846 (
    .a(rs1_data[20]),
    .b(_al_u7141_o),
    .o(_al_u7846_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7847 (
    .a(_al_u7845_o),
    .b(_al_u7846_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[20]),
    .o(\ins_dec/n272 [20]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7848 (
    .a(csr_data[18]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[18]),
    .o(_al_u7848_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7849 (
    .a(rs1_data[18]),
    .b(_al_u7141_o),
    .o(_al_u7849_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7850 (
    .a(_al_u7848_o),
    .b(_al_u7849_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[18]),
    .o(\ins_dec/n272 [18]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7851 (
    .a(csr_data[17]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[17]),
    .o(_al_u7851_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7852 (
    .a(rs1_data[17]),
    .b(_al_u7141_o),
    .o(_al_u7852_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7853 (
    .a(_al_u7851_o),
    .b(_al_u7852_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(id_ins[17]),
    .o(\ins_dec/n272 [17]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u7854 (
    .a(csr_data[12]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[12]),
    .o(_al_u7854_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7855 (
    .a(rs1_data[12]),
    .b(_al_u7141_o),
    .o(_al_u7855_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~B*~A)*~(D)*~(C)+~(~B*~A)*D*~(C)+~(~(~B*~A))*D*C+~(~B*~A)*D*C)"),
    .INIT(16'hfe0e))
    _al_u7856 (
    .a(_al_u7854_o),
    .b(_al_u7855_o),
    .c(\ins_dec/op_lui_lutinv ),
    .d(_al_u3384_o),
    .o(\ins_dec/n272 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7857 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[1]),
    .d(\cu_ru/sscratch [1]),
    .o(_al_u7857_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7858 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_sepc_sel_lutinv ),
    .c(\cu_ru/sepc [1]),
    .d(\cu_ru/mtval [1]),
    .o(_al_u7858_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7859 (
    .a(_al_u7857_o),
    .b(_al_u7858_o),
    .c(\cu_ru/read_mepc_sel_lutinv ),
    .d(\cu_ru/mepc [1]),
    .o(_al_u7859_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7860 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/mcycle [1]),
    .d(\cu_ru/scause [1]),
    .o(_al_u7860_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7861 (
    .a(_al_u7860_o),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcause [1]),
    .o(_al_u7861_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7862 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mcycle [1]),
    .d(\cu_ru/mscratch [1]),
    .o(_al_u7862_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7863 (
    .a(_al_u7807_o),
    .b(\cu_ru/m_sip [1]),
    .o(_al_u7863_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7864 (
    .a(\cu_ru/read_medeleg_sel_lutinv ),
    .b(_al_u7863_o),
    .c(_al_u7478_o),
    .d(\cu_ru/medeleg [1]),
    .o(_al_u7864_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7865 (
    .a(_al_u7859_o),
    .b(_al_u7861_o),
    .c(_al_u7862_o),
    .d(_al_u7864_o),
    .o(_al_u7865_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7866 (
    .a(\cu_ru/read_time_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(mtime_pad[1]),
    .d(\cu_ru/stvec [1]),
    .o(_al_u7866_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u7867 (
    .a(_al_u7866_o),
    .b(\cu_ru/read_mtvec_sel_lutinv ),
    .c(\cu_ru/mtvec [1]),
    .o(_al_u7867_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7868 (
    .a(_al_u7401_o),
    .b(\cu_ru/read_stval_sel_lutinv ),
    .c(\cu_ru/mstatus [1]),
    .d(\cu_ru/stval [1]),
    .o(_al_u7868_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7869 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mideleg_sel_lutinv ),
    .c(\cu_ru/minstret [1]),
    .d(\cu_ru/mideleg [1]),
    .o(_al_u7869_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7870 (
    .a(_al_u7865_o),
    .b(_al_u7867_o),
    .c(_al_u7868_o),
    .d(_al_u7869_o),
    .o(csr_data[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7871 (
    .a(csr_data[8]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[8]),
    .o(_al_u7871_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7872 (
    .a(_al_u7871_o),
    .b(rs1_data[8]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u7873 (
    .a(\cu_ru/n84 [10]),
    .b(_al_u6769_o),
    .c(_al_u7478_o),
    .d(\cu_ru/m_sip [5]),
    .o(_al_u7873_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u7874 (
    .a(_al_u7873_o),
    .b(\cu_ru/n64 [32]),
    .c(\cu_ru/n90 [32]),
    .d(\cu_ru/mstatus [5]),
    .o(_al_u7874_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u7875 (
    .a(_al_u6763_o),
    .b(\cu_ru/read_mideleg_sel_lutinv ),
    .c(\cu_ru/minstret [5]),
    .d(\cu_ru/mideleg [5]),
    .o(_al_u7875_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7876 (
    .a(\cu_ru/read_mcycle_sel_lutinv ),
    .b(\cu_ru/read_mcause_sel_lutinv ),
    .c(\cu_ru/mcycle [5]),
    .d(\cu_ru/mcause [5]),
    .o(_al_u7876_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7877 (
    .a(\cu_ru/read_cycle_sel_lutinv ),
    .b(\cu_ru/read_scause_sel_lutinv ),
    .c(\cu_ru/mcycle [5]),
    .d(\cu_ru/scause [5]),
    .o(_al_u7877_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7878 (
    .a(\cu_ru/read_sscratch_sel_lutinv ),
    .b(\cu_ru/read_mscratch_sel_lutinv ),
    .c(\cu_ru/mscratch [5]),
    .d(\cu_ru/sscratch [5]),
    .o(_al_u7878_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7879 (
    .a(\cu_ru/read_medeleg_sel_lutinv ),
    .b(\cu_ru/read_satp_sel_lutinv ),
    .c(satp[5]),
    .d(\cu_ru/medeleg [5]),
    .o(_al_u7879_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7880 (
    .a(_al_u7876_o),
    .b(_al_u7877_o),
    .c(_al_u7878_o),
    .d(_al_u7879_o),
    .o(_al_u7880_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7881 (
    .a(\cu_ru/read_mtval_sel_lutinv ),
    .b(\cu_ru/read_mip_sel_lutinv ),
    .c(\cu_ru/m_sip [5]),
    .d(\cu_ru/mtval [5]),
    .o(_al_u7881_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7882 (
    .a(\cu_ru/read_stval_sel_lutinv ),
    .b(\cu_ru/read_mepc_sel_lutinv ),
    .c(\cu_ru/mepc [5]),
    .d(\cu_ru/stval [5]),
    .o(_al_u7882_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u7883 (
    .a(\cu_ru/read_mtvec_sel_lutinv ),
    .b(\cu_ru/read_time_sel_lutinv ),
    .c(mtime_pad[5]),
    .d(\cu_ru/mtvec [5]),
    .o(_al_u7883_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7884 (
    .a(\cu_ru/read_sepc_sel_lutinv ),
    .b(\cu_ru/read_stvec_sel_lutinv ),
    .c(\cu_ru/sepc [5]),
    .d(\cu_ru/stvec [5]),
    .o(_al_u7884_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u7885 (
    .a(_al_u7881_o),
    .b(_al_u7882_o),
    .c(_al_u7883_o),
    .d(_al_u7884_o),
    .o(_al_u7885_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u7886 (
    .a(_al_u7874_o),
    .b(_al_u7875_o),
    .c(_al_u7880_o),
    .d(_al_u7885_o),
    .o(csr_data[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7887 (
    .a(csr_data[2]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[2]),
    .o(_al_u7887_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7888 (
    .a(_al_u7887_o),
    .b(rs1_data[2]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [2]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7889 (
    .a(csr_data[0]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[0]),
    .o(_al_u7889_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7890 (
    .a(_al_u7889_o),
    .b(rs1_data[0]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [0]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7891 (
    .a(csr_data[9]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[9]),
    .o(_al_u7891_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7892 (
    .a(_al_u7891_o),
    .b(rs1_data[9]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [9]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7893 (
    .a(csr_data[1]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[1]),
    .o(_al_u7893_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7894 (
    .a(_al_u7893_o),
    .b(rs1_data[1]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [1]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h404c))
    _al_u7895 (
    .a(csr_data[5]),
    .b(_al_u7141_o),
    .c(id_system),
    .d(id_ins_pc[5]),
    .o(_al_u7895_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(~C*~B))"),
    .INIT(16'h0054))
    _al_u7896 (
    .a(_al_u7895_o),
    .b(rs1_data[5]),
    .c(_al_u7141_o),
    .d(\ins_dec/op_lui_lutinv ),
    .o(\ins_dec/n272 [5]));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u7897 (
    .a(\biu/l1d_out [15]),
    .b(uncache_data[15]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n2_lutinv ),
    .o(_al_u7897_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u7898 (
    .a(uncache_data[7]),
    .b(_al_u3224_o),
    .c(\exu/lsu/n0_lutinv ),
    .o(_al_u7898_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u7899 (
    .a(_al_u7898_o),
    .b(\biu/l1d_out [7]),
    .c(_al_u3224_o),
    .o(_al_u7899_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u7900 (
    .a(\biu/l1d_out [31]),
    .b(uncache_data[31]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u7900_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u7901 (
    .a(\biu/l1d_out [23]),
    .b(uncache_data[23]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u7901_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u7902 (
    .a(_al_u7897_o),
    .b(_al_u7899_o),
    .c(_al_u7900_o),
    .d(_al_u7901_o),
    .o(_al_u7902_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*(D@B))"),
    .INIT(16'h0208))
    _al_u7903 (
    .a(\exu/main_state [0]),
    .b(\exu/main_state [1]),
    .c(\exu/main_state [2]),
    .d(\exu/main_state [3]),
    .o(\exu/n60_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7904 (
    .a(ex_size[0]),
    .b(unsign),
    .o(\exu/lsu/n51 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u7905 (
    .a(_al_u7902_o),
    .b(\exu/n60_lutinv ),
    .c(\exu/lsu/n51 ),
    .o(_al_u7905_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u7906 (
    .a(\biu/l1d_out [33]),
    .b(_al_u3224_o),
    .c(uncache_data[33]),
    .o(_al_u7906_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u7907 (
    .a(\biu/l1d_out [25]),
    .b(_al_u3224_o),
    .c(uncache_data[25]),
    .o(_al_u7907_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h5300))
    _al_u7908 (
    .a(_al_u7906_o),
    .b(_al_u7907_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7908_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u7909 (
    .a(\biu/l1d_out [9]),
    .b(_al_u3224_o),
    .c(uncache_data[9]),
    .o(_al_u7909_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u7910 (
    .a(uncache_data[17]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [17]),
    .o(_al_u7910_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h00ca))
    _al_u7911 (
    .a(_al_u7909_o),
    .b(_al_u7910_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7911_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u7912 (
    .a(ex_size[2]),
    .b(unsign),
    .o(_al_u7912_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u7913 (
    .a(_al_u7908_o),
    .b(_al_u7911_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u7913_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7914 (
    .a(uncache_data[7]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n22 [7]));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u7915 (
    .a(uncache_data[31]),
    .b(uncache_data[15]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7915_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u7916 (
    .a(\exu/lsu/n22 [7]),
    .b(_al_u7915_o),
    .c(uncache_data[23]),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u7916_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7917 (
    .a(_al_u7916_o),
    .b(\exu/lsu/n51 ),
    .o(\exu/lsu/n52 [10]));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u7918 (
    .a(uncache_data[33]),
    .b(uncache_data[17]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7918_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u7919 (
    .a(uncache_data[9]),
    .b(uncache_data[25]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7919_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u7920 (
    .a(_al_u7918_o),
    .b(_al_u7919_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u7920_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u7921 (
    .a(\exu/lsu/n52 [10]),
    .b(_al_u7920_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u7921_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u7922 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[9]),
    .o(_al_u7922_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*A)))"),
    .INIT(16'h20f0))
    _al_u7923 (
    .a(_al_u7905_o),
    .b(_al_u7913_o),
    .c(_al_u7921_o),
    .d(_al_u7922_o),
    .o(_al_u7923_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u7924 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[9]),
    .d(ds2[9]),
    .o(_al_u7924_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7925 (
    .a(\exu/alu_au/sub_64 [9]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[9]),
    .o(_al_u7925_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7926 (
    .a(_al_u7924_o),
    .b(_al_u7925_o),
    .c(\exu/alu_au/add_64 [9]),
    .d(rd_data_add),
    .o(_al_u7926_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u7927 (
    .a(_al_u7926_o),
    .b(rd_data_xor),
    .c(ds1[9]),
    .d(ds2[9]),
    .o(_al_u7927_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(D*C)))"),
    .INIT(16'h3111))
    _al_u7928 (
    .a(_al_u7927_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/alu_and [9]),
    .d(rd_data_and),
    .o(_al_u7928_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u7929 (
    .a(data_rd[10]),
    .b(data_rd[9]),
    .c(shift_r),
    .o(\exu/n57 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u7930 (
    .a(_al_u2855_o),
    .b(\exu/n57 [9]),
    .c(data_rd[8]),
    .d(shift_l),
    .o(_al_u7930_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*~A))"),
    .INIT(8'hf4))
    _al_u7931 (
    .a(_al_u7923_o),
    .b(_al_u7928_o),
    .c(_al_u7930_o),
    .o(\exu/n64 [9]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u7932 (
    .a(\biu/l1d_out [24]),
    .b(_al_u3224_o),
    .c(uncache_data[24]),
    .o(_al_u7932_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u7933 (
    .a(\biu/l1d_out [16]),
    .b(_al_u3224_o),
    .c(uncache_data[16]),
    .o(_al_u7933_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u7934 (
    .a(_al_u7932_o),
    .b(_al_u7933_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7934_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u7935 (
    .a(uncache_data[8]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [8]),
    .o(_al_u7935_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u7936 (
    .a(\biu/l1d_out [32]),
    .b(_al_u3224_o),
    .c(uncache_data[32]),
    .o(_al_u7936_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ffa))
    _al_u7937 (
    .a(_al_u7935_o),
    .b(_al_u7936_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7937_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*A))"),
    .INIT(16'h7707))
    _al_u7938 (
    .a(_al_u7934_o),
    .b(_al_u7937_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u7938_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u7939 (
    .a(uncache_data[32]),
    .b(uncache_data[16]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7939_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u7940 (
    .a(uncache_data[8]),
    .b(uncache_data[24]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7940_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u7941 (
    .a(_al_u7939_o),
    .b(_al_u7940_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u7941_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u7942 (
    .a(\exu/lsu/n52 [10]),
    .b(_al_u7941_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u7942_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u7943 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[8]),
    .o(_al_u7943_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*A)))"),
    .INIT(16'h20f0))
    _al_u7944 (
    .a(_al_u7905_o),
    .b(_al_u7938_o),
    .c(_al_u7942_o),
    .d(_al_u7943_o),
    .o(_al_u7944_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u7945 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[8]),
    .d(ds2[8]),
    .o(_al_u7945_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7946 (
    .a(\exu/alu_au/sub_64 [8]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[8]),
    .o(_al_u7946_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7947 (
    .a(_al_u7945_o),
    .b(_al_u7946_o),
    .c(\exu/alu_au/add_64 [8]),
    .d(rd_data_add),
    .o(_al_u7947_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u7948 (
    .a(_al_u7947_o),
    .b(rd_data_xor),
    .c(ds1[8]),
    .d(ds2[8]),
    .o(_al_u7948_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(D*C)))"),
    .INIT(16'h3111))
    _al_u7949 (
    .a(_al_u7948_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/alu_and [8]),
    .d(rd_data_and),
    .o(_al_u7949_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u7950 (
    .a(data_rd[8]),
    .b(data_rd[9]),
    .c(shift_r),
    .o(\exu/n57 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u7951 (
    .a(_al_u2855_o),
    .b(\exu/n57 [8]),
    .c(data_rd[7]),
    .d(shift_l),
    .o(_al_u7951_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*~A))"),
    .INIT(8'hf4))
    _al_u7952 (
    .a(_al_u7944_o),
    .b(_al_u7949_o),
    .c(_al_u7951_o),
    .o(\exu/n64 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7953 (
    .a(_al_u3415_o),
    .b(\exu/n60_lutinv ),
    .c(_al_u7912_o),
    .o(_al_u7953_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7954 (
    .a(\exu/n60_lutinv ),
    .b(data_rd[7]),
    .o(_al_u7954_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(B*~A)))"),
    .INIT(16'h00f4))
    _al_u7955 (
    .a(_al_u7902_o),
    .b(_al_u7953_o),
    .c(_al_u7954_o),
    .d(\exu/n59_lutinv ),
    .o(_al_u7955_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7956 (
    .a(_al_u3415_o),
    .b(\exu/n59_lutinv ),
    .c(_al_u7912_o),
    .o(_al_u7956_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u7957 (
    .a(_al_u7916_o),
    .b(_al_u7956_o),
    .c(\exu/c_stb_lutinv ),
    .o(_al_u7957_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u7958 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[7]),
    .d(ds2[7]),
    .o(_al_u7958_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u7959 (
    .a(\exu/alu_au/sub_64 [7]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[7]),
    .o(_al_u7959_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u7960 (
    .a(_al_u7958_o),
    .b(_al_u7959_o),
    .c(\exu/alu_au/add_64 [7]),
    .d(rd_data_add),
    .o(_al_u7960_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u7961 (
    .a(_al_u7960_o),
    .b(rd_data_xor),
    .c(ds1[7]),
    .d(ds2[7]),
    .o(_al_u7961_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u7962 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[7]),
    .d(ds2[7]),
    .o(\exu/alu_au/n33 [7]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u7963 (
    .a(_al_u7961_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [7]),
    .o(_al_u7963_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u7964 (
    .a(data_rd[7]),
    .b(data_rd[8]),
    .c(shift_r),
    .o(\exu/n57 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u7965 (
    .a(_al_u2855_o),
    .b(\exu/n57 [7]),
    .c(data_rd[6]),
    .d(shift_l),
    .o(_al_u7965_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u7966 (
    .a(_al_u7955_o),
    .b(_al_u7957_o),
    .c(_al_u7963_o),
    .d(_al_u7965_o),
    .o(\exu/n64 [7]));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u7967 (
    .a(\biu/l1d_out [31]),
    .b(uncache_data[31]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u7967_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u7968 (
    .a(\biu/l1d_out [23]),
    .b(uncache_data[23]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n2_lutinv ),
    .o(_al_u7968_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u7969 (
    .a(\biu/l1d_out [15]),
    .b(uncache_data[15]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n0_lutinv ),
    .o(_al_u7969_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u7970 (
    .a(\biu/l1d_out [39]),
    .b(uncache_data[39]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u7970_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u7971 (
    .a(_al_u7967_o),
    .b(_al_u7968_o),
    .c(_al_u7969_o),
    .d(_al_u7970_o),
    .o(_al_u7971_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7972 (
    .a(ex_size[1]),
    .b(unsign),
    .o(\exu/lsu/n53 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7973 (
    .a(_al_u7971_o),
    .b(\exu/lsu/n53 ),
    .o(_al_u7973_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7974 (
    .a(uncache_data[47]),
    .b(_al_u3224_o),
    .o(_al_u7974_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~(~B*A)))"),
    .INIT(16'hf200))
    _al_u7975 (
    .a(\biu/l1d_out [47]),
    .b(_al_u3224_o),
    .c(_al_u7974_o),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u7975_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u7976 (
    .a(\biu/l1d_out [31]),
    .b(uncache_data[31]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n0_lutinv ),
    .o(_al_u7976_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u7977 (
    .a(\biu/l1d_out [39]),
    .b(uncache_data[39]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n2_lutinv ),
    .o(_al_u7977_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u7978 (
    .a(\biu/l1d_out [55]),
    .b(uncache_data[55]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u7978_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u7979 (
    .a(_al_u7975_o),
    .b(_al_u7976_o),
    .c(_al_u7977_o),
    .d(_al_u7978_o),
    .o(_al_u7979_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u7980 (
    .a(\biu/l1d_out [63]),
    .b(_al_u3224_o),
    .o(_al_u7980_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7981 (
    .a(uncache_data[63]),
    .b(_al_u3224_o),
    .o(_al_u7981_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u7982 (
    .a(_al_u7980_o),
    .b(_al_u7981_o),
    .o(_al_u7982_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7983 (
    .a(\exu/lsu/n0_lutinv ),
    .b(unsign),
    .o(\exu/lsu/mux27_b56_sel_is_3_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u7984 (
    .a(ex_size[2]),
    .b(unsign),
    .o(\exu/lsu/n56 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u7985 (
    .a(_al_u7979_o),
    .b(_al_u7982_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/lsu/n56 ),
    .o(_al_u7985_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u7986 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[63]),
    .o(_al_u7986_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u7987 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u7985_o),
    .d(_al_u7986_o),
    .o(_al_u7987_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u7988 (
    .a(uncache_data[31]),
    .b(uncache_data[23]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7988_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7989 (
    .a(uncache_data[15]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n22 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u7990 (
    .a(_al_u7988_o),
    .b(\exu/lsu/n22 [15]),
    .c(uncache_data[39]),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u7990_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u7991 (
    .a(\exu/lsu/n52 [10]),
    .b(_al_u7990_o),
    .c(\exu/lsu/n53 ),
    .o(_al_u7991_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7992 (
    .a(uncache_data[47]),
    .b(\exu/lsu/n5_lutinv ),
    .o(\exu/lsu/n25 [31]));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u7993 (
    .a(uncache_data[55]),
    .b(uncache_data[39]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u7993_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D*C))"),
    .INIT(16'h0111))
    _al_u7994 (
    .a(\exu/lsu/n25 [31]),
    .b(_al_u7993_o),
    .c(uncache_data[31]),
    .d(\exu/lsu/n0_lutinv ),
    .o(_al_u7994_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u7995 (
    .a(_al_u7991_o),
    .b(_al_u7994_o),
    .c(\exu/lsu/n56 ),
    .o(_al_u7995_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u7996 (
    .a(uncache_data[63]),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [63]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u7997 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [63]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u7997_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u7998 (
    .a(ex_size[2]),
    .b(shift_r),
    .o(\exu/mux27_b32_sel_is_1_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u7999 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[63]),
    .c(unsign),
    .o(\exu/n57 [63]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u8000 (
    .a(_al_u2855_o),
    .b(data_rd[63]),
    .c(ex_size[2]),
    .o(_al_u8000_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u8001 (
    .a(data_rd[62]),
    .b(ex_size[2]),
    .o(_al_u8001_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8002 (
    .a(\exu/n57 [63]),
    .b(_al_u8000_o),
    .c(_al_u8001_o),
    .d(shift_l),
    .o(_al_u8002_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u8003 (
    .a(rd_data_xor),
    .b(ds1[63]),
    .c(ds2[63]),
    .o(\exu/alu_au/n37 [63]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8004 (
    .a(\exu/alu_au/add_64 [63]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [63]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*~A))"),
    .INIT(16'h0203))
    _al_u8005 (
    .a(_al_u3459_o),
    .b(\exu/alu_au/n37 [63]),
    .c(\exu/alu_au/n31 [63]),
    .d(rd_data_add),
    .o(_al_u8005_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u8006 (
    .a(rd_data_or),
    .b(ds1[63]),
    .c(ds2[63]),
    .o(\exu/alu_au/n35 [63]));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u8007 (
    .a(\exu/c_stb_lutinv ),
    .b(\exu/alu_au/n35 [63]),
    .c(rd_data_ds1),
    .d(ds1[63]),
    .o(_al_u8007_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8008 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[63]),
    .d(ds2[63]),
    .o(\exu/alu_au/n33 [63]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*B*A))"),
    .INIT(16'h0f07))
    _al_u8009 (
    .a(_al_u8005_o),
    .b(_al_u8007_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [63]),
    .o(_al_u8009_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B*~A)))"),
    .INIT(16'hfbf0))
    _al_u8010 (
    .a(_al_u7987_o),
    .b(_al_u7997_o),
    .c(_al_u8002_o),
    .d(_al_u8009_o),
    .o(\exu/n64 [63]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u8011 (
    .a(uncache_data[62]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [62]),
    .o(_al_u8011_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u8012 (
    .a(_al_u7979_o),
    .b(_al_u8011_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/lsu/n56 ),
    .o(_al_u8012_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8013 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[62]),
    .o(_al_u8013_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u8014 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8012_o),
    .d(_al_u8013_o),
    .o(_al_u8014_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8015 (
    .a(uncache_data[62]),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [62]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8016 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [62]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8016_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8017 (
    .a(\exu/alu_au/add_64 [62]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [62]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8018 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3467_o),
    .c(\exu/alu_au/n31 [62]),
    .d(rd_data_add),
    .o(_al_u8018_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8019 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[62]),
    .o(_al_u8019_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8020 (
    .a(_al_u8019_o),
    .b(rd_data_xor),
    .c(ds1[62]),
    .d(ds2[62]),
    .o(_al_u8020_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8021 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[62]),
    .d(ds2[62]),
    .o(\exu/alu_au/n33 [62]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8022 (
    .a(_al_u8018_o),
    .b(_al_u8020_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [62]),
    .o(_al_u8022_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8023 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[62]),
    .c(data_rd[63]),
    .o(\exu/n57 [62]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8024 (
    .a(data_rd[61]),
    .b(data_rd[62]),
    .c(ex_size[2]),
    .o(\exu/n54 [30]));
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    .INIT(16'hc088))
    _al_u8025 (
    .a(\exu/n57 [62]),
    .b(_al_u2855_o),
    .c(\exu/n54 [30]),
    .d(shift_l),
    .o(_al_u8025_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8026 (
    .a(_al_u8014_o),
    .b(_al_u8016_o),
    .c(_al_u8022_o),
    .d(_al_u8025_o),
    .o(\exu/n64 [62]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u8027 (
    .a(\biu/l1d_out [61]),
    .b(_al_u3224_o),
    .o(_al_u8027_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8028 (
    .a(uncache_data[61]),
    .b(_al_u3224_o),
    .o(_al_u8028_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u8029 (
    .a(_al_u8027_o),
    .b(_al_u8028_o),
    .o(_al_u8029_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u8030 (
    .a(_al_u7979_o),
    .b(_al_u8029_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/lsu/n56 ),
    .o(_al_u8030_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8031 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[61]),
    .o(_al_u8031_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u8032 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8030_o),
    .d(_al_u8031_o),
    .o(_al_u8032_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8033 (
    .a(uncache_data[61]),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [61]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8034 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [61]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8034_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8035 (
    .a(\exu/alu_au/add_64 [61]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [61]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8036 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3475_o),
    .c(\exu/alu_au/n31 [61]),
    .d(rd_data_add),
    .o(_al_u8036_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8037 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[61]),
    .o(_al_u8037_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8038 (
    .a(_al_u8037_o),
    .b(rd_data_xor),
    .c(ds1[61]),
    .d(ds2[61]),
    .o(_al_u8038_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8039 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[61]),
    .d(ds2[61]),
    .o(\exu/alu_au/n33 [61]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8040 (
    .a(_al_u8036_o),
    .b(_al_u8038_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [61]),
    .o(_al_u8040_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u8041 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[61]),
    .c(data_rd[62]),
    .o(_al_u8041_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8042 (
    .a(data_rd[60]),
    .b(data_rd[61]),
    .c(ex_size[2]),
    .o(_al_u8042_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    .INIT(16'h0c44))
    _al_u8043 (
    .a(_al_u8041_o),
    .b(_al_u2855_o),
    .c(_al_u8042_o),
    .d(shift_l),
    .o(_al_u8043_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8044 (
    .a(_al_u8032_o),
    .b(_al_u8034_o),
    .c(_al_u8040_o),
    .d(_al_u8043_o),
    .o(\exu/n64 [61]));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8045 (
    .a(\biu/l1d_out [60]),
    .b(uncache_data[60]),
    .c(_al_u3224_o),
    .d(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(_al_u8045_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8046 (
    .a(_al_u7979_o),
    .b(_al_u8045_o),
    .c(\exu/lsu/n56 ),
    .o(_al_u8046_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8047 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[60]),
    .o(_al_u8047_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u8048 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8046_o),
    .d(_al_u8047_o),
    .o(_al_u8048_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8049 (
    .a(uncache_data[60]),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [60]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8050 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [60]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8050_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8051 (
    .a(\exu/alu_au/add_64 [60]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [60]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8052 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3483_o),
    .c(\exu/alu_au/n31 [60]),
    .d(rd_data_add),
    .o(_al_u8052_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8053 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[60]),
    .o(_al_u8053_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8054 (
    .a(_al_u8053_o),
    .b(rd_data_xor),
    .c(ds1[60]),
    .d(ds2[60]),
    .o(_al_u8054_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8055 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[60]),
    .d(ds2[60]),
    .o(\exu/alu_au/n33 [60]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8056 (
    .a(_al_u8052_o),
    .b(_al_u8054_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [60]),
    .o(_al_u8056_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u8057 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[60]),
    .c(data_rd[61]),
    .o(_al_u8057_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8058 (
    .a(data_rd[59]),
    .b(data_rd[60]),
    .c(ex_size[2]),
    .o(_al_u8058_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    .INIT(16'h0c44))
    _al_u8059 (
    .a(_al_u8057_o),
    .b(_al_u2855_o),
    .c(_al_u8058_o),
    .d(shift_l),
    .o(_al_u8059_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8060 (
    .a(_al_u8048_o),
    .b(_al_u8050_o),
    .c(_al_u8056_o),
    .d(_al_u8059_o),
    .o(\exu/n64 [60]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8061 (
    .a(uncache_data[59]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [59]),
    .o(_al_u8061_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u8062 (
    .a(_al_u7979_o),
    .b(_al_u8061_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/lsu/n56 ),
    .o(_al_u8062_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8063 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[59]),
    .o(_al_u8063_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u8064 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8062_o),
    .d(_al_u8063_o),
    .o(_al_u8064_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8065 (
    .a(uncache_data[59]),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [59]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8066 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [59]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8066_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8067 (
    .a(\exu/alu_au/add_64 [59]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [59]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8068 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3498_o),
    .c(\exu/alu_au/n31 [59]),
    .d(rd_data_add),
    .o(_al_u8068_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8069 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[59]),
    .o(_al_u8069_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8070 (
    .a(_al_u8069_o),
    .b(rd_data_xor),
    .c(ds1[59]),
    .d(ds2[59]),
    .o(_al_u8070_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8071 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[59]),
    .d(ds2[59]),
    .o(\exu/alu_au/n33 [59]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8072 (
    .a(_al_u8068_o),
    .b(_al_u8070_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [59]),
    .o(_al_u8072_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8073 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[59]),
    .c(data_rd[60]),
    .o(\exu/n57 [59]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8074 (
    .a(data_rd[58]),
    .b(data_rd[59]),
    .c(ex_size[2]),
    .o(_al_u8074_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8075 (
    .a(\exu/n57 [59]),
    .b(_al_u2855_o),
    .c(_al_u8074_o),
    .d(shift_l),
    .o(_al_u8075_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8076 (
    .a(_al_u8064_o),
    .b(_al_u8066_o),
    .c(_al_u8072_o),
    .d(_al_u8075_o),
    .o(\exu/n64 [59]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8077 (
    .a(uncache_data[58]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [58]),
    .o(_al_u8077_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u8078 (
    .a(_al_u7979_o),
    .b(_al_u8077_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/lsu/n56 ),
    .o(_al_u8078_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8079 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[58]),
    .o(_al_u8079_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u8080 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8078_o),
    .d(_al_u8079_o),
    .o(_al_u8080_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8081 (
    .a(uncache_data[58]),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [58]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8082 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [58]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8082_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8083 (
    .a(\exu/alu_au/add_64 [58]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [58]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8084 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3506_o),
    .c(\exu/alu_au/n31 [58]),
    .d(rd_data_add),
    .o(_al_u8084_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8085 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[58]),
    .o(_al_u8085_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8086 (
    .a(_al_u8085_o),
    .b(rd_data_xor),
    .c(ds1[58]),
    .d(ds2[58]),
    .o(_al_u8086_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8087 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[58]),
    .d(ds2[58]),
    .o(\exu/alu_au/n33 [58]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8088 (
    .a(_al_u8084_o),
    .b(_al_u8086_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [58]),
    .o(_al_u8088_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8089 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[58]),
    .c(data_rd[59]),
    .o(\exu/n57 [58]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8090 (
    .a(data_rd[57]),
    .b(data_rd[58]),
    .c(ex_size[2]),
    .o(_al_u8090_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8091 (
    .a(\exu/n57 [58]),
    .b(_al_u2855_o),
    .c(_al_u8090_o),
    .d(shift_l),
    .o(_al_u8091_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8092 (
    .a(_al_u8080_o),
    .b(_al_u8082_o),
    .c(_al_u8088_o),
    .d(_al_u8091_o),
    .o(\exu/n64 [58]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u8093 (
    .a(\biu/l1d_out [57]),
    .b(_al_u3224_o),
    .c(uncache_data[57]),
    .o(_al_u8093_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u8094 (
    .a(_al_u7979_o),
    .b(_al_u8093_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/lsu/n56 ),
    .o(_al_u8094_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8095 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[57]),
    .o(_al_u8095_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u8096 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8094_o),
    .d(_al_u8095_o),
    .o(_al_u8096_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8097 (
    .a(uncache_data[57]),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [57]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8098 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [57]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8098_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8099 (
    .a(\exu/alu_au/add_64 [57]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [57]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8100 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3514_o),
    .c(\exu/alu_au/n31 [57]),
    .d(rd_data_add),
    .o(_al_u8100_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8101 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[57]),
    .o(_al_u8101_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8102 (
    .a(_al_u8101_o),
    .b(rd_data_xor),
    .c(ds1[57]),
    .d(ds2[57]),
    .o(_al_u8102_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8103 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[57]),
    .d(ds2[57]),
    .o(\exu/alu_au/n33 [57]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8104 (
    .a(_al_u8100_o),
    .b(_al_u8102_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [57]),
    .o(_al_u8104_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8105 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[57]),
    .c(data_rd[58]),
    .o(\exu/n57 [57]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8106 (
    .a(data_rd[56]),
    .b(data_rd[57]),
    .c(ex_size[2]),
    .o(_al_u8106_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8107 (
    .a(\exu/n57 [57]),
    .b(_al_u2855_o),
    .c(_al_u8106_o),
    .d(shift_l),
    .o(_al_u8107_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8108 (
    .a(_al_u8096_o),
    .b(_al_u8098_o),
    .c(_al_u8104_o),
    .d(_al_u8107_o),
    .o(\exu/n64 [57]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8109 (
    .a(uncache_data[56]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [56]),
    .o(_al_u8109_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u8110 (
    .a(_al_u7979_o),
    .b(_al_u8109_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/lsu/n56 ),
    .o(_al_u8110_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8111 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[56]),
    .o(_al_u8111_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u8112 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8110_o),
    .d(_al_u8111_o),
    .o(_al_u8112_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8113 (
    .a(uncache_data[56]),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [56]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8114 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [56]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8114_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8115 (
    .a(\exu/alu_au/add_64 [56]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [56]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8116 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3522_o),
    .c(\exu/alu_au/n31 [56]),
    .d(rd_data_add),
    .o(_al_u8116_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8117 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[56]),
    .o(_al_u8117_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8118 (
    .a(_al_u8117_o),
    .b(rd_data_xor),
    .c(ds1[56]),
    .d(ds2[56]),
    .o(_al_u8118_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8119 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[56]),
    .d(ds2[56]),
    .o(\exu/alu_au/n33 [56]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8120 (
    .a(_al_u8116_o),
    .b(_al_u8118_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [56]),
    .o(_al_u8120_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8121 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[56]),
    .c(data_rd[57]),
    .o(\exu/n57 [56]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8122 (
    .a(data_rd[55]),
    .b(data_rd[56]),
    .c(ex_size[2]),
    .o(_al_u8122_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8123 (
    .a(\exu/n57 [56]),
    .b(_al_u2855_o),
    .c(_al_u8122_o),
    .d(shift_l),
    .o(_al_u8123_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8124 (
    .a(_al_u8112_o),
    .b(_al_u8114_o),
    .c(_al_u8120_o),
    .d(_al_u8123_o),
    .o(\exu/n64 [56]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8125 (
    .a(_al_u7979_o),
    .b(\exu/lsu/n56 ),
    .o(_al_u8125_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u8126 (
    .a(_al_u7902_o),
    .b(_al_u7971_o),
    .c(\exu/lsu/n51 ),
    .d(\exu/lsu/n53 ),
    .o(_al_u8126_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8127 (
    .a(\exu/lsu/n2_lutinv ),
    .b(unsign),
    .o(_al_u8127_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u8128 (
    .a(_al_u7980_o),
    .b(_al_u7981_o),
    .c(_al_u8127_o),
    .o(_al_u8128_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8129 (
    .a(\biu/l1d_out [55]),
    .b(uncache_data[55]),
    .c(_al_u3224_o),
    .o(_al_u8129_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*~B))"),
    .INIT(16'h4500))
    _al_u8130 (
    .a(_al_u8128_o),
    .b(_al_u8129_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/n60_lutinv ),
    .o(_al_u8130_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8131 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[55]),
    .o(_al_u8131_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8132 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8130_o),
    .d(_al_u8131_o),
    .o(_al_u8132_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u8133 (
    .a(uncache_data[63]),
    .b(uncache_data[55]),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(_al_u8127_o),
    .o(_al_u8133_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u8134 (
    .a(_al_u7995_o),
    .b(_al_u8133_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8134_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8135 (
    .a(\exu/alu_au/add_64 [55]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [55]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8136 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3530_o),
    .c(\exu/alu_au/n31 [55]),
    .d(rd_data_add),
    .o(_al_u8136_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8137 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[55]),
    .o(_al_u8137_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8138 (
    .a(_al_u8137_o),
    .b(rd_data_xor),
    .c(ds1[55]),
    .d(ds2[55]),
    .o(_al_u8138_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8139 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[55]),
    .d(ds2[55]),
    .o(\exu/alu_au/n33 [55]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8140 (
    .a(_al_u8136_o),
    .b(_al_u8138_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [55]),
    .o(_al_u8140_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8141 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[55]),
    .c(data_rd[56]),
    .o(\exu/n57 [55]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8142 (
    .a(data_rd[54]),
    .b(data_rd[55]),
    .c(ex_size[2]),
    .o(_al_u8142_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8143 (
    .a(\exu/n57 [55]),
    .b(_al_u2855_o),
    .c(_al_u8142_o),
    .d(shift_l),
    .o(_al_u8143_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8144 (
    .a(_al_u8132_o),
    .b(_al_u8134_o),
    .c(_al_u8140_o),
    .d(_al_u8143_o),
    .o(\exu/n64 [55]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u8145 (
    .a(_al_u8011_o),
    .b(_al_u8127_o),
    .c(\exu/n60_lutinv ),
    .o(_al_u8145_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u8146 (
    .a(\biu/l1d_out [54]),
    .b(_al_u3224_o),
    .c(uncache_data[54]),
    .o(_al_u8146_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u8147 (
    .a(_al_u8145_o),
    .b(_al_u8146_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(_al_u8147_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8148 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[54]),
    .o(_al_u8148_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8149 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8147_o),
    .d(_al_u8148_o),
    .o(_al_u8149_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u8150 (
    .a(uncache_data[62]),
    .b(uncache_data[54]),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(_al_u8127_o),
    .o(_al_u8150_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u8151 (
    .a(_al_u7995_o),
    .b(_al_u8150_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8151_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8152 (
    .a(\exu/alu_au/add_64 [54]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [54]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8153 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3538_o),
    .c(\exu/alu_au/n31 [54]),
    .d(rd_data_add),
    .o(_al_u8153_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8154 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[54]),
    .o(_al_u8154_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8155 (
    .a(_al_u8154_o),
    .b(rd_data_xor),
    .c(ds1[54]),
    .d(ds2[54]),
    .o(_al_u8155_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8156 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[54]),
    .d(ds2[54]),
    .o(\exu/alu_au/n33 [54]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8157 (
    .a(_al_u8153_o),
    .b(_al_u8155_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [54]),
    .o(_al_u8157_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8158 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[54]),
    .c(data_rd[55]),
    .o(\exu/n57 [54]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8159 (
    .a(data_rd[53]),
    .b(data_rd[54]),
    .c(ex_size[2]),
    .o(_al_u8159_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8160 (
    .a(\exu/n57 [54]),
    .b(_al_u2855_o),
    .c(_al_u8159_o),
    .d(shift_l),
    .o(_al_u8160_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8161 (
    .a(_al_u8149_o),
    .b(_al_u8151_o),
    .c(_al_u8157_o),
    .d(_al_u8160_o),
    .o(\exu/n64 [54]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u8162 (
    .a(_al_u8027_o),
    .b(_al_u8028_o),
    .c(_al_u8127_o),
    .o(_al_u8162_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8163 (
    .a(uncache_data[53]),
    .b(_al_u3224_o),
    .o(_al_u8163_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8164 (
    .a(\biu/l1d_out [53]),
    .b(_al_u3224_o),
    .c(_al_u8163_o),
    .o(_al_u8164_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u8165 (
    .a(_al_u8162_o),
    .b(_al_u8164_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/n60_lutinv ),
    .o(_al_u8165_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8166 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[53]),
    .o(_al_u8166_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8167 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8165_o),
    .d(_al_u8166_o),
    .o(_al_u8167_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u8168 (
    .a(uncache_data[61]),
    .b(uncache_data[53]),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(_al_u8127_o),
    .o(_al_u8168_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u8169 (
    .a(_al_u7995_o),
    .b(_al_u8168_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8169_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8170 (
    .a(\exu/alu_au/add_64 [53]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [53]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8171 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3546_o),
    .c(\exu/alu_au/n31 [53]),
    .d(rd_data_add),
    .o(_al_u8171_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8172 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[53]),
    .o(_al_u8172_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8173 (
    .a(_al_u8172_o),
    .b(rd_data_xor),
    .c(ds1[53]),
    .d(ds2[53]),
    .o(_al_u8173_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8174 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[53]),
    .d(ds2[53]),
    .o(\exu/alu_au/n33 [53]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8175 (
    .a(_al_u8171_o),
    .b(_al_u8173_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [53]),
    .o(_al_u8175_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8176 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[53]),
    .c(data_rd[54]),
    .o(\exu/n57 [53]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8177 (
    .a(data_rd[52]),
    .b(data_rd[53]),
    .c(ex_size[2]),
    .o(_al_u8177_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8178 (
    .a(\exu/n57 [53]),
    .b(_al_u2855_o),
    .c(_al_u8177_o),
    .d(shift_l),
    .o(_al_u8178_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8179 (
    .a(_al_u8167_o),
    .b(_al_u8169_o),
    .c(_al_u8175_o),
    .d(_al_u8178_o),
    .o(\exu/n64 [53]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8180 (
    .a(\biu/l1d_out [52]),
    .b(uncache_data[52]),
    .c(_al_u3224_o),
    .o(_al_u8180_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8181 (
    .a(\biu/l1d_out [60]),
    .b(uncache_data[60]),
    .c(_al_u3224_o),
    .d(_al_u8127_o),
    .o(_al_u8181_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(C*A))"),
    .INIT(16'h1300))
    _al_u8182 (
    .a(_al_u8180_o),
    .b(_al_u8181_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/n60_lutinv ),
    .o(_al_u8182_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8183 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[52]),
    .o(_al_u8183_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8184 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8182_o),
    .d(_al_u8183_o),
    .o(_al_u8184_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u8185 (
    .a(uncache_data[60]),
    .b(uncache_data[52]),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(_al_u8127_o),
    .o(_al_u8185_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u8186 (
    .a(_al_u7995_o),
    .b(_al_u8185_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8186_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8187 (
    .a(\exu/alu_au/add_64 [52]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [52]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8188 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3554_o),
    .c(\exu/alu_au/n31 [52]),
    .d(rd_data_add),
    .o(_al_u8188_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8189 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[52]),
    .o(_al_u8189_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8190 (
    .a(_al_u8189_o),
    .b(rd_data_xor),
    .c(ds1[52]),
    .d(ds2[52]),
    .o(_al_u8190_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8191 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[52]),
    .d(ds2[52]),
    .o(\exu/alu_au/n33 [52]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8192 (
    .a(_al_u8188_o),
    .b(_al_u8190_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [52]),
    .o(_al_u8192_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8193 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[52]),
    .c(data_rd[53]),
    .o(\exu/n57 [52]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8194 (
    .a(data_rd[51]),
    .b(data_rd[52]),
    .c(ex_size[2]),
    .o(_al_u8194_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8195 (
    .a(\exu/n57 [52]),
    .b(_al_u2855_o),
    .c(_al_u8194_o),
    .d(shift_l),
    .o(_al_u8195_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8196 (
    .a(_al_u8184_o),
    .b(_al_u8186_o),
    .c(_al_u8192_o),
    .d(_al_u8195_o),
    .o(\exu/n64 [52]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8197 (
    .a(_al_u8061_o),
    .b(_al_u8127_o),
    .c(\exu/n60_lutinv ),
    .o(_al_u8197_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u8198 (
    .a(uncache_data[51]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [51]),
    .o(_al_u8198_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u8199 (
    .a(_al_u8197_o),
    .b(_al_u8198_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(_al_u8199_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8200 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[51]),
    .o(_al_u8200_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8201 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8199_o),
    .d(_al_u8200_o),
    .o(_al_u8201_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u8202 (
    .a(uncache_data[59]),
    .b(uncache_data[51]),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(_al_u8127_o),
    .o(_al_u8202_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u8203 (
    .a(_al_u7995_o),
    .b(_al_u8202_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8203_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8204 (
    .a(\exu/alu_au/add_64 [51]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [51]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8205 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3562_o),
    .c(\exu/alu_au/n31 [51]),
    .d(rd_data_add),
    .o(_al_u8205_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8206 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[51]),
    .o(_al_u8206_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8207 (
    .a(_al_u8206_o),
    .b(rd_data_xor),
    .c(ds1[51]),
    .d(ds2[51]),
    .o(_al_u8207_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8208 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[51]),
    .d(ds2[51]),
    .o(\exu/alu_au/n33 [51]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8209 (
    .a(_al_u8205_o),
    .b(_al_u8207_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [51]),
    .o(_al_u8209_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8210 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[51]),
    .c(data_rd[52]),
    .o(\exu/n57 [51]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8211 (
    .a(data_rd[50]),
    .b(data_rd[51]),
    .c(ex_size[2]),
    .o(_al_u8211_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8212 (
    .a(\exu/n57 [51]),
    .b(_al_u2855_o),
    .c(_al_u8211_o),
    .d(shift_l),
    .o(_al_u8212_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8213 (
    .a(_al_u8201_o),
    .b(_al_u8203_o),
    .c(_al_u8209_o),
    .d(_al_u8212_o),
    .o(\exu/n64 [51]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8214 (
    .a(_al_u8077_o),
    .b(_al_u8127_o),
    .c(\exu/n60_lutinv ),
    .o(_al_u8214_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u8215 (
    .a(\biu/l1d_out [50]),
    .b(_al_u3224_o),
    .c(uncache_data[50]),
    .o(_al_u8215_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u8216 (
    .a(_al_u8214_o),
    .b(_al_u8215_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(_al_u8216_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8217 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[50]),
    .o(_al_u8217_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8218 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8216_o),
    .d(_al_u8217_o),
    .o(_al_u8218_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u8219 (
    .a(uncache_data[58]),
    .b(uncache_data[50]),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(_al_u8127_o),
    .o(_al_u8219_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u8220 (
    .a(_al_u7995_o),
    .b(_al_u8219_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8220_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8221 (
    .a(\exu/alu_au/add_64 [50]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [50]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8222 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3570_o),
    .c(\exu/alu_au/n31 [50]),
    .d(rd_data_add),
    .o(_al_u8222_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8223 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[50]),
    .o(_al_u8223_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8224 (
    .a(_al_u8223_o),
    .b(rd_data_xor),
    .c(ds1[50]),
    .d(ds2[50]),
    .o(_al_u8224_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8225 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[50]),
    .d(ds2[50]),
    .o(\exu/alu_au/n33 [50]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8226 (
    .a(_al_u8222_o),
    .b(_al_u8224_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [50]),
    .o(_al_u8226_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8227 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[50]),
    .c(data_rd[51]),
    .o(\exu/n57 [50]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8228 (
    .a(data_rd[49]),
    .b(data_rd[50]),
    .c(ex_size[2]),
    .o(_al_u8228_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8229 (
    .a(\exu/n57 [50]),
    .b(_al_u2855_o),
    .c(_al_u8228_o),
    .d(shift_l),
    .o(_al_u8229_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8230 (
    .a(_al_u8218_o),
    .b(_al_u8220_o),
    .c(_al_u8226_o),
    .d(_al_u8229_o),
    .o(\exu/n64 [50]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8231 (
    .a(_al_u8093_o),
    .b(_al_u8127_o),
    .o(_al_u8231_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8232 (
    .a(uncache_data[49]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [49]),
    .o(_al_u8232_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*~B))"),
    .INIT(16'h4500))
    _al_u8233 (
    .a(_al_u8231_o),
    .b(_al_u8232_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/n60_lutinv ),
    .o(_al_u8233_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8234 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[49]),
    .o(_al_u8234_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8235 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8233_o),
    .d(_al_u8234_o),
    .o(_al_u8235_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u8236 (
    .a(uncache_data[57]),
    .b(uncache_data[49]),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(_al_u8127_o),
    .o(_al_u8236_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u8237 (
    .a(_al_u7995_o),
    .b(_al_u8236_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8237_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8238 (
    .a(\exu/alu_au/add_64 [49]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [49]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8239 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3585_o),
    .c(\exu/alu_au/n31 [49]),
    .d(rd_data_add),
    .o(_al_u8239_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8240 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[49]),
    .o(_al_u8240_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8241 (
    .a(_al_u8240_o),
    .b(rd_data_xor),
    .c(ds1[49]),
    .d(ds2[49]),
    .o(_al_u8241_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8242 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[49]),
    .d(ds2[49]),
    .o(\exu/alu_au/n33 [49]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8243 (
    .a(_al_u8239_o),
    .b(_al_u8241_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [49]),
    .o(_al_u8243_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8244 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[49]),
    .c(data_rd[50]),
    .o(\exu/n57 [49]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8245 (
    .a(data_rd[48]),
    .b(data_rd[49]),
    .c(ex_size[2]),
    .o(_al_u8245_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8246 (
    .a(\exu/n57 [49]),
    .b(_al_u2855_o),
    .c(_al_u8245_o),
    .d(shift_l),
    .o(_al_u8246_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8247 (
    .a(_al_u8235_o),
    .b(_al_u8237_o),
    .c(_al_u8243_o),
    .d(_al_u8246_o),
    .o(\exu/n64 [49]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8248 (
    .a(_al_u8109_o),
    .b(_al_u8127_o),
    .c(\exu/n60_lutinv ),
    .o(_al_u8248_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u8249 (
    .a(\biu/l1d_out [48]),
    .b(_al_u3224_o),
    .c(uncache_data[48]),
    .o(_al_u8249_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u8250 (
    .a(_al_u8248_o),
    .b(_al_u8249_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(_al_u8250_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8251 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[48]),
    .o(_al_u8251_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8252 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8250_o),
    .d(_al_u8251_o),
    .o(_al_u8252_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u8253 (
    .a(uncache_data[56]),
    .b(uncache_data[48]),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(_al_u8127_o),
    .o(_al_u8253_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*A)))"),
    .INIT(16'h080f))
    _al_u8254 (
    .a(_al_u7995_o),
    .b(_al_u8253_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8254_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8255 (
    .a(\exu/alu_au/add_64 [48]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [48]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8256 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3593_o),
    .c(\exu/alu_au/n31 [48]),
    .d(rd_data_add),
    .o(_al_u8256_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8257 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[48]),
    .o(_al_u8257_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8258 (
    .a(_al_u8257_o),
    .b(rd_data_xor),
    .c(ds1[48]),
    .d(ds2[48]),
    .o(_al_u8258_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8259 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[48]),
    .d(ds2[48]),
    .o(\exu/alu_au/n33 [48]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8260 (
    .a(_al_u8256_o),
    .b(_al_u8258_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [48]),
    .o(_al_u8260_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8261 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[48]),
    .c(data_rd[49]),
    .o(\exu/n57 [48]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8262 (
    .a(data_rd[47]),
    .b(data_rd[48]),
    .c(ex_size[2]),
    .o(_al_u8262_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8263 (
    .a(\exu/n57 [48]),
    .b(_al_u2855_o),
    .c(_al_u8262_o),
    .d(shift_l),
    .o(_al_u8263_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8264 (
    .a(_al_u8252_o),
    .b(_al_u8254_o),
    .c(_al_u8260_o),
    .d(_al_u8263_o),
    .o(\exu/n64 [48]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u8265 (
    .a(_al_u7980_o),
    .b(_al_u7981_o),
    .c(\exu/lsu/n5_lutinv ),
    .o(_al_u8265_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8266 (
    .a(_al_u8129_o),
    .b(\exu/lsu/n2_lutinv ),
    .o(_al_u8266_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u8267 (
    .a(\biu/l1d_out [47]),
    .b(_al_u3224_o),
    .c(_al_u7974_o),
    .o(_al_u8267_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8268 (
    .a(_al_u8267_o),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .c(\exu/n60_lutinv ),
    .o(_al_u8268_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*~A)))"),
    .INIT(16'h10f0))
    _al_u8269 (
    .a(_al_u8265_o),
    .b(_al_u8266_o),
    .c(_al_u8268_o),
    .d(unsign),
    .o(_al_u8269_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8270 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[47]),
    .o(_al_u8270_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8271 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8269_o),
    .d(_al_u8270_o),
    .o(_al_u8271_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8272 (
    .a(uncache_data[63]),
    .b(uncache_data[47]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8272_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u8273 (
    .a(_al_u8272_o),
    .b(uncache_data[55]),
    .c(\exu/lsu/n2_lutinv ),
    .d(unsign),
    .o(\exu/lsu/n59 [47]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8274 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [47]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8274_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8275 (
    .a(\exu/alu_au/add_64 [47]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [47]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8276 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3601_o),
    .c(\exu/alu_au/n31 [47]),
    .d(rd_data_add),
    .o(_al_u8276_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8277 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[47]),
    .o(_al_u8277_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8278 (
    .a(_al_u8277_o),
    .b(rd_data_xor),
    .c(ds1[47]),
    .d(ds2[47]),
    .o(_al_u8278_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8279 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[47]),
    .d(ds2[47]),
    .o(\exu/alu_au/n33 [47]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8280 (
    .a(_al_u8276_o),
    .b(_al_u8278_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [47]),
    .o(_al_u8280_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8281 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[47]),
    .c(data_rd[48]),
    .o(\exu/n57 [47]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8282 (
    .a(data_rd[46]),
    .b(data_rd[47]),
    .c(ex_size[2]),
    .o(_al_u8282_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8283 (
    .a(\exu/n57 [47]),
    .b(_al_u2855_o),
    .c(_al_u8282_o),
    .d(shift_l),
    .o(_al_u8283_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8284 (
    .a(_al_u8271_o),
    .b(_al_u8274_o),
    .c(_al_u8280_o),
    .d(_al_u8283_o),
    .o(\exu/n64 [47]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf5cf))
    _al_u8285 (
    .a(_al_u8011_o),
    .b(_al_u8146_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8285_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8286 (
    .a(uncache_data[46]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [46]),
    .o(_al_u8286_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8287 (
    .a(_al_u8286_o),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .c(\exu/n60_lutinv ),
    .o(_al_u8287_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u8288 (
    .a(_al_u8285_o),
    .b(_al_u8287_o),
    .c(unsign),
    .o(_al_u8288_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8289 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[46]),
    .o(_al_u8289_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8290 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8288_o),
    .d(_al_u8289_o),
    .o(_al_u8290_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8291 (
    .a(uncache_data[62]),
    .b(uncache_data[46]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8291_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u8292 (
    .a(_al_u8291_o),
    .b(uncache_data[54]),
    .c(\exu/lsu/n2_lutinv ),
    .d(unsign),
    .o(\exu/lsu/n59 [46]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8293 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [46]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8293_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8294 (
    .a(\exu/alu_au/add_64 [46]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [46]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8295 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3609_o),
    .c(\exu/alu_au/n31 [46]),
    .d(rd_data_add),
    .o(_al_u8295_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8296 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[46]),
    .o(_al_u8296_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8297 (
    .a(_al_u8296_o),
    .b(rd_data_xor),
    .c(ds1[46]),
    .d(ds2[46]),
    .o(_al_u8297_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8298 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[46]),
    .d(ds2[46]),
    .o(\exu/alu_au/n33 [46]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8299 (
    .a(_al_u8295_o),
    .b(_al_u8297_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [46]),
    .o(_al_u8299_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8300 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[46]),
    .c(data_rd[47]),
    .o(\exu/n57 [46]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8301 (
    .a(data_rd[45]),
    .b(data_rd[46]),
    .c(ex_size[2]),
    .o(_al_u8301_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8302 (
    .a(\exu/n57 [46]),
    .b(_al_u2855_o),
    .c(_al_u8301_o),
    .d(shift_l),
    .o(_al_u8302_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8303 (
    .a(_al_u8290_o),
    .b(_al_u8293_o),
    .c(_al_u8299_o),
    .d(_al_u8302_o),
    .o(\exu/n64 [46]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u8304 (
    .a(_al_u8027_o),
    .b(_al_u8028_o),
    .c(\exu/lsu/n5_lutinv ),
    .o(_al_u8304_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8305 (
    .a(_al_u8164_o),
    .b(\exu/lsu/n2_lutinv ),
    .o(_al_u8305_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8306 (
    .a(\biu/l1d_out [45]),
    .b(uncache_data[45]),
    .c(_al_u3224_o),
    .o(_al_u8306_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u8307 (
    .a(_al_u8306_o),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .c(\exu/n60_lutinv ),
    .o(_al_u8307_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*~A)))"),
    .INIT(16'h10f0))
    _al_u8308 (
    .a(_al_u8304_o),
    .b(_al_u8305_o),
    .c(_al_u8307_o),
    .d(unsign),
    .o(_al_u8308_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8309 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[45]),
    .o(_al_u8309_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8310 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8308_o),
    .d(_al_u8309_o),
    .o(_al_u8310_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8311 (
    .a(uncache_data[61]),
    .b(uncache_data[45]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8311_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u8312 (
    .a(_al_u8311_o),
    .b(uncache_data[53]),
    .c(\exu/lsu/n2_lutinv ),
    .d(unsign),
    .o(\exu/lsu/n59 [45]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8313 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [45]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8313_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8314 (
    .a(\exu/alu_au/add_64 [45]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [45]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8315 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3617_o),
    .c(\exu/alu_au/n31 [45]),
    .d(rd_data_add),
    .o(_al_u8315_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8316 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[45]),
    .o(_al_u8316_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8317 (
    .a(_al_u8316_o),
    .b(rd_data_xor),
    .c(ds1[45]),
    .d(ds2[45]),
    .o(_al_u8317_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8318 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[45]),
    .d(ds2[45]),
    .o(\exu/alu_au/n33 [45]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8319 (
    .a(_al_u8315_o),
    .b(_al_u8317_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [45]),
    .o(_al_u8319_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8320 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[45]),
    .c(data_rd[46]),
    .o(\exu/n57 [45]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8321 (
    .a(data_rd[44]),
    .b(data_rd[45]),
    .c(ex_size[2]),
    .o(_al_u8321_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8322 (
    .a(\exu/n57 [45]),
    .b(_al_u2855_o),
    .c(_al_u8321_o),
    .d(shift_l),
    .o(_al_u8322_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8323 (
    .a(_al_u8310_o),
    .b(_al_u8313_o),
    .c(_al_u8319_o),
    .d(_al_u8322_o),
    .o(\exu/n64 [45]));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8324 (
    .a(\biu/l1d_out [60]),
    .b(uncache_data[60]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u8324_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(C*A)))"),
    .INIT(16'hec00))
    _al_u8325 (
    .a(_al_u8180_o),
    .b(_al_u8324_o),
    .c(\exu/lsu/n2_lutinv ),
    .d(unsign),
    .o(_al_u8325_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8326 (
    .a(uncache_data[44]),
    .b(_al_u3224_o),
    .o(_al_u8326_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8327 (
    .a(\biu/l1d_out [44]),
    .b(_al_u3224_o),
    .c(_al_u8326_o),
    .o(_al_u8327_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u8328 (
    .a(_al_u8325_o),
    .b(_al_u8327_o),
    .c(\exu/lsu/mux27_b56_sel_is_3_o ),
    .d(\exu/n60_lutinv ),
    .o(_al_u8328_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8329 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[44]),
    .o(_al_u8329_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8330 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8328_o),
    .d(_al_u8329_o),
    .o(_al_u8330_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8331 (
    .a(uncache_data[60]),
    .b(uncache_data[44]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8331_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u8332 (
    .a(_al_u8331_o),
    .b(uncache_data[52]),
    .c(\exu/lsu/n2_lutinv ),
    .d(unsign),
    .o(\exu/lsu/n59 [44]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8333 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [44]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8333_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8334 (
    .a(\exu/alu_au/add_64 [44]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [44]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8335 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3625_o),
    .c(\exu/alu_au/n31 [44]),
    .d(rd_data_add),
    .o(_al_u8335_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8336 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[44]),
    .o(_al_u8336_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8337 (
    .a(_al_u8336_o),
    .b(rd_data_xor),
    .c(ds1[44]),
    .d(ds2[44]),
    .o(_al_u8337_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8338 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[44]),
    .d(ds2[44]),
    .o(\exu/alu_au/n33 [44]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8339 (
    .a(_al_u8335_o),
    .b(_al_u8337_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [44]),
    .o(_al_u8339_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8340 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[44]),
    .c(data_rd[45]),
    .o(\exu/n57 [44]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8341 (
    .a(data_rd[43]),
    .b(data_rd[44]),
    .c(ex_size[2]),
    .o(_al_u8341_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8342 (
    .a(\exu/n57 [44]),
    .b(_al_u2855_o),
    .c(_al_u8341_o),
    .d(shift_l),
    .o(_al_u8342_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8343 (
    .a(_al_u8330_o),
    .b(_al_u8333_o),
    .c(_al_u8339_o),
    .d(_al_u8342_o),
    .o(\exu/n64 [44]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfa3f))
    _al_u8344 (
    .a(_al_u8061_o),
    .b(_al_u8198_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8344_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8345 (
    .a(uncache_data[43]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [43]),
    .o(_al_u8345_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8346 (
    .a(_al_u8345_o),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .c(\exu/n60_lutinv ),
    .o(_al_u8346_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u8347 (
    .a(_al_u8344_o),
    .b(_al_u8346_o),
    .c(unsign),
    .o(_al_u8347_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8348 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[43]),
    .o(_al_u8348_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8349 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8347_o),
    .d(_al_u8348_o),
    .o(_al_u8349_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8350 (
    .a(uncache_data[59]),
    .b(uncache_data[43]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8350_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u8351 (
    .a(_al_u8350_o),
    .b(uncache_data[51]),
    .c(\exu/lsu/n2_lutinv ),
    .d(unsign),
    .o(\exu/lsu/n59 [43]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8352 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [43]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8352_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8353 (
    .a(\exu/alu_au/add_64 [43]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [43]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8354 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3633_o),
    .c(\exu/alu_au/n31 [43]),
    .d(rd_data_add),
    .o(_al_u8354_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8355 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[43]),
    .o(_al_u8355_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8356 (
    .a(_al_u8355_o),
    .b(rd_data_xor),
    .c(ds1[43]),
    .d(ds2[43]),
    .o(_al_u8356_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8357 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[43]),
    .d(ds2[43]),
    .o(\exu/alu_au/n33 [43]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8358 (
    .a(_al_u8354_o),
    .b(_al_u8356_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [43]),
    .o(_al_u8358_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8359 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[43]),
    .c(data_rd[44]),
    .o(\exu/n57 [43]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8360 (
    .a(data_rd[42]),
    .b(data_rd[43]),
    .c(ex_size[2]),
    .o(_al_u8360_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8361 (
    .a(\exu/n57 [43]),
    .b(_al_u2855_o),
    .c(_al_u8360_o),
    .d(shift_l),
    .o(_al_u8361_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8362 (
    .a(_al_u8349_o),
    .b(_al_u8352_o),
    .c(_al_u8358_o),
    .d(_al_u8361_o),
    .o(\exu/n64 [43]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfacf))
    _al_u8363 (
    .a(_al_u8077_o),
    .b(_al_u8215_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8363_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8364 (
    .a(uncache_data[42]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [42]),
    .o(_al_u8364_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8365 (
    .a(_al_u8364_o),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .c(\exu/n60_lutinv ),
    .o(_al_u8365_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u8366 (
    .a(_al_u8363_o),
    .b(_al_u8365_o),
    .c(unsign),
    .o(_al_u8366_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8367 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[42]),
    .o(_al_u8367_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8368 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8366_o),
    .d(_al_u8367_o),
    .o(_al_u8368_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8369 (
    .a(uncache_data[58]),
    .b(uncache_data[42]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8369_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u8370 (
    .a(_al_u8369_o),
    .b(uncache_data[50]),
    .c(\exu/lsu/n2_lutinv ),
    .d(unsign),
    .o(\exu/lsu/n59 [42]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8371 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [42]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8371_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8372 (
    .a(\exu/alu_au/add_64 [42]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [42]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8373 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3641_o),
    .c(\exu/alu_au/n31 [42]),
    .d(rd_data_add),
    .o(_al_u8373_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8374 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[42]),
    .o(_al_u8374_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8375 (
    .a(_al_u8374_o),
    .b(rd_data_xor),
    .c(ds1[42]),
    .d(ds2[42]),
    .o(_al_u8375_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8376 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[42]),
    .d(ds2[42]),
    .o(\exu/alu_au/n33 [42]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8377 (
    .a(_al_u8373_o),
    .b(_al_u8375_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [42]),
    .o(_al_u8377_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8378 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[42]),
    .c(data_rd[43]),
    .o(\exu/n57 [42]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8379 (
    .a(data_rd[41]),
    .b(data_rd[42]),
    .c(ex_size[2]),
    .o(_al_u8379_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8380 (
    .a(\exu/n57 [42]),
    .b(_al_u2855_o),
    .c(_al_u8379_o),
    .d(shift_l),
    .o(_al_u8380_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8381 (
    .a(_al_u8368_o),
    .b(_al_u8371_o),
    .c(_al_u8377_o),
    .d(_al_u8380_o),
    .o(\exu/n64 [42]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf5cf))
    _al_u8382 (
    .a(_al_u8093_o),
    .b(_al_u8232_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8382_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u8383 (
    .a(\biu/l1d_out [41]),
    .b(_al_u3224_o),
    .c(uncache_data[41]),
    .o(_al_u8383_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u8384 (
    .a(_al_u8383_o),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .c(\exu/n60_lutinv ),
    .o(_al_u8384_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u8385 (
    .a(_al_u8382_o),
    .b(_al_u8384_o),
    .c(unsign),
    .o(_al_u8385_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8386 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[41]),
    .o(_al_u8386_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8387 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8385_o),
    .d(_al_u8386_o),
    .o(_al_u8387_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8388 (
    .a(uncache_data[57]),
    .b(uncache_data[41]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8388_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u8389 (
    .a(_al_u8388_o),
    .b(uncache_data[49]),
    .c(\exu/lsu/n2_lutinv ),
    .d(unsign),
    .o(\exu/lsu/n59 [41]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8390 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [41]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8390_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'h00e4))
    _al_u8391 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[41]),
    .c(data_rd[42]),
    .d(shift_l),
    .o(_al_u8391_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8392 (
    .a(data_rd[40]),
    .b(data_rd[41]),
    .c(ex_size[2]),
    .d(shift_l),
    .o(_al_u8392_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u8393 (
    .a(_al_u8391_o),
    .b(_al_u2855_o),
    .c(_al_u8392_o),
    .o(_al_u8393_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8394 (
    .a(\exu/alu_au/add_64 [41]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [41]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8395 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3649_o),
    .c(\exu/alu_au/n31 [41]),
    .d(rd_data_add),
    .o(_al_u8395_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8396 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[41]),
    .o(_al_u8396_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8397 (
    .a(_al_u8396_o),
    .b(rd_data_xor),
    .c(ds1[41]),
    .d(ds2[41]),
    .o(_al_u8397_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8398 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[41]),
    .d(ds2[41]),
    .o(\exu/alu_au/n33 [41]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8399 (
    .a(_al_u8395_o),
    .b(_al_u8397_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [41]),
    .o(_al_u8399_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B*~A)))"),
    .INIT(16'hfbf0))
    _al_u8400 (
    .a(_al_u8387_o),
    .b(_al_u8390_o),
    .c(_al_u8393_o),
    .d(_al_u8399_o),
    .o(\exu/n64 [41]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfa3f))
    _al_u8401 (
    .a(_al_u8109_o),
    .b(_al_u8249_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8401_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8402 (
    .a(uncache_data[40]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [40]),
    .o(_al_u8402_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8403 (
    .a(_al_u8402_o),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .c(\exu/n60_lutinv ),
    .o(_al_u8403_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u8404 (
    .a(_al_u8401_o),
    .b(_al_u8403_o),
    .c(unsign),
    .o(_al_u8404_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8405 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[40]),
    .o(_al_u8405_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8406 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8404_o),
    .d(_al_u8405_o),
    .o(_al_u8406_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8407 (
    .a(uncache_data[56]),
    .b(uncache_data[40]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8407_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u8408 (
    .a(_al_u8407_o),
    .b(uncache_data[48]),
    .c(\exu/lsu/n2_lutinv ),
    .d(unsign),
    .o(\exu/lsu/n59 [40]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8409 (
    .a(_al_u7995_o),
    .b(\exu/lsu/n59 [40]),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8409_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'h00e4))
    _al_u8410 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[40]),
    .c(data_rd[41]),
    .d(shift_l),
    .o(_al_u8410_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8411 (
    .a(data_rd[39]),
    .b(data_rd[40]),
    .c(ex_size[2]),
    .d(shift_l),
    .o(_al_u8411_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u8412 (
    .a(_al_u8410_o),
    .b(_al_u2855_o),
    .c(_al_u8411_o),
    .o(_al_u8412_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8413 (
    .a(\exu/alu_au/add_64 [40]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [40]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8414 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3657_o),
    .c(\exu/alu_au/n31 [40]),
    .d(rd_data_add),
    .o(_al_u8414_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8415 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[40]),
    .o(_al_u8415_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8416 (
    .a(_al_u8415_o),
    .b(rd_data_xor),
    .c(ds1[40]),
    .d(ds2[40]),
    .o(_al_u8416_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8417 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[40]),
    .d(ds2[40]),
    .o(\exu/alu_au/n33 [40]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8418 (
    .a(_al_u8414_o),
    .b(_al_u8416_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [40]),
    .o(_al_u8418_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B*~A)))"),
    .INIT(16'hfbf0))
    _al_u8419 (
    .a(_al_u8406_o),
    .b(_al_u8409_o),
    .c(_al_u8412_o),
    .d(_al_u8418_o),
    .o(\exu/n64 [40]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~(~B*A)))"),
    .INIT(16'hf200))
    _al_u8420 (
    .a(\biu/l1d_out [47]),
    .b(_al_u3224_o),
    .c(_al_u7974_o),
    .d(\exu/lsu/n2_lutinv ),
    .o(_al_u8420_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(~B*~A))"),
    .INIT(16'h0e00))
    _al_u8421 (
    .a(\biu/l1d_out [63]),
    .b(_al_u3224_o),
    .c(_al_u7981_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u8421_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8422 (
    .a(\biu/l1d_out [55]),
    .b(uncache_data[55]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u8422_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8423 (
    .a(\biu/l1d_out [39]),
    .b(uncache_data[39]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n0_lutinv ),
    .o(_al_u8423_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u8424 (
    .a(_al_u8420_o),
    .b(_al_u8421_o),
    .c(_al_u8422_o),
    .d(_al_u8423_o),
    .o(_al_u8424_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~A)*~(B)*~(D)+~(C*~A)*B*~(D)+~(~(C*~A))*B*D+~(C*~A)*B*D)"),
    .INIT(16'hccaf))
    _al_u8425 (
    .a(_al_u7979_o),
    .b(_al_u8424_o),
    .c(ex_size[2]),
    .d(unsign),
    .o(_al_u8425_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8426 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[39]),
    .o(_al_u8426_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u8427 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8425_o),
    .d(_al_u8426_o),
    .o(_al_u8427_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8428 (
    .a(uncache_data[63]),
    .b(uncache_data[47]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8428_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8429 (
    .a(uncache_data[55]),
    .b(uncache_data[39]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8429_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u8430 (
    .a(_al_u7995_o),
    .b(_al_u8428_o),
    .c(_al_u8429_o),
    .d(unsign),
    .o(_al_u8430_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8431 (
    .a(_al_u8430_o),
    .b(\exu/c_stb_lutinv ),
    .c(\exu/n59_lutinv ),
    .o(_al_u8431_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'h00e4))
    _al_u8432 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[39]),
    .c(data_rd[40]),
    .d(shift_l),
    .o(_al_u8432_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8433 (
    .a(data_rd[38]),
    .b(data_rd[39]),
    .c(ex_size[2]),
    .d(shift_l),
    .o(_al_u8433_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u8434 (
    .a(_al_u8432_o),
    .b(_al_u2855_o),
    .c(_al_u8433_o),
    .o(_al_u8434_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8435 (
    .a(\exu/alu_au/add_64 [39]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [39]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8436 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3672_o),
    .c(\exu/alu_au/n31 [39]),
    .d(rd_data_add),
    .o(_al_u8436_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8437 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[39]),
    .o(_al_u8437_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8438 (
    .a(_al_u8437_o),
    .b(rd_data_xor),
    .c(ds1[39]),
    .d(ds2[39]),
    .o(_al_u8438_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8439 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[39]),
    .d(ds2[39]),
    .o(\exu/alu_au/n33 [39]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8440 (
    .a(_al_u8436_o),
    .b(_al_u8438_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [39]),
    .o(_al_u8440_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B*~A)))"),
    .INIT(16'hfbf0))
    _al_u8441 (
    .a(_al_u8427_o),
    .b(_al_u8431_o),
    .c(_al_u8434_o),
    .d(_al_u8440_o),
    .o(\exu/n64 [39]));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'ha300))
    _al_u8442 (
    .a(_al_u8011_o),
    .b(_al_u8146_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8442_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8443 (
    .a(_al_u8286_o),
    .b(_al_u8127_o),
    .o(_al_u8443_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u8444 (
    .a(uncache_data[38]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [38]),
    .o(_al_u8444_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u8445 (
    .a(_al_u8444_o),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .c(\exu/n60_lutinv ),
    .o(_al_u8445_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*A))"),
    .INIT(16'h1030))
    _al_u8446 (
    .a(_al_u8442_o),
    .b(_al_u8443_o),
    .c(_al_u8445_o),
    .d(unsign),
    .o(_al_u8446_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8447 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[38]),
    .o(_al_u8447_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8448 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8446_o),
    .d(_al_u8447_o),
    .o(_al_u8448_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8449 (
    .a(uncache_data[62]),
    .b(uncache_data[38]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8449_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8450 (
    .a(uncache_data[54]),
    .b(uncache_data[46]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8450_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u8451 (
    .a(_al_u7995_o),
    .b(_al_u8449_o),
    .c(_al_u8450_o),
    .d(unsign),
    .o(_al_u8451_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8452 (
    .a(_al_u8451_o),
    .b(\exu/c_stb_lutinv ),
    .c(\exu/n59_lutinv ),
    .o(_al_u8452_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8453 (
    .a(\exu/alu_au/add_64 [38]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [38]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8454 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3680_o),
    .c(\exu/alu_au/n31 [38]),
    .d(rd_data_add),
    .o(_al_u8454_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8455 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[38]),
    .o(_al_u8455_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8456 (
    .a(_al_u8455_o),
    .b(rd_data_xor),
    .c(ds1[38]),
    .d(ds2[38]),
    .o(_al_u8456_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8457 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[38]),
    .d(ds2[38]),
    .o(\exu/alu_au/n33 [38]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8458 (
    .a(_al_u8454_o),
    .b(_al_u8456_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [38]),
    .o(_al_u8458_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u8459 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[38]),
    .c(data_rd[39]),
    .o(_al_u8459_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8460 (
    .a(data_rd[37]),
    .b(data_rd[38]),
    .c(ex_size[2]),
    .o(_al_u8460_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    .INIT(16'h0c44))
    _al_u8461 (
    .a(_al_u8459_o),
    .b(_al_u2855_o),
    .c(_al_u8460_o),
    .d(shift_l),
    .o(_al_u8461_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8462 (
    .a(_al_u8448_o),
    .b(_al_u8452_o),
    .c(_al_u8458_o),
    .d(_al_u8461_o),
    .o(\exu/n64 [38]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(~B*~A))"),
    .INIT(16'h0e00))
    _al_u8463 (
    .a(\biu/l1d_out [61]),
    .b(_al_u3224_o),
    .c(_al_u8028_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u8463_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(~B*~A))"),
    .INIT(16'h0e00))
    _al_u8464 (
    .a(\biu/l1d_out [53]),
    .b(_al_u3224_o),
    .c(_al_u8163_o),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u8464_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8465 (
    .a(\biu/l1d_out [45]),
    .b(uncache_data[45]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n2_lutinv ),
    .o(_al_u8465_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8466 (
    .a(\biu/l1d_out [37]),
    .b(uncache_data[37]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n0_lutinv ),
    .o(_al_u8466_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u8467 (
    .a(_al_u8463_o),
    .b(_al_u8464_o),
    .c(_al_u8465_o),
    .d(_al_u8466_o),
    .o(_al_u8467_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~A)*~(B)*~(D)+~(C*~A)*B*~(D)+~(~(C*~A))*B*D+~(C*~A)*B*D)"),
    .INIT(16'hccaf))
    _al_u8468 (
    .a(_al_u7979_o),
    .b(_al_u8467_o),
    .c(ex_size[2]),
    .d(unsign),
    .o(_al_u8468_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8469 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[37]),
    .o(_al_u8469_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u8470 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8468_o),
    .d(_al_u8469_o),
    .o(_al_u8470_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8471 (
    .a(uncache_data[53]),
    .b(uncache_data[45]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8471_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8472 (
    .a(uncache_data[61]),
    .b(uncache_data[37]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8472_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u8473 (
    .a(_al_u7995_o),
    .b(_al_u8471_o),
    .c(_al_u8472_o),
    .d(unsign),
    .o(_al_u8473_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8474 (
    .a(_al_u8473_o),
    .b(\exu/c_stb_lutinv ),
    .c(\exu/n59_lutinv ),
    .o(_al_u8474_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8475 (
    .a(\exu/alu_au/add_64 [37]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [37]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8476 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3688_o),
    .c(\exu/alu_au/n31 [37]),
    .d(rd_data_add),
    .o(_al_u8476_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8477 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[37]),
    .o(_al_u8477_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8478 (
    .a(_al_u8477_o),
    .b(rd_data_xor),
    .c(ds1[37]),
    .d(ds2[37]),
    .o(_al_u8478_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8479 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[37]),
    .d(ds2[37]),
    .o(\exu/alu_au/n33 [37]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8480 (
    .a(_al_u8476_o),
    .b(_al_u8478_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [37]),
    .o(_al_u8480_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u8481 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[37]),
    .c(data_rd[38]),
    .o(_al_u8481_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8482 (
    .a(data_rd[36]),
    .b(data_rd[37]),
    .c(ex_size[2]),
    .o(_al_u8482_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    .INIT(16'h0c44))
    _al_u8483 (
    .a(_al_u8481_o),
    .b(_al_u2855_o),
    .c(_al_u8482_o),
    .d(shift_l),
    .o(_al_u8483_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8484 (
    .a(_al_u8470_o),
    .b(_al_u8474_o),
    .c(_al_u8480_o),
    .d(_al_u8483_o),
    .o(\exu/n64 [37]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(~B*~A))"),
    .INIT(16'h0e00))
    _al_u8485 (
    .a(\biu/l1d_out [44]),
    .b(_al_u3224_o),
    .c(_al_u8326_o),
    .d(\exu/lsu/n2_lutinv ),
    .o(_al_u8485_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8486 (
    .a(\biu/l1d_out [60]),
    .b(uncache_data[60]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u8486_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8487 (
    .a(\biu/l1d_out [52]),
    .b(uncache_data[52]),
    .c(_al_u3224_o),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u8487_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8488 (
    .a(uncache_data[36]),
    .b(_al_u3224_o),
    .o(_al_u8488_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~(~B*A)))"),
    .INIT(16'hf200))
    _al_u8489 (
    .a(\biu/l1d_out [36]),
    .b(_al_u3224_o),
    .c(_al_u8488_o),
    .d(\exu/lsu/n0_lutinv ),
    .o(_al_u8489_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u8490 (
    .a(_al_u8485_o),
    .b(_al_u8486_o),
    .c(_al_u8487_o),
    .d(_al_u8489_o),
    .o(_al_u8490_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~A)*~(B)*~(D)+~(C*~A)*B*~(D)+~(~(C*~A))*B*D+~(C*~A)*B*D)"),
    .INIT(16'hccaf))
    _al_u8491 (
    .a(_al_u7979_o),
    .b(_al_u8490_o),
    .c(ex_size[2]),
    .d(unsign),
    .o(_al_u8491_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8492 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[36]),
    .o(_al_u8492_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u8493 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8491_o),
    .d(_al_u8492_o),
    .o(_al_u8493_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8494 (
    .a(uncache_data[52]),
    .b(uncache_data[44]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8494_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8495 (
    .a(uncache_data[60]),
    .b(uncache_data[36]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8495_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u8496 (
    .a(_al_u7995_o),
    .b(_al_u8494_o),
    .c(_al_u8495_o),
    .d(unsign),
    .o(_al_u8496_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8497 (
    .a(_al_u8496_o),
    .b(\exu/c_stb_lutinv ),
    .c(\exu/n59_lutinv ),
    .o(_al_u8497_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8498 (
    .a(\exu/alu_au/add_64 [36]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [36]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8499 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3696_o),
    .c(\exu/alu_au/n31 [36]),
    .d(rd_data_add),
    .o(_al_u8499_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8500 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[36]),
    .o(_al_u8500_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8501 (
    .a(_al_u8500_o),
    .b(rd_data_xor),
    .c(ds1[36]),
    .d(ds2[36]),
    .o(_al_u8501_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8502 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[36]),
    .d(ds2[36]),
    .o(\exu/alu_au/n33 [36]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8503 (
    .a(_al_u8499_o),
    .b(_al_u8501_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [36]),
    .o(_al_u8503_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8504 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[36]),
    .c(data_rd[37]),
    .o(\exu/n57 [36]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8505 (
    .a(data_rd[35]),
    .b(data_rd[36]),
    .c(ex_size[2]),
    .o(_al_u8505_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8506 (
    .a(\exu/n57 [36]),
    .b(_al_u2855_o),
    .c(_al_u8505_o),
    .d(shift_l),
    .o(_al_u8506_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8507 (
    .a(_al_u8493_o),
    .b(_al_u8497_o),
    .c(_al_u8503_o),
    .d(_al_u8506_o),
    .o(\exu/n64 [36]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u8508 (
    .a(\biu/l1d_out [35]),
    .b(_al_u3224_o),
    .c(uncache_data[35]),
    .o(_al_u8508_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8509 (
    .a(_al_u8508_o),
    .b(\exu/lsu/n0_lutinv ),
    .o(_al_u8509_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h5c00))
    _al_u8510 (
    .a(_al_u8061_o),
    .b(_al_u8198_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8510_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8511 (
    .a(_al_u8345_o),
    .b(_al_u8127_o),
    .c(\exu/n60_lutinv ),
    .o(_al_u8511_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*~A)))"),
    .INIT(16'h10f0))
    _al_u8512 (
    .a(_al_u8509_o),
    .b(_al_u8510_o),
    .c(_al_u8511_o),
    .d(unsign),
    .o(_al_u8512_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8513 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[35]),
    .o(_al_u8513_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8514 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8512_o),
    .d(_al_u8513_o),
    .o(_al_u8514_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8515 (
    .a(uncache_data[51]),
    .b(uncache_data[43]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8515_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8516 (
    .a(uncache_data[59]),
    .b(uncache_data[35]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8516_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u8517 (
    .a(_al_u7995_o),
    .b(_al_u8515_o),
    .c(_al_u8516_o),
    .d(unsign),
    .o(_al_u8517_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8518 (
    .a(_al_u8517_o),
    .b(\exu/c_stb_lutinv ),
    .c(\exu/n59_lutinv ),
    .o(_al_u8518_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'h00e4))
    _al_u8519 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[35]),
    .c(data_rd[36]),
    .d(shift_l),
    .o(_al_u8519_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8520 (
    .a(data_rd[34]),
    .b(data_rd[35]),
    .c(ex_size[2]),
    .d(shift_l),
    .o(_al_u8520_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u8521 (
    .a(_al_u8519_o),
    .b(_al_u2855_o),
    .c(_al_u8520_o),
    .o(_al_u8521_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8522 (
    .a(\exu/alu_au/add_64 [35]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [35]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8523 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3704_o),
    .c(\exu/alu_au/n31 [35]),
    .d(rd_data_add),
    .o(_al_u8523_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8524 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[35]),
    .o(_al_u8524_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8525 (
    .a(_al_u8524_o),
    .b(rd_data_xor),
    .c(ds1[35]),
    .d(ds2[35]),
    .o(_al_u8525_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8526 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[35]),
    .d(ds2[35]),
    .o(\exu/alu_au/n33 [35]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8527 (
    .a(_al_u8523_o),
    .b(_al_u8525_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [35]),
    .o(_al_u8527_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B*~A)))"),
    .INIT(16'hfbf0))
    _al_u8528 (
    .a(_al_u8514_o),
    .b(_al_u8518_o),
    .c(_al_u8521_o),
    .d(_al_u8527_o),
    .o(\exu/n64 [35]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h5300))
    _al_u8529 (
    .a(_al_u8077_o),
    .b(_al_u8215_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8529_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8530 (
    .a(_al_u8364_o),
    .b(_al_u8127_o),
    .o(_al_u8530_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u8531 (
    .a(uncache_data[34]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [34]),
    .o(_al_u8531_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u8532 (
    .a(_al_u8531_o),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .c(\exu/n60_lutinv ),
    .o(_al_u8532_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*A))"),
    .INIT(16'h1030))
    _al_u8533 (
    .a(_al_u8529_o),
    .b(_al_u8530_o),
    .c(_al_u8532_o),
    .d(unsign),
    .o(_al_u8533_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8534 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[34]),
    .o(_al_u8534_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8535 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8533_o),
    .d(_al_u8534_o),
    .o(_al_u8535_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8536 (
    .a(uncache_data[50]),
    .b(uncache_data[34]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8536_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8537 (
    .a(uncache_data[58]),
    .b(uncache_data[42]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8537_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u8538 (
    .a(_al_u7995_o),
    .b(_al_u8536_o),
    .c(_al_u8537_o),
    .d(unsign),
    .o(_al_u8538_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8539 (
    .a(_al_u8538_o),
    .b(\exu/c_stb_lutinv ),
    .c(\exu/n59_lutinv ),
    .o(_al_u8539_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .INIT(16'h00e4))
    _al_u8540 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[34]),
    .c(data_rd[35]),
    .d(shift_l),
    .o(_al_u8540_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8541 (
    .a(data_rd[33]),
    .b(data_rd[34]),
    .c(ex_size[2]),
    .d(shift_l),
    .o(_al_u8541_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u8542 (
    .a(_al_u8540_o),
    .b(_al_u2855_o),
    .c(_al_u8541_o),
    .o(_al_u8542_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8543 (
    .a(\exu/alu_au/add_64 [34]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [34]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8544 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3712_o),
    .c(\exu/alu_au/n31 [34]),
    .d(rd_data_add),
    .o(_al_u8544_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8545 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[34]),
    .o(_al_u8545_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8546 (
    .a(_al_u8545_o),
    .b(rd_data_xor),
    .c(ds1[34]),
    .d(ds2[34]),
    .o(_al_u8546_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8547 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[34]),
    .d(ds2[34]),
    .o(\exu/alu_au/n33 [34]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8548 (
    .a(_al_u8544_o),
    .b(_al_u8546_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [34]),
    .o(_al_u8548_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B*~A)))"),
    .INIT(16'hfbf0))
    _al_u8549 (
    .a(_al_u8535_o),
    .b(_al_u8539_o),
    .c(_al_u8542_o),
    .d(_al_u8548_o),
    .o(\exu/n64 [34]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8550 (
    .a(_al_u8383_o),
    .b(\exu/lsu/n2_lutinv ),
    .o(_al_u8550_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'ha300))
    _al_u8551 (
    .a(_al_u8093_o),
    .b(_al_u8232_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8551_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8552 (
    .a(_al_u7906_o),
    .b(\exu/lsu/mux27_b56_sel_is_3_o ),
    .c(\exu/n60_lutinv ),
    .o(_al_u8552_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*~A)))"),
    .INIT(16'h10f0))
    _al_u8553 (
    .a(_al_u8550_o),
    .b(_al_u8551_o),
    .c(_al_u8552_o),
    .d(unsign),
    .o(_al_u8553_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8554 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[33]),
    .o(_al_u8554_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8555 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8553_o),
    .d(_al_u8554_o),
    .o(_al_u8555_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8556 (
    .a(uncache_data[49]),
    .b(uncache_data[41]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8556_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8557 (
    .a(uncache_data[57]),
    .b(uncache_data[33]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8557_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u8558 (
    .a(_al_u7995_o),
    .b(_al_u8556_o),
    .c(_al_u8557_o),
    .d(unsign),
    .o(_al_u8558_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8559 (
    .a(_al_u8558_o),
    .b(\exu/c_stb_lutinv ),
    .c(\exu/n59_lutinv ),
    .o(_al_u8559_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8560 (
    .a(\exu/alu_au/add_64 [33]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [33]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8561 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3720_o),
    .c(\exu/alu_au/n31 [33]),
    .d(rd_data_add),
    .o(_al_u8561_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8562 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[33]),
    .o(_al_u8562_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8563 (
    .a(_al_u8562_o),
    .b(rd_data_xor),
    .c(ds1[33]),
    .d(ds2[33]),
    .o(_al_u8563_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8564 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[33]),
    .d(ds2[33]),
    .o(\exu/alu_au/n33 [33]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8565 (
    .a(_al_u8561_o),
    .b(_al_u8563_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [33]),
    .o(_al_u8565_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8566 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[33]),
    .c(data_rd[34]),
    .o(\exu/n57 [33]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8567 (
    .a(data_rd[32]),
    .b(data_rd[33]),
    .c(ex_size[2]),
    .o(_al_u8567_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'h0c88))
    _al_u8568 (
    .a(\exu/n57 [33]),
    .b(_al_u2855_o),
    .c(_al_u8567_o),
    .d(shift_l),
    .o(_al_u8568_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8569 (
    .a(_al_u8555_o),
    .b(_al_u8559_o),
    .c(_al_u8565_o),
    .d(_al_u8568_o),
    .o(\exu/n64 [33]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u8570 (
    .a(_al_u7936_o),
    .b(\exu/lsu/n0_lutinv ),
    .o(_al_u8570_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h5c00))
    _al_u8571 (
    .a(_al_u8109_o),
    .b(_al_u8249_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8571_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8572 (
    .a(_al_u8402_o),
    .b(_al_u8127_o),
    .c(\exu/n60_lutinv ),
    .o(_al_u8572_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*~A)))"),
    .INIT(16'h10f0))
    _al_u8573 (
    .a(_al_u8570_o),
    .b(_al_u8571_o),
    .c(_al_u8572_o),
    .d(unsign),
    .o(_al_u8573_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8574 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[32]),
    .o(_al_u8574_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*~A))"),
    .INIT(16'hbf00))
    _al_u8575 (
    .a(_al_u8125_o),
    .b(_al_u8126_o),
    .c(_al_u8573_o),
    .d(_al_u8574_o),
    .o(_al_u8575_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8576 (
    .a(uncache_data[48]),
    .b(uncache_data[40]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8576_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8577 (
    .a(uncache_data[56]),
    .b(uncache_data[32]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8577_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u8578 (
    .a(_al_u7995_o),
    .b(_al_u8576_o),
    .c(_al_u8577_o),
    .d(unsign),
    .o(_al_u8578_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8579 (
    .a(_al_u8578_o),
    .b(\exu/c_stb_lutinv ),
    .c(\exu/n59_lutinv ),
    .o(_al_u8579_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8580 (
    .a(\exu/alu_au/add_64 [32]),
    .b(\exu/alu_au/sub_64 [31]),
    .c(rd_data_sub),
    .d(ex_size[2]),
    .o(\exu/alu_au/n31 [32]));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u8581 (
    .a(\exu/c_stb_lutinv ),
    .b(_al_u3728_o),
    .c(\exu/alu_au/n31 [32]),
    .d(rd_data_add),
    .o(_al_u8581_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u8582 (
    .a(rd_data_ds1),
    .b(rd_data_or),
    .c(ds1[32]),
    .o(_al_u8582_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5dd0))
    _al_u8583 (
    .a(_al_u8582_o),
    .b(rd_data_xor),
    .c(ds1[32]),
    .d(ds2[32]),
    .o(_al_u8583_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8584 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[32]),
    .d(ds2[32]),
    .o(\exu/alu_au/n33 [32]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u8585 (
    .a(_al_u8581_o),
    .b(_al_u8583_o),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [32]),
    .o(_al_u8585_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u8586 (
    .a(\exu/mux27_b32_sel_is_1_o ),
    .b(data_rd[32]),
    .c(data_rd[33]),
    .o(\exu/n57 [32]));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u8587 (
    .a(data_rd[31]),
    .b(data_rd[32]),
    .c(ex_size[2]),
    .d(shift_l),
    .o(_al_u8587_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(~D*A)))"),
    .INIT(16'hc0c8))
    _al_u8588 (
    .a(\exu/n57 [32]),
    .b(_al_u2855_o),
    .c(_al_u8587_o),
    .d(shift_l),
    .o(_al_u8588_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8589 (
    .a(_al_u8575_o),
    .b(_al_u8579_o),
    .c(_al_u8585_o),
    .d(_al_u8588_o),
    .o(\exu/n64 [32]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u8590 (
    .a(_al_u7979_o),
    .b(_al_u7912_o),
    .o(_al_u8590_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8591 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[31]),
    .o(_al_u8591_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8592 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8590_o),
    .d(_al_u8591_o),
    .o(_al_u8592_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u8593 (
    .a(_al_u7991_o),
    .b(_al_u7994_o),
    .c(_al_u7912_o),
    .o(_al_u8593_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8594 (
    .a(_al_u8593_o),
    .b(\exu/c_stb_lutinv ),
    .c(\exu/n59_lutinv ),
    .o(_al_u8594_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8595 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[31]),
    .d(ds2[31]),
    .o(_al_u8595_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8596 (
    .a(\exu/alu_au/sub_64 [31]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[31]),
    .o(_al_u8596_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8597 (
    .a(_al_u8595_o),
    .b(_al_u8596_o),
    .c(\exu/alu_au/add_64 [31]),
    .d(rd_data_add),
    .o(_al_u8597_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8598 (
    .a(_al_u8597_o),
    .b(rd_data_xor),
    .c(ds1[31]),
    .d(ds2[31]),
    .o(_al_u8598_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8599 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[31]),
    .d(ds2[31]),
    .o(\exu/alu_au/n33 [31]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8600 (
    .a(_al_u8598_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [31]),
    .o(_al_u8600_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~B*A))"),
    .INIT(16'h0d0f))
    _al_u8601 (
    .a(data_rd[32]),
    .b(ex_size[2]),
    .c(shift_l),
    .d(shift_r),
    .o(_al_u8601_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D*~A)))"),
    .INIT(16'h4c0c))
    _al_u8602 (
    .a(\exu/lsu/n56 ),
    .b(_al_u8601_o),
    .c(data_rd[31]),
    .d(shift_r),
    .o(_al_u8602_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*~C))"),
    .INIT(16'h4044))
    _al_u8603 (
    .a(_al_u8602_o),
    .b(_al_u2855_o),
    .c(data_rd[30]),
    .d(shift_l),
    .o(_al_u8603_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8604 (
    .a(_al_u8592_o),
    .b(_al_u8594_o),
    .c(_al_u8600_o),
    .d(_al_u8603_o),
    .o(\exu/n64 [31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u8605 (
    .a(uncache_data[30]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [30]),
    .o(_al_u8605_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u8606 (
    .a(_al_u8444_o),
    .b(_al_u8605_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8606_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h5300))
    _al_u8607 (
    .a(_al_u8146_o),
    .b(_al_u8286_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8607_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8608 (
    .a(_al_u8606_o),
    .b(_al_u8607_o),
    .c(_al_u7912_o),
    .o(_al_u8608_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8609 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[30]),
    .o(_al_u8609_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8610 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8608_o),
    .d(_al_u8609_o),
    .o(_al_u8610_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8611 (
    .a(uncache_data[46]),
    .b(uncache_data[38]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8611_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8612 (
    .a(uncache_data[54]),
    .b(uncache_data[30]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8612_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8613 (
    .a(_al_u8611_o),
    .b(_al_u8612_o),
    .c(_al_u7912_o),
    .o(_al_u8613_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8614 (
    .a(_al_u7991_o),
    .b(_al_u8613_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8614_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8615 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[30]),
    .d(ds2[30]),
    .o(_al_u8615_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8616 (
    .a(\exu/alu_au/sub_64 [30]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[30]),
    .o(_al_u8616_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8617 (
    .a(_al_u8615_o),
    .b(_al_u8616_o),
    .c(\exu/alu_au/add_64 [30]),
    .d(rd_data_add),
    .o(_al_u8617_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8618 (
    .a(_al_u8617_o),
    .b(rd_data_xor),
    .c(ds1[30]),
    .d(ds2[30]),
    .o(_al_u8618_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8619 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[30]),
    .d(ds2[30]),
    .o(\exu/alu_au/n33 [30]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8620 (
    .a(_al_u8618_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [30]),
    .o(_al_u8620_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8621 (
    .a(data_rd[30]),
    .b(data_rd[31]),
    .c(shift_r),
    .o(\exu/n57 [30]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8622 (
    .a(_al_u2855_o),
    .b(\exu/n57 [30]),
    .c(data_rd[29]),
    .d(shift_l),
    .o(_al_u8622_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8623 (
    .a(_al_u8610_o),
    .b(_al_u8614_o),
    .c(_al_u8620_o),
    .d(_al_u8622_o),
    .o(\exu/n64 [30]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8624 (
    .a(\biu/l1d_out [37]),
    .b(uncache_data[37]),
    .c(_al_u3224_o),
    .o(_al_u8624_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u8625 (
    .a(\biu/l1d_out [29]),
    .b(_al_u3224_o),
    .c(uncache_data[29]),
    .o(_al_u8625_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h0053))
    _al_u8626 (
    .a(_al_u8624_o),
    .b(_al_u8625_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8626_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u8627 (
    .a(_al_u8164_o),
    .b(_al_u8306_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8627_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8628 (
    .a(_al_u8626_o),
    .b(_al_u8627_o),
    .c(_al_u7912_o),
    .o(_al_u8628_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8629 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[29]),
    .o(_al_u8629_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8630 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8628_o),
    .d(_al_u8629_o),
    .o(_al_u8630_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8631 (
    .a(uncache_data[45]),
    .b(uncache_data[29]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8631_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8632 (
    .a(uncache_data[53]),
    .b(uncache_data[37]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8632_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8633 (
    .a(_al_u8631_o),
    .b(_al_u8632_o),
    .c(_al_u7912_o),
    .o(_al_u8633_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8634 (
    .a(_al_u7991_o),
    .b(_al_u8633_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8634_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8635 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[29]),
    .d(ds2[29]),
    .o(_al_u8635_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8636 (
    .a(\exu/alu_au/sub_64 [29]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[29]),
    .o(_al_u8636_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8637 (
    .a(_al_u8635_o),
    .b(_al_u8636_o),
    .c(\exu/alu_au/add_64 [29]),
    .d(rd_data_add),
    .o(_al_u8637_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8638 (
    .a(_al_u8637_o),
    .b(rd_data_xor),
    .c(ds1[29]),
    .d(ds2[29]),
    .o(_al_u8638_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8639 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[29]),
    .d(ds2[29]),
    .o(\exu/alu_au/n33 [29]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8640 (
    .a(_al_u8638_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [29]),
    .o(_al_u8640_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8641 (
    .a(data_rd[29]),
    .b(data_rd[30]),
    .c(shift_r),
    .o(\exu/n57 [29]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8642 (
    .a(_al_u2855_o),
    .b(\exu/n57 [29]),
    .c(data_rd[28]),
    .d(shift_l),
    .o(_al_u8642_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8643 (
    .a(_al_u8630_o),
    .b(_al_u8634_o),
    .c(_al_u8640_o),
    .d(_al_u8642_o),
    .o(\exu/n64 [29]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u8644 (
    .a(\biu/l1d_out [36]),
    .b(_al_u3224_o),
    .c(_al_u8488_o),
    .o(_al_u8644_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8645 (
    .a(uncache_data[28]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [28]),
    .o(_al_u8645_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h0053))
    _al_u8646 (
    .a(_al_u8644_o),
    .b(_al_u8645_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8646_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u8647 (
    .a(_al_u8180_o),
    .b(_al_u8327_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8647_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8648 (
    .a(_al_u8646_o),
    .b(_al_u8647_o),
    .c(_al_u7912_o),
    .o(_al_u8648_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8649 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[28]),
    .o(_al_u8649_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8650 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8648_o),
    .d(_al_u8649_o),
    .o(_al_u8650_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8651 (
    .a(uncache_data[52]),
    .b(uncache_data[36]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8651_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8652 (
    .a(uncache_data[44]),
    .b(uncache_data[28]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8652_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8653 (
    .a(_al_u8651_o),
    .b(_al_u8652_o),
    .c(_al_u7912_o),
    .o(_al_u8653_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8654 (
    .a(_al_u7991_o),
    .b(_al_u8653_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8654_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8655 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[28]),
    .d(ds2[28]),
    .o(_al_u8655_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8656 (
    .a(\exu/alu_au/sub_64 [28]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[28]),
    .o(_al_u8656_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8657 (
    .a(_al_u8655_o),
    .b(_al_u8656_o),
    .c(\exu/alu_au/add_64 [28]),
    .d(rd_data_add),
    .o(_al_u8657_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8658 (
    .a(_al_u8657_o),
    .b(rd_data_xor),
    .c(ds1[28]),
    .d(ds2[28]),
    .o(_al_u8658_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8659 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[28]),
    .d(ds2[28]),
    .o(\exu/alu_au/n33 [28]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8660 (
    .a(_al_u8658_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [28]),
    .o(_al_u8660_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8661 (
    .a(data_rd[28]),
    .b(data_rd[29]),
    .c(shift_r),
    .o(\exu/n57 [28]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8662 (
    .a(_al_u2855_o),
    .b(\exu/n57 [28]),
    .c(data_rd[27]),
    .d(shift_l),
    .o(_al_u8662_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8663 (
    .a(_al_u8650_o),
    .b(_al_u8654_o),
    .c(_al_u8660_o),
    .d(_al_u8662_o),
    .o(\exu/n64 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfacf))
    _al_u8664 (
    .a(_al_u8345_o),
    .b(_al_u8508_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8664_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8665 (
    .a(uncache_data[27]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [27]),
    .o(_al_u8665_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ffc))
    _al_u8666 (
    .a(_al_u8198_o),
    .b(_al_u8665_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8666_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8667 (
    .a(_al_u8664_o),
    .b(_al_u8666_o),
    .c(_al_u7912_o),
    .o(_al_u8667_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8668 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[27]),
    .o(_al_u8668_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8669 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8667_o),
    .d(_al_u8668_o),
    .o(_al_u8669_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8670 (
    .a(uncache_data[51]),
    .b(uncache_data[27]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8670_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8671 (
    .a(uncache_data[43]),
    .b(uncache_data[35]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8671_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8672 (
    .a(_al_u8670_o),
    .b(_al_u8671_o),
    .c(_al_u7912_o),
    .o(_al_u8672_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8673 (
    .a(_al_u7991_o),
    .b(_al_u8672_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8673_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8674 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[27]),
    .d(ds2[27]),
    .o(_al_u8674_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8675 (
    .a(\exu/alu_au/sub_64 [27]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[27]),
    .o(_al_u8675_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8676 (
    .a(_al_u8674_o),
    .b(_al_u8675_o),
    .c(\exu/alu_au/add_64 [27]),
    .d(rd_data_add),
    .o(_al_u8676_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8677 (
    .a(_al_u8676_o),
    .b(rd_data_xor),
    .c(ds1[27]),
    .d(ds2[27]),
    .o(_al_u8677_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8678 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[27]),
    .d(ds2[27]),
    .o(\exu/alu_au/n33 [27]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8679 (
    .a(_al_u8677_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [27]),
    .o(_al_u8679_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8680 (
    .a(data_rd[27]),
    .b(data_rd[28]),
    .c(shift_r),
    .o(\exu/n57 [27]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8681 (
    .a(_al_u2855_o),
    .b(\exu/n57 [27]),
    .c(data_rd[26]),
    .d(shift_l),
    .o(_al_u8681_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8682 (
    .a(_al_u8669_o),
    .b(_al_u8673_o),
    .c(_al_u8679_o),
    .d(_al_u8681_o),
    .o(\exu/n64 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfa3f))
    _al_u8683 (
    .a(_al_u8364_o),
    .b(_al_u8531_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8683_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u8684 (
    .a(uncache_data[26]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [26]),
    .o(_al_u8684_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haff3))
    _al_u8685 (
    .a(_al_u8215_o),
    .b(_al_u8684_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8685_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8686 (
    .a(_al_u8683_o),
    .b(_al_u8685_o),
    .c(_al_u7912_o),
    .o(_al_u8686_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8687 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[26]),
    .o(_al_u8687_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8688 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8686_o),
    .d(_al_u8687_o),
    .o(_al_u8688_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8689 (
    .a(uncache_data[50]),
    .b(uncache_data[34]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8689_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8690 (
    .a(uncache_data[42]),
    .b(uncache_data[26]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8690_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8691 (
    .a(_al_u8689_o),
    .b(_al_u8690_o),
    .c(_al_u7912_o),
    .o(_al_u8691_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8692 (
    .a(_al_u7991_o),
    .b(_al_u8691_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8692_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8693 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[26]),
    .d(ds2[26]),
    .o(_al_u8693_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8694 (
    .a(\exu/alu_au/sub_64 [26]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[26]),
    .o(_al_u8694_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8695 (
    .a(_al_u8693_o),
    .b(_al_u8694_o),
    .c(\exu/alu_au/add_64 [26]),
    .d(rd_data_add),
    .o(_al_u8695_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8696 (
    .a(_al_u8695_o),
    .b(rd_data_xor),
    .c(ds1[26]),
    .d(ds2[26]),
    .o(_al_u8696_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8697 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[26]),
    .d(ds2[26]),
    .o(\exu/alu_au/n33 [26]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8698 (
    .a(_al_u8696_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [26]),
    .o(_al_u8698_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8699 (
    .a(data_rd[26]),
    .b(data_rd[27]),
    .c(shift_r),
    .o(\exu/n57 [26]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8700 (
    .a(_al_u2855_o),
    .b(\exu/n57 [26]),
    .c(data_rd[25]),
    .d(shift_l),
    .o(_al_u8700_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8701 (
    .a(_al_u8688_o),
    .b(_al_u8692_o),
    .c(_al_u8698_o),
    .d(_al_u8700_o),
    .o(\exu/n64 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf3af))
    _al_u8702 (
    .a(_al_u7906_o),
    .b(_al_u8383_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8702_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcffa))
    _al_u8703 (
    .a(_al_u7907_o),
    .b(_al_u8232_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8703_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8704 (
    .a(_al_u8702_o),
    .b(_al_u8703_o),
    .c(_al_u7912_o),
    .o(_al_u8704_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8705 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[25]),
    .o(_al_u8705_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8706 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8704_o),
    .d(_al_u8705_o),
    .o(_al_u8706_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8707 (
    .a(uncache_data[49]),
    .b(uncache_data[33]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8707_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8708 (
    .a(uncache_data[41]),
    .b(uncache_data[25]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8708_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8709 (
    .a(_al_u8707_o),
    .b(_al_u8708_o),
    .c(_al_u7912_o),
    .o(_al_u8709_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8710 (
    .a(_al_u7991_o),
    .b(_al_u8709_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8710_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8711 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[25]),
    .d(ds2[25]),
    .o(_al_u8711_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8712 (
    .a(\exu/alu_au/sub_64 [25]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[25]),
    .o(_al_u8712_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8713 (
    .a(_al_u8711_o),
    .b(_al_u8712_o),
    .c(\exu/alu_au/add_64 [25]),
    .d(rd_data_add),
    .o(_al_u8713_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8714 (
    .a(_al_u8713_o),
    .b(rd_data_xor),
    .c(ds1[25]),
    .d(ds2[25]),
    .o(_al_u8714_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8715 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[25]),
    .d(ds2[25]),
    .o(\exu/alu_au/n33 [25]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8716 (
    .a(_al_u8714_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [25]),
    .o(_al_u8716_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8717 (
    .a(data_rd[25]),
    .b(data_rd[26]),
    .c(shift_r),
    .o(\exu/n57 [25]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8718 (
    .a(_al_u2855_o),
    .b(\exu/n57 [25]),
    .c(data_rd[24]),
    .d(shift_l),
    .o(_al_u8718_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8719 (
    .a(_al_u8706_o),
    .b(_al_u8710_o),
    .c(_al_u8716_o),
    .d(_al_u8718_o),
    .o(\exu/n64 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D))"),
    .INIT(16'h030a))
    _al_u8720 (
    .a(_al_u7932_o),
    .b(_al_u8402_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8720_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u8721 (
    .a(_al_u7936_o),
    .b(_al_u8249_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8721_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8722 (
    .a(_al_u8720_o),
    .b(_al_u8721_o),
    .c(_al_u7912_o),
    .o(_al_u8722_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8723 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[24]),
    .o(_al_u8723_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8724 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8722_o),
    .d(_al_u8723_o),
    .o(_al_u8724_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8725 (
    .a(uncache_data[40]),
    .b(uncache_data[24]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8725_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8726 (
    .a(uncache_data[48]),
    .b(uncache_data[32]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8726_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8727 (
    .a(_al_u8725_o),
    .b(_al_u8726_o),
    .c(_al_u7912_o),
    .o(_al_u8727_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8728 (
    .a(_al_u7991_o),
    .b(_al_u8727_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8728_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8729 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[24]),
    .d(ds2[24]),
    .o(_al_u8729_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8730 (
    .a(\exu/alu_au/sub_64 [24]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[24]),
    .o(_al_u8730_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8731 (
    .a(_al_u8729_o),
    .b(_al_u8730_o),
    .c(\exu/alu_au/add_64 [24]),
    .d(rd_data_add),
    .o(_al_u8731_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8732 (
    .a(_al_u8731_o),
    .b(rd_data_xor),
    .c(ds1[24]),
    .d(ds2[24]),
    .o(_al_u8732_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8733 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[24]),
    .d(ds2[24]),
    .o(\exu/alu_au/n33 [24]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8734 (
    .a(_al_u8732_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [24]),
    .o(_al_u8734_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8735 (
    .a(data_rd[24]),
    .b(data_rd[25]),
    .c(shift_r),
    .o(\exu/n57 [24]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8736 (
    .a(_al_u2855_o),
    .b(\exu/n57 [24]),
    .c(data_rd[23]),
    .d(shift_l),
    .o(_al_u8736_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8737 (
    .a(_al_u8724_o),
    .b(_al_u8728_o),
    .c(_al_u8734_o),
    .d(_al_u8736_o),
    .o(\exu/n64 [24]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8738 (
    .a(\biu/l1d_out [31]),
    .b(uncache_data[31]),
    .c(_al_u3224_o),
    .o(_al_u8738_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8739 (
    .a(\biu/l1d_out [23]),
    .b(uncache_data[23]),
    .c(_al_u3224_o),
    .o(_al_u8739_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h0053))
    _al_u8740 (
    .a(_al_u8738_o),
    .b(_al_u8739_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8740_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u8741 (
    .a(\biu/l1d_out [39]),
    .b(uncache_data[39]),
    .c(_al_u3224_o),
    .o(_al_u8741_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    _al_u8742 (
    .a(_al_u8741_o),
    .b(_al_u8267_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8742_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8743 (
    .a(_al_u8740_o),
    .b(_al_u8742_o),
    .c(_al_u7912_o),
    .o(_al_u8743_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8744 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[23]),
    .o(_al_u8744_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8745 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8743_o),
    .d(_al_u8744_o),
    .o(_al_u8745_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8746 (
    .a(uncache_data[39]),
    .b(uncache_data[23]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8746_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8747 (
    .a(uncache_data[47]),
    .b(uncache_data[31]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8747_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8748 (
    .a(_al_u8746_o),
    .b(_al_u8747_o),
    .c(_al_u7912_o),
    .o(_al_u8748_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8749 (
    .a(_al_u7991_o),
    .b(_al_u8748_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8749_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8750 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[23]),
    .d(ds2[23]),
    .o(_al_u8750_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8751 (
    .a(\exu/alu_au/sub_64 [23]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[23]),
    .o(_al_u8751_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8752 (
    .a(_al_u8750_o),
    .b(_al_u8751_o),
    .c(\exu/alu_au/add_64 [23]),
    .d(rd_data_add),
    .o(_al_u8752_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8753 (
    .a(_al_u8752_o),
    .b(rd_data_xor),
    .c(ds1[23]),
    .d(ds2[23]),
    .o(_al_u8753_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8754 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[23]),
    .d(ds2[23]),
    .o(\exu/alu_au/n33 [23]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8755 (
    .a(_al_u8753_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [23]),
    .o(_al_u8755_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8756 (
    .a(data_rd[23]),
    .b(data_rd[24]),
    .c(shift_r),
    .o(\exu/n57 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8757 (
    .a(_al_u2855_o),
    .b(\exu/n57 [23]),
    .c(data_rd[22]),
    .d(shift_l),
    .o(_al_u8757_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8758 (
    .a(_al_u8745_o),
    .b(_al_u8749_o),
    .c(_al_u8755_o),
    .d(_al_u8757_o),
    .o(\exu/n64 [23]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8759 (
    .a(uncache_data[22]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [22]),
    .o(_al_u8759_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h00a3))
    _al_u8760 (
    .a(_al_u8605_o),
    .b(_al_u8759_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8760_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h5c00))
    _al_u8761 (
    .a(_al_u8286_o),
    .b(_al_u8444_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8761_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8762 (
    .a(_al_u8760_o),
    .b(_al_u8761_o),
    .c(_al_u7912_o),
    .o(_al_u8762_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8763 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[22]),
    .o(_al_u8763_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8764 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8762_o),
    .d(_al_u8763_o),
    .o(_al_u8764_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8765 (
    .a(uncache_data[46]),
    .b(uncache_data[22]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8765_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8766 (
    .a(uncache_data[38]),
    .b(uncache_data[30]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8766_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8767 (
    .a(_al_u8765_o),
    .b(_al_u8766_o),
    .c(_al_u7912_o),
    .o(_al_u8767_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8768 (
    .a(_al_u7991_o),
    .b(_al_u8767_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8768_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8769 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[22]),
    .d(ds2[22]),
    .o(_al_u8769_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8770 (
    .a(\exu/alu_au/sub_64 [22]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[22]),
    .o(_al_u8770_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8771 (
    .a(_al_u8769_o),
    .b(_al_u8770_o),
    .c(\exu/alu_au/add_64 [22]),
    .d(rd_data_add),
    .o(_al_u8771_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8772 (
    .a(_al_u8771_o),
    .b(rd_data_xor),
    .c(ds1[22]),
    .d(ds2[22]),
    .o(_al_u8772_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8773 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[22]),
    .d(ds2[22]),
    .o(\exu/alu_au/n33 [22]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8774 (
    .a(_al_u8772_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [22]),
    .o(_al_u8774_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8775 (
    .a(data_rd[22]),
    .b(data_rd[23]),
    .c(shift_r),
    .o(\exu/n57 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8776 (
    .a(_al_u2855_o),
    .b(\exu/n57 [22]),
    .c(data_rd[21]),
    .d(shift_l),
    .o(_al_u8776_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8777 (
    .a(_al_u8764_o),
    .b(_al_u8768_o),
    .c(_al_u8774_o),
    .d(_al_u8776_o),
    .o(\exu/n64 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfacf))
    _al_u8778 (
    .a(_al_u8624_o),
    .b(_al_u8625_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8778_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u8779 (
    .a(\biu/l1d_out [21]),
    .b(_al_u3224_o),
    .c(uncache_data[21]),
    .o(_al_u8779_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8780 (
    .a(_al_u8306_o),
    .b(_al_u8779_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8780_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8781 (
    .a(_al_u8778_o),
    .b(_al_u8780_o),
    .c(_al_u7912_o),
    .o(_al_u8781_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8782 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[21]),
    .o(_al_u8782_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8783 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8781_o),
    .d(_al_u8782_o),
    .o(_al_u8783_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8784 (
    .a(uncache_data[37]),
    .b(uncache_data[21]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8784_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8785 (
    .a(uncache_data[45]),
    .b(uncache_data[29]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8785_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8786 (
    .a(_al_u8784_o),
    .b(_al_u8785_o),
    .c(_al_u7912_o),
    .o(_al_u8786_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8787 (
    .a(_al_u7991_o),
    .b(_al_u8786_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8787_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8788 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[21]),
    .d(ds2[21]),
    .o(_al_u8788_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8789 (
    .a(\exu/alu_au/sub_64 [21]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[21]),
    .o(_al_u8789_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8790 (
    .a(_al_u8788_o),
    .b(_al_u8789_o),
    .c(\exu/alu_au/add_64 [21]),
    .d(rd_data_add),
    .o(_al_u8790_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8791 (
    .a(_al_u8790_o),
    .b(rd_data_xor),
    .c(ds1[21]),
    .d(ds2[21]),
    .o(_al_u8791_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8792 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[21]),
    .d(ds2[21]),
    .o(\exu/alu_au/n33 [21]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8793 (
    .a(_al_u8791_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [21]),
    .o(_al_u8793_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8794 (
    .a(data_rd[21]),
    .b(data_rd[22]),
    .c(shift_r),
    .o(\exu/n57 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8795 (
    .a(_al_u2855_o),
    .b(\exu/n57 [21]),
    .c(data_rd[20]),
    .d(shift_l),
    .o(_al_u8795_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8796 (
    .a(_al_u8783_o),
    .b(_al_u8787_o),
    .c(_al_u8793_o),
    .d(_al_u8795_o),
    .o(\exu/n64 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfacf))
    _al_u8797 (
    .a(_al_u8644_o),
    .b(_al_u8645_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8797_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u8798 (
    .a(uncache_data[20]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [20]),
    .o(_al_u8798_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8799 (
    .a(_al_u8327_o),
    .b(_al_u8798_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8799_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8800 (
    .a(_al_u8797_o),
    .b(_al_u8799_o),
    .c(_al_u7912_o),
    .o(_al_u8800_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8801 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[20]),
    .o(_al_u8801_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8802 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8800_o),
    .d(_al_u8801_o),
    .o(_al_u8802_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8803 (
    .a(uncache_data[44]),
    .b(uncache_data[28]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8803_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8804 (
    .a(uncache_data[36]),
    .b(uncache_data[20]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8804_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8805 (
    .a(_al_u8803_o),
    .b(_al_u8804_o),
    .c(_al_u7912_o),
    .o(_al_u8805_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8806 (
    .a(_al_u7991_o),
    .b(_al_u8805_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8806_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8807 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[20]),
    .d(ds2[20]),
    .o(_al_u8807_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8808 (
    .a(\exu/alu_au/sub_64 [20]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[20]),
    .o(_al_u8808_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8809 (
    .a(_al_u8807_o),
    .b(_al_u8808_o),
    .c(\exu/alu_au/add_64 [20]),
    .d(rd_data_add),
    .o(_al_u8809_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8810 (
    .a(_al_u8809_o),
    .b(rd_data_xor),
    .c(ds1[20]),
    .d(ds2[20]),
    .o(_al_u8810_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8811 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[20]),
    .d(ds2[20]),
    .o(\exu/alu_au/n33 [20]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8812 (
    .a(_al_u8810_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [20]),
    .o(_al_u8812_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8813 (
    .a(data_rd[20]),
    .b(data_rd[21]),
    .c(shift_r),
    .o(\exu/n57 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8814 (
    .a(_al_u2855_o),
    .b(\exu/n57 [20]),
    .c(data_rd[19]),
    .d(shift_l),
    .o(_al_u8814_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8815 (
    .a(_al_u8802_o),
    .b(_al_u8806_o),
    .c(_al_u8812_o),
    .d(_al_u8814_o),
    .o(\exu/n64 [20]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u8816 (
    .a(uncache_data[19]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [19]),
    .o(_al_u8816_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h0053))
    _al_u8817 (
    .a(_al_u8665_o),
    .b(_al_u8816_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8817_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h5300))
    _al_u8818 (
    .a(_al_u8345_o),
    .b(_al_u8508_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8818_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8819 (
    .a(_al_u8817_o),
    .b(_al_u8818_o),
    .c(_al_u7912_o),
    .o(_al_u8819_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8820 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[19]),
    .o(_al_u8820_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8821 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8819_o),
    .d(_al_u8820_o),
    .o(_al_u8821_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8822 (
    .a(uncache_data[35]),
    .b(uncache_data[27]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8822_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8823 (
    .a(uncache_data[43]),
    .b(uncache_data[19]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8823_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8824 (
    .a(_al_u8822_o),
    .b(_al_u8823_o),
    .c(_al_u7912_o),
    .o(_al_u8824_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8825 (
    .a(_al_u7991_o),
    .b(_al_u8824_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8825_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8826 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[19]),
    .d(ds2[19]),
    .o(_al_u8826_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8827 (
    .a(\exu/alu_au/sub_64 [19]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[19]),
    .o(_al_u8827_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8828 (
    .a(_al_u8826_o),
    .b(_al_u8827_o),
    .c(\exu/alu_au/add_64 [19]),
    .d(rd_data_add),
    .o(_al_u8828_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8829 (
    .a(_al_u8828_o),
    .b(rd_data_xor),
    .c(ds1[19]),
    .d(ds2[19]),
    .o(_al_u8829_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8830 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[19]),
    .d(ds2[19]),
    .o(\exu/alu_au/n33 [19]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8831 (
    .a(_al_u8829_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [19]),
    .o(_al_u8831_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8832 (
    .a(data_rd[19]),
    .b(data_rd[20]),
    .c(shift_r),
    .o(\exu/n57 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8833 (
    .a(_al_u2855_o),
    .b(\exu/n57 [19]),
    .c(data_rd[18]),
    .d(shift_l),
    .o(_al_u8833_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8834 (
    .a(_al_u8821_o),
    .b(_al_u8825_o),
    .c(_al_u8831_o),
    .d(_al_u8833_o),
    .o(\exu/n64 [19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u8835 (
    .a(\biu/l1d_out [18]),
    .b(_al_u3224_o),
    .c(uncache_data[18]),
    .o(_al_u8835_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u8836 (
    .a(_al_u8684_o),
    .b(_al_u8835_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8836_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h5c00))
    _al_u8837 (
    .a(_al_u8364_o),
    .b(_al_u8531_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8837_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8838 (
    .a(_al_u8836_o),
    .b(_al_u8837_o),
    .c(_al_u7912_o),
    .o(_al_u8838_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8839 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[18]),
    .o(_al_u8839_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8840 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8838_o),
    .d(_al_u8839_o),
    .o(_al_u8840_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8841 (
    .a(uncache_data[42]),
    .b(uncache_data[26]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8841_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8842 (
    .a(uncache_data[34]),
    .b(uncache_data[18]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8842_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8843 (
    .a(_al_u8841_o),
    .b(_al_u8842_o),
    .c(_al_u7912_o),
    .o(_al_u8843_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8844 (
    .a(_al_u7991_o),
    .b(_al_u8843_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8844_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8845 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[18]),
    .d(ds2[18]),
    .o(_al_u8845_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8846 (
    .a(\exu/alu_au/sub_64 [18]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[18]),
    .o(_al_u8846_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8847 (
    .a(_al_u8845_o),
    .b(_al_u8846_o),
    .c(\exu/alu_au/add_64 [18]),
    .d(rd_data_add),
    .o(_al_u8847_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8848 (
    .a(_al_u8847_o),
    .b(rd_data_xor),
    .c(ds1[18]),
    .d(ds2[18]),
    .o(_al_u8848_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8849 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[18]),
    .d(ds2[18]),
    .o(\exu/alu_au/n33 [18]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8850 (
    .a(_al_u8848_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [18]),
    .o(_al_u8850_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8851 (
    .a(data_rd[18]),
    .b(data_rd[19]),
    .c(shift_r),
    .o(\exu/n57 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8852 (
    .a(_al_u2855_o),
    .b(\exu/n57 [18]),
    .c(data_rd[17]),
    .d(shift_l),
    .o(_al_u8852_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8853 (
    .a(_al_u8840_o),
    .b(_al_u8844_o),
    .c(_al_u8850_o),
    .d(_al_u8852_o),
    .o(\exu/n64 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfacf))
    _al_u8854 (
    .a(_al_u7906_o),
    .b(_al_u7907_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8854_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u8855 (
    .a(_al_u7910_o),
    .b(_al_u8383_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8855_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8856 (
    .a(_al_u8854_o),
    .b(_al_u8855_o),
    .c(_al_u7912_o),
    .o(_al_u8856_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8857 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[17]),
    .o(_al_u8857_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8858 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8856_o),
    .d(_al_u8857_o),
    .o(_al_u8858_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8859 (
    .a(uncache_data[41]),
    .b(uncache_data[17]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8859_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8860 (
    .a(uncache_data[33]),
    .b(uncache_data[25]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8860_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u8861 (
    .a(_al_u8859_o),
    .b(_al_u8860_o),
    .c(_al_u7912_o),
    .o(_al_u8861_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8862 (
    .a(_al_u7991_o),
    .b(_al_u8861_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8862_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8863 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[17]),
    .d(ds2[17]),
    .o(_al_u8863_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8864 (
    .a(\exu/alu_au/sub_64 [17]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[17]),
    .o(_al_u8864_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8865 (
    .a(_al_u8863_o),
    .b(_al_u8864_o),
    .c(\exu/alu_au/add_64 [17]),
    .d(rd_data_add),
    .o(_al_u8865_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8866 (
    .a(_al_u8865_o),
    .b(rd_data_xor),
    .c(ds1[17]),
    .d(ds2[17]),
    .o(_al_u8866_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8867 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[17]),
    .d(ds2[17]),
    .o(\exu/alu_au/n33 [17]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8868 (
    .a(_al_u8866_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [17]),
    .o(_al_u8868_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8869 (
    .a(data_rd[17]),
    .b(data_rd[18]),
    .c(shift_r),
    .o(\exu/n57 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8870 (
    .a(_al_u2855_o),
    .b(\exu/n57 [17]),
    .c(data_rd[16]),
    .d(shift_l),
    .o(_al_u8870_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8871 (
    .a(_al_u8858_o),
    .b(_al_u8862_o),
    .c(_al_u8868_o),
    .d(_al_u8870_o),
    .o(\exu/n64 [17]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'h3a00))
    _al_u8872 (
    .a(_al_u7936_o),
    .b(_al_u8402_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8872_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u8873 (
    .a(_al_u7932_o),
    .b(_al_u7933_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8873_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8874 (
    .a(_al_u8872_o),
    .b(_al_u8873_o),
    .c(_al_u7912_o),
    .o(_al_u8874_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8875 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[16]),
    .o(_al_u8875_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8876 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8874_o),
    .d(_al_u8875_o),
    .o(_al_u8876_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8877 (
    .a(uncache_data[32]),
    .b(uncache_data[16]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8877_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8878 (
    .a(uncache_data[40]),
    .b(uncache_data[24]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8878_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u8879 (
    .a(_al_u8877_o),
    .b(_al_u8878_o),
    .c(_al_u7912_o),
    .o(_al_u8879_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*A)))"),
    .INIT(16'h020f))
    _al_u8880 (
    .a(_al_u7991_o),
    .b(_al_u8879_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8880_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8881 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[16]),
    .d(ds2[16]),
    .o(_al_u8881_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8882 (
    .a(\exu/alu_au/sub_64 [16]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[16]),
    .o(_al_u8882_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8883 (
    .a(_al_u8881_o),
    .b(_al_u8882_o),
    .c(\exu/alu_au/add_64 [16]),
    .d(rd_data_add),
    .o(_al_u8883_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8884 (
    .a(_al_u8883_o),
    .b(rd_data_xor),
    .c(ds1[16]),
    .d(ds2[16]),
    .o(_al_u8884_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8885 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[16]),
    .d(ds2[16]),
    .o(\exu/alu_au/n33 [16]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8886 (
    .a(_al_u8884_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [16]),
    .o(_al_u8886_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8887 (
    .a(data_rd[16]),
    .b(data_rd[17]),
    .c(shift_r),
    .o(\exu/n57 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8888 (
    .a(_al_u2855_o),
    .b(\exu/n57 [16]),
    .c(data_rd[15]),
    .d(shift_l),
    .o(_al_u8888_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8889 (
    .a(_al_u8876_o),
    .b(_al_u8880_o),
    .c(_al_u8886_o),
    .d(_al_u8888_o),
    .o(\exu/n64 [16]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u8890 (
    .a(_al_u7971_o),
    .b(_al_u7912_o),
    .o(_al_u8890_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8891 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[15]),
    .o(_al_u8891_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u8892 (
    .a(_al_u7905_o),
    .b(_al_u7973_o),
    .c(_al_u8890_o),
    .d(_al_u8891_o),
    .o(_al_u8892_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u8893 (
    .a(_al_u7991_o),
    .b(_al_u7990_o),
    .c(_al_u7912_o),
    .o(_al_u8893_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u8894 (
    .a(_al_u8893_o),
    .b(\exu/c_stb_lutinv ),
    .c(\exu/n59_lutinv ),
    .o(_al_u8894_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8895 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[15]),
    .d(ds2[15]),
    .o(_al_u8895_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8896 (
    .a(\exu/alu_au/sub_64 [15]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[15]),
    .o(_al_u8896_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8897 (
    .a(_al_u8895_o),
    .b(_al_u8896_o),
    .c(\exu/alu_au/add_64 [15]),
    .d(rd_data_add),
    .o(_al_u8897_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8898 (
    .a(_al_u8897_o),
    .b(rd_data_xor),
    .c(ds1[15]),
    .d(ds2[15]),
    .o(_al_u8898_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8899 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[15]),
    .d(ds2[15]),
    .o(\exu/alu_au/n33 [15]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8900 (
    .a(_al_u8898_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [15]),
    .o(_al_u8900_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8901 (
    .a(data_rd[15]),
    .b(data_rd[16]),
    .c(shift_r),
    .o(\exu/n57 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8902 (
    .a(_al_u2855_o),
    .b(\exu/n57 [15]),
    .c(data_rd[14]),
    .d(shift_l),
    .o(_al_u8902_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8903 (
    .a(_al_u8892_o),
    .b(_al_u8894_o),
    .c(_al_u8900_o),
    .d(_al_u8902_o),
    .o(\exu/n64 [15]));
  AL_MAP_LUT4 #(
    .EQN("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'hb080))
    _al_u8904 (
    .a(uncache_data[6]),
    .b(_al_u3224_o),
    .c(\exu/lsu/n0_lutinv ),
    .d(\biu/l1d_out [6]),
    .o(_al_u8904_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u8905 (
    .a(uncache_data[14]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [14]),
    .o(_al_u8905_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfa3f))
    _al_u8906 (
    .a(_al_u8759_o),
    .b(_al_u8905_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8906_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u8907 (
    .a(_al_u8904_o),
    .b(_al_u8906_o),
    .c(_al_u8605_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u8907_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8908 (
    .a(\exu/n60_lutinv ),
    .b(data_rd[6]),
    .o(_al_u8908_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(B*~A)))"),
    .INIT(16'h00f4))
    _al_u8909 (
    .a(_al_u8907_o),
    .b(_al_u7953_o),
    .c(_al_u8908_o),
    .d(\exu/n59_lutinv ),
    .o(_al_u8909_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u8910 (
    .a(uncache_data[6]),
    .b(uncache_data[30]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8910_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8911 (
    .a(uncache_data[22]),
    .b(uncache_data[14]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8911_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*A)))"),
    .INIT(16'h008f))
    _al_u8912 (
    .a(_al_u8910_o),
    .b(_al_u8911_o),
    .c(_al_u7956_o),
    .d(\exu/c_stb_lutinv ),
    .o(_al_u8912_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8913 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[6]),
    .d(ds2[6]),
    .o(_al_u8913_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8914 (
    .a(\exu/alu_au/sub_64 [6]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[6]),
    .o(_al_u8914_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8915 (
    .a(_al_u8913_o),
    .b(_al_u8914_o),
    .c(\exu/alu_au/add_64 [6]),
    .d(rd_data_add),
    .o(_al_u8915_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8916 (
    .a(_al_u8915_o),
    .b(rd_data_xor),
    .c(ds1[6]),
    .d(ds2[6]),
    .o(_al_u8916_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8917 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[6]),
    .d(ds2[6]),
    .o(\exu/alu_au/n33 [6]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8918 (
    .a(_al_u8916_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [6]),
    .o(_al_u8918_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8919 (
    .a(data_rd[6]),
    .b(data_rd[7]),
    .c(shift_r),
    .o(\exu/n57 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8920 (
    .a(_al_u2855_o),
    .b(\exu/n57 [6]),
    .c(data_rd[5]),
    .d(shift_l),
    .o(_al_u8920_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8921 (
    .a(_al_u8909_o),
    .b(_al_u8912_o),
    .c(_al_u8918_o),
    .d(_al_u8920_o),
    .o(\exu/n64 [6]));
  AL_MAP_LUT4 #(
    .EQN("(C*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'ha030))
    _al_u8922 (
    .a(_al_u8444_o),
    .b(_al_u8759_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8922_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8923 (
    .a(_al_u8605_o),
    .b(_al_u8905_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8923_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u8924 (
    .a(_al_u8922_o),
    .b(_al_u8923_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u8924_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8925 (
    .a(uncache_data[38]),
    .b(uncache_data[14]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8925_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8926 (
    .a(uncache_data[30]),
    .b(uncache_data[22]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8926_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*A))"),
    .INIT(16'h7707))
    _al_u8927 (
    .a(_al_u8925_o),
    .b(_al_u8926_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u8927_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u8928 (
    .a(\exu/lsu/n52 [10]),
    .b(_al_u8927_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8928_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8929 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[14]),
    .o(_al_u8929_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*A)))"),
    .INIT(16'h20f0))
    _al_u8930 (
    .a(_al_u7905_o),
    .b(_al_u8924_o),
    .c(_al_u8928_o),
    .d(_al_u8929_o),
    .o(_al_u8930_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8931 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[14]),
    .d(ds2[14]),
    .o(_al_u8931_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8932 (
    .a(\exu/alu_au/sub_64 [14]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[14]),
    .o(_al_u8932_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8933 (
    .a(_al_u8931_o),
    .b(_al_u8932_o),
    .c(\exu/alu_au/add_64 [14]),
    .d(rd_data_add),
    .o(_al_u8933_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8934 (
    .a(_al_u8933_o),
    .b(rd_data_xor),
    .c(ds1[14]),
    .d(ds2[14]),
    .o(_al_u8934_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(D*C)))"),
    .INIT(16'h3111))
    _al_u8935 (
    .a(_al_u8934_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/alu_and [14]),
    .d(rd_data_and),
    .o(_al_u8935_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8936 (
    .a(data_rd[14]),
    .b(data_rd[15]),
    .c(shift_r),
    .o(\exu/n57 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8937 (
    .a(_al_u2855_o),
    .b(\exu/n57 [14]),
    .c(data_rd[13]),
    .d(shift_l),
    .o(_al_u8937_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*~A))"),
    .INIT(8'hf4))
    _al_u8938 (
    .a(_al_u8930_o),
    .b(_al_u8935_o),
    .c(_al_u8937_o),
    .o(\exu/n64 [14]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u8939 (
    .a(_al_u3224_o),
    .b(\biu/l1d_out [5]),
    .o(_al_u8939_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u8940 (
    .a(uncache_data[5]),
    .b(_al_u3224_o),
    .c(\exu/lsu/n0_lutinv ),
    .o(_al_u8940_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u8941 (
    .a(_al_u8625_o),
    .b(_al_u8939_o),
    .c(_al_u8940_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u8941_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'h1d))
    _al_u8942 (
    .a(\biu/l1d_out [13]),
    .b(_al_u3224_o),
    .c(uncache_data[13]),
    .o(_al_u8942_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8943 (
    .a(_al_u8942_o),
    .b(\exu/lsu/n2_lutinv ),
    .o(_al_u8943_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u8944 (
    .a(_al_u8941_o),
    .b(_al_u8943_o),
    .c(_al_u8779_o),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u8944_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8945 (
    .a(\exu/n60_lutinv ),
    .b(data_rd[5]),
    .o(_al_u8945_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(B*~A)))"),
    .INIT(16'h00f4))
    _al_u8946 (
    .a(_al_u8944_o),
    .b(_al_u7953_o),
    .c(_al_u8945_o),
    .d(\exu/n59_lutinv ),
    .o(_al_u8946_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u8947 (
    .a(uncache_data[5]),
    .b(uncache_data[21]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8947_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8948 (
    .a(uncache_data[29]),
    .b(uncache_data[13]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8948_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(~B*~A)))"),
    .INIT(16'h001f))
    _al_u8949 (
    .a(_al_u8947_o),
    .b(_al_u8948_o),
    .c(_al_u7956_o),
    .d(\exu/c_stb_lutinv ),
    .o(_al_u8949_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8950 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[5]),
    .d(ds2[5]),
    .o(_al_u8950_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8951 (
    .a(\exu/alu_au/sub_64 [5]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[5]),
    .o(_al_u8951_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8952 (
    .a(_al_u8950_o),
    .b(_al_u8951_o),
    .c(\exu/alu_au/add_64 [5]),
    .d(rd_data_add),
    .o(_al_u8952_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8953 (
    .a(_al_u8952_o),
    .b(rd_data_xor),
    .c(ds1[5]),
    .d(ds2[5]),
    .o(_al_u8953_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8954 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[5]),
    .d(ds2[5]),
    .o(\exu/alu_au/n33 [5]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8955 (
    .a(_al_u8953_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [5]),
    .o(_al_u8955_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8956 (
    .a(data_rd[5]),
    .b(data_rd[6]),
    .c(shift_r),
    .o(\exu/n57 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8957 (
    .a(_al_u2855_o),
    .b(\exu/n57 [5]),
    .c(data_rd[4]),
    .d(shift_l),
    .o(_al_u8957_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8958 (
    .a(_al_u8946_o),
    .b(_al_u8949_o),
    .c(_al_u8955_o),
    .d(_al_u8957_o),
    .o(\exu/n64 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0503))
    _al_u8959 (
    .a(_al_u8625_o),
    .b(_al_u8942_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8959_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'h50c0))
    _al_u8960 (
    .a(_al_u8624_o),
    .b(_al_u8779_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8960_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u8961 (
    .a(_al_u8959_o),
    .b(_al_u8960_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u8961_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8962 (
    .a(uncache_data[29]),
    .b(uncache_data[21]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8962_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u8963 (
    .a(uncache_data[37]),
    .b(uncache_data[13]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8963_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*A))"),
    .INIT(16'h7707))
    _al_u8964 (
    .a(_al_u8962_o),
    .b(_al_u8963_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u8964_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u8965 (
    .a(\exu/lsu/n52 [10]),
    .b(_al_u8964_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u8965_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u8966 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[13]),
    .o(_al_u8966_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*A)))"),
    .INIT(16'h20f0))
    _al_u8967 (
    .a(_al_u7905_o),
    .b(_al_u8961_o),
    .c(_al_u8965_o),
    .d(_al_u8966_o),
    .o(_al_u8967_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8968 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[13]),
    .d(ds2[13]),
    .o(_al_u8968_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8969 (
    .a(\exu/alu_au/sub_64 [13]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[13]),
    .o(_al_u8969_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8970 (
    .a(_al_u8968_o),
    .b(_al_u8969_o),
    .c(\exu/alu_au/add_64 [13]),
    .d(rd_data_add),
    .o(_al_u8970_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8971 (
    .a(_al_u8970_o),
    .b(rd_data_xor),
    .c(ds1[13]),
    .d(ds2[13]),
    .o(_al_u8971_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(D*C)))"),
    .INIT(16'h3111))
    _al_u8972 (
    .a(_al_u8971_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/alu_and [13]),
    .d(rd_data_and),
    .o(_al_u8972_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8973 (
    .a(data_rd[13]),
    .b(data_rd[14]),
    .c(shift_r),
    .o(\exu/n57 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8974 (
    .a(_al_u2855_o),
    .b(\exu/n57 [13]),
    .c(data_rd[12]),
    .d(shift_l),
    .o(_al_u8974_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*~A))"),
    .INIT(8'hf4))
    _al_u8975 (
    .a(_al_u8967_o),
    .b(_al_u8972_o),
    .c(_al_u8974_o),
    .o(\exu/n64 [13]));
  AL_MAP_LUT4 #(
    .EQN("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'hb080))
    _al_u8976 (
    .a(uncache_data[4]),
    .b(_al_u3224_o),
    .c(\exu/lsu/n0_lutinv ),
    .d(\biu/l1d_out [4]),
    .o(_al_u8976_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u8977 (
    .a(uncache_data[12]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [12]),
    .o(_al_u8977_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8978 (
    .a(_al_u8798_o),
    .b(_al_u8977_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8978_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*~C))"),
    .INIT(16'h4044))
    _al_u8979 (
    .a(_al_u8976_o),
    .b(_al_u8978_o),
    .c(_al_u8645_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u8979_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u8980 (
    .a(\exu/n60_lutinv ),
    .b(data_rd[4]),
    .o(_al_u8980_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(B*~A)))"),
    .INIT(16'h00f4))
    _al_u8981 (
    .a(_al_u8979_o),
    .b(_al_u7953_o),
    .c(_al_u8980_o),
    .d(\exu/n59_lutinv ),
    .o(_al_u8981_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u8982 (
    .a(uncache_data[20]),
    .b(uncache_data[12]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8982_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u8983 (
    .a(uncache_data[4]),
    .b(uncache_data[28]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8983_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*A)))"),
    .INIT(16'h008f))
    _al_u8984 (
    .a(_al_u8982_o),
    .b(_al_u8983_o),
    .c(_al_u7956_o),
    .d(\exu/c_stb_lutinv ),
    .o(_al_u8984_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u8985 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[4]),
    .d(ds2[4]),
    .o(_al_u8985_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u8986 (
    .a(\exu/alu_au/sub_64 [4]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[4]),
    .o(_al_u8986_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u8987 (
    .a(_al_u8985_o),
    .b(_al_u8986_o),
    .c(\exu/alu_au/add_64 [4]),
    .d(rd_data_add),
    .o(_al_u8987_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u8988 (
    .a(_al_u8987_o),
    .b(rd_data_xor),
    .c(ds1[4]),
    .d(ds2[4]),
    .o(_al_u8988_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u8989 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[4]),
    .d(ds2[4]),
    .o(\exu/alu_au/n33 [4]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u8990 (
    .a(_al_u8988_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [4]),
    .o(_al_u8990_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u8991 (
    .a(data_rd[4]),
    .b(data_rd[5]),
    .c(shift_r),
    .o(\exu/n57 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u8992 (
    .a(_al_u2855_o),
    .b(\exu/n57 [4]),
    .c(data_rd[3]),
    .d(shift_l),
    .o(_al_u8992_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u8993 (
    .a(_al_u8981_o),
    .b(_al_u8984_o),
    .c(_al_u8990_o),
    .d(_al_u8992_o),
    .o(\exu/n64 [4]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'h50c0))
    _al_u8994 (
    .a(_al_u8644_o),
    .b(_al_u8798_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8994_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'h050c))
    _al_u8995 (
    .a(_al_u8645_o),
    .b(_al_u8977_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8995_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u8996 (
    .a(_al_u8994_o),
    .b(_al_u8995_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u8996_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u8997 (
    .a(uncache_data[36]),
    .b(uncache_data[20]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8997_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u8998 (
    .a(uncache_data[28]),
    .b(uncache_data[12]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u8998_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u8999 (
    .a(_al_u8997_o),
    .b(_al_u8998_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u8999_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u9000 (
    .a(\exu/lsu/n52 [10]),
    .b(_al_u8999_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u9000_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u9001 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[12]),
    .o(_al_u9001_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*A)))"),
    .INIT(16'h20f0))
    _al_u9002 (
    .a(_al_u7905_o),
    .b(_al_u8996_o),
    .c(_al_u9000_o),
    .d(_al_u9001_o),
    .o(_al_u9002_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u9003 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[12]),
    .d(ds2[12]),
    .o(_al_u9003_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u9004 (
    .a(\exu/alu_au/sub_64 [12]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[12]),
    .o(_al_u9004_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u9005 (
    .a(_al_u9003_o),
    .b(_al_u9004_o),
    .c(\exu/alu_au/add_64 [12]),
    .d(rd_data_add),
    .o(_al_u9005_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u9006 (
    .a(_al_u9005_o),
    .b(rd_data_xor),
    .c(ds1[12]),
    .d(ds2[12]),
    .o(_al_u9006_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(D*C)))"),
    .INIT(16'h3111))
    _al_u9007 (
    .a(_al_u9006_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/alu_and [12]),
    .d(rd_data_and),
    .o(_al_u9007_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u9008 (
    .a(data_rd[12]),
    .b(data_rd[13]),
    .c(shift_r),
    .o(\exu/n57 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u9009 (
    .a(_al_u2855_o),
    .b(\exu/n57 [12]),
    .c(data_rd[11]),
    .d(shift_l),
    .o(_al_u9009_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*~A))"),
    .INIT(8'hf4))
    _al_u9010 (
    .a(_al_u9002_o),
    .b(_al_u9007_o),
    .c(_al_u9009_o),
    .o(\exu/n64 [12]));
  AL_MAP_LUT4 #(
    .EQN("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'hb080))
    _al_u9011 (
    .a(uncache_data[3]),
    .b(_al_u3224_o),
    .c(\exu/lsu/n0_lutinv ),
    .d(\biu/l1d_out [3]),
    .o(_al_u9011_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u9012 (
    .a(uncache_data[11]),
    .b(_al_u3224_o),
    .c(\biu/l1d_out [11]),
    .o(_al_u9012_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfacf))
    _al_u9013 (
    .a(_al_u8816_o),
    .b(_al_u9012_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9013_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*~C))"),
    .INIT(16'h4044))
    _al_u9014 (
    .a(_al_u9011_o),
    .b(_al_u9013_o),
    .c(_al_u8665_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u9014_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9015 (
    .a(\exu/n60_lutinv ),
    .b(data_rd[3]),
    .o(_al_u9015_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(B*~A)))"),
    .INIT(16'h00f4))
    _al_u9016 (
    .a(_al_u9014_o),
    .b(_al_u7953_o),
    .c(_al_u9015_o),
    .d(\exu/n59_lutinv ),
    .o(_al_u9016_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u9017 (
    .a(uncache_data[19]),
    .b(uncache_data[11]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9017_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ff5))
    _al_u9018 (
    .a(uncache_data[3]),
    .b(uncache_data[27]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9018_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*A)))"),
    .INIT(16'h008f))
    _al_u9019 (
    .a(_al_u9017_o),
    .b(_al_u9018_o),
    .c(_al_u7956_o),
    .d(\exu/c_stb_lutinv ),
    .o(_al_u9019_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u9020 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[3]),
    .d(ds2[3]),
    .o(_al_u9020_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u9021 (
    .a(\exu/alu_au/sub_64 [3]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[3]),
    .o(_al_u9021_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u9022 (
    .a(_al_u9020_o),
    .b(_al_u9021_o),
    .c(\exu/alu_au/add_64 [3]),
    .d(rd_data_add),
    .o(_al_u9022_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u9023 (
    .a(_al_u9022_o),
    .b(rd_data_xor),
    .c(ds1[3]),
    .d(ds2[3]),
    .o(_al_u9023_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u9024 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[3]),
    .d(ds2[3]),
    .o(\exu/alu_au/n33 [3]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9025 (
    .a(_al_u9023_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [3]),
    .o(_al_u9025_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u9026 (
    .a(data_rd[3]),
    .b(data_rd[4]),
    .c(shift_r),
    .o(\exu/n57 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u9027 (
    .a(_al_u2855_o),
    .b(\exu/n57 [3]),
    .c(data_rd[2]),
    .d(shift_l),
    .o(_al_u9027_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u9028 (
    .a(_al_u9016_o),
    .b(_al_u9019_o),
    .c(_al_u9025_o),
    .d(_al_u9027_o),
    .o(\exu/n64 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0503))
    _al_u9029 (
    .a(_al_u8665_o),
    .b(_al_u9012_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9029_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u9030 (
    .a(_al_u8508_o),
    .b(_al_u8816_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9030_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u9031 (
    .a(_al_u9029_o),
    .b(_al_u9030_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u9031_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u9032 (
    .a(uncache_data[27]),
    .b(uncache_data[11]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9032_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u9033 (
    .a(uncache_data[35]),
    .b(uncache_data[19]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9033_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u9034 (
    .a(_al_u9032_o),
    .b(_al_u9033_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u9034_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u9035 (
    .a(\exu/lsu/n52 [10]),
    .b(_al_u9034_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u9035_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u9036 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[11]),
    .o(_al_u9036_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*A)))"),
    .INIT(16'h20f0))
    _al_u9037 (
    .a(_al_u7905_o),
    .b(_al_u9031_o),
    .c(_al_u9035_o),
    .d(_al_u9036_o),
    .o(_al_u9037_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u9038 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[11]),
    .d(ds2[11]),
    .o(_al_u9038_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u9039 (
    .a(\exu/alu_au/sub_64 [11]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[11]),
    .o(_al_u9039_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u9040 (
    .a(_al_u9038_o),
    .b(_al_u9039_o),
    .c(\exu/alu_au/add_64 [11]),
    .d(rd_data_add),
    .o(_al_u9040_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u9041 (
    .a(_al_u9040_o),
    .b(rd_data_xor),
    .c(ds1[11]),
    .d(ds2[11]),
    .o(_al_u9041_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(D*C)))"),
    .INIT(16'h3111))
    _al_u9042 (
    .a(_al_u9041_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/alu_and [11]),
    .d(rd_data_and),
    .o(_al_u9042_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u9043 (
    .a(data_rd[11]),
    .b(data_rd[12]),
    .c(shift_r),
    .o(\exu/n57 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u9044 (
    .a(_al_u2855_o),
    .b(\exu/n57 [11]),
    .c(data_rd[10]),
    .d(shift_l),
    .o(_al_u9044_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*~A))"),
    .INIT(8'hf4))
    _al_u9045 (
    .a(_al_u9037_o),
    .b(_al_u9042_o),
    .c(_al_u9044_o),
    .o(\exu/n64 [11]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9046 (
    .a(_al_u3224_o),
    .b(\biu/l1d_out [2]),
    .o(_al_u9046_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u9047 (
    .a(uncache_data[2]),
    .b(_al_u3224_o),
    .c(\exu/lsu/n0_lutinv ),
    .o(_al_u9047_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u9048 (
    .a(_al_u8684_o),
    .b(_al_u9046_o),
    .c(_al_u9047_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u9048_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u9049 (
    .a(\biu/l1d_out [10]),
    .b(_al_u3224_o),
    .c(uncache_data[10]),
    .o(_al_u9049_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9050 (
    .a(_al_u9049_o),
    .b(\exu/lsu/n2_lutinv ),
    .o(_al_u9050_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u9051 (
    .a(_al_u9048_o),
    .b(_al_u9050_o),
    .c(_al_u8835_o),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u9051_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9052 (
    .a(\exu/n60_lutinv ),
    .b(data_rd[2]),
    .o(_al_u9052_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(B*~A)))"),
    .INIT(16'h00f4))
    _al_u9053 (
    .a(_al_u9051_o),
    .b(_al_u7953_o),
    .c(_al_u9052_o),
    .d(\exu/n59_lutinv ),
    .o(_al_u9053_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u9054 (
    .a(uncache_data[26]),
    .b(uncache_data[2]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9054_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf53f))
    _al_u9055 (
    .a(uncache_data[18]),
    .b(uncache_data[10]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9055_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*A)))"),
    .INIT(16'h008f))
    _al_u9056 (
    .a(_al_u9054_o),
    .b(_al_u9055_o),
    .c(_al_u7956_o),
    .d(\exu/c_stb_lutinv ),
    .o(_al_u9056_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u9057 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[2]),
    .d(ds2[2]),
    .o(_al_u9057_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u9058 (
    .a(\exu/alu_au/sub_64 [2]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[2]),
    .o(_al_u9058_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u9059 (
    .a(_al_u9057_o),
    .b(_al_u9058_o),
    .c(\exu/alu_au/add_64 [2]),
    .d(rd_data_add),
    .o(_al_u9059_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u9060 (
    .a(_al_u9059_o),
    .b(rd_data_xor),
    .c(ds1[2]),
    .d(ds2[2]),
    .o(_al_u9060_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u9061 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[2]),
    .d(ds2[2]),
    .o(\exu/alu_au/n33 [2]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9062 (
    .a(_al_u9060_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [2]),
    .o(_al_u9062_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u9063 (
    .a(data_rd[2]),
    .b(data_rd[3]),
    .c(shift_r),
    .o(\exu/n57 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u9064 (
    .a(_al_u2855_o),
    .b(\exu/n57 [2]),
    .c(data_rd[1]),
    .d(shift_l),
    .o(_al_u9064_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u9065 (
    .a(_al_u9053_o),
    .b(_al_u9056_o),
    .c(_al_u9062_o),
    .d(_al_u9064_o),
    .o(\exu/n64 [2]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u9066 (
    .a(_al_u8531_o),
    .b(_al_u8684_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9066_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u9067 (
    .a(_al_u8835_o),
    .b(_al_u9049_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9067_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u9068 (
    .a(_al_u9066_o),
    .b(_al_u9067_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u9068_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u9069 (
    .a(uncache_data[34]),
    .b(uncache_data[18]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9069_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u9070 (
    .a(uncache_data[26]),
    .b(uncache_data[10]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9070_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(~B*~A))"),
    .INIT(16'hee0e))
    _al_u9071 (
    .a(_al_u9069_o),
    .b(_al_u9070_o),
    .c(_al_u7912_o),
    .d(ex_size[1]),
    .o(_al_u9071_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u9072 (
    .a(\exu/lsu/n52 [10]),
    .b(_al_u9071_o),
    .c(\exu/c_stb_lutinv ),
    .d(\exu/n59_lutinv ),
    .o(_al_u9072_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u9073 (
    .a(\exu/n59_lutinv ),
    .b(\exu/n60_lutinv ),
    .c(data_rd[10]),
    .o(_al_u9073_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*A)))"),
    .INIT(16'h20f0))
    _al_u9074 (
    .a(_al_u7905_o),
    .b(_al_u9068_o),
    .c(_al_u9072_o),
    .d(_al_u9073_o),
    .o(_al_u9074_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u9075 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[10]),
    .d(ds2[10]),
    .o(_al_u9075_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u9076 (
    .a(\exu/alu_au/sub_64 [10]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[10]),
    .o(_al_u9076_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u9077 (
    .a(_al_u9075_o),
    .b(_al_u9076_o),
    .c(\exu/alu_au/add_64 [10]),
    .d(rd_data_add),
    .o(_al_u9077_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u9078 (
    .a(_al_u9077_o),
    .b(rd_data_xor),
    .c(ds1[10]),
    .d(ds2[10]),
    .o(_al_u9078_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(A*~(D*C)))"),
    .INIT(16'h3111))
    _al_u9079 (
    .a(_al_u9078_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/alu_and [10]),
    .d(rd_data_and),
    .o(_al_u9079_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u9080 (
    .a(data_rd[10]),
    .b(data_rd[11]),
    .c(shift_r),
    .o(\exu/n57 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u9081 (
    .a(_al_u2855_o),
    .b(\exu/n57 [10]),
    .c(data_rd[9]),
    .d(shift_l),
    .o(_al_u9081_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*~A))"),
    .INIT(8'hf4))
    _al_u9082 (
    .a(_al_u9074_o),
    .b(_al_u9079_o),
    .c(_al_u9081_o),
    .o(\exu/n64 [10]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9083 (
    .a(_al_u3224_o),
    .b(\biu/l1d_out [1]),
    .o(_al_u9083_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    _al_u9084 (
    .a(uncache_data[1]),
    .b(_al_u3224_o),
    .c(\exu/lsu/n0_lutinv ),
    .o(_al_u9084_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u9085 (
    .a(_al_u7907_o),
    .b(_al_u9083_o),
    .c(_al_u9084_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u9085_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9086 (
    .a(_al_u7909_o),
    .b(\exu/lsu/n2_lutinv ),
    .o(_al_u9086_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u9087 (
    .a(_al_u9085_o),
    .b(_al_u9086_o),
    .c(_al_u7910_o),
    .d(\exu/lsu/n5_lutinv ),
    .o(_al_u9087_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9088 (
    .a(\exu/n60_lutinv ),
    .b(data_rd[1]),
    .o(_al_u9088_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(B*~A)))"),
    .INIT(16'h00f4))
    _al_u9089 (
    .a(_al_u9087_o),
    .b(_al_u7953_o),
    .c(_al_u9088_o),
    .d(\exu/n59_lutinv ),
    .o(_al_u9089_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5ff3))
    _al_u9090 (
    .a(uncache_data[25]),
    .b(uncache_data[1]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9090_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u9091 (
    .a(uncache_data[9]),
    .b(uncache_data[17]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9091_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*A)))"),
    .INIT(16'h008f))
    _al_u9092 (
    .a(_al_u9090_o),
    .b(_al_u9091_o),
    .c(_al_u7956_o),
    .d(\exu/c_stb_lutinv ),
    .o(_al_u9092_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u9093 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[1]),
    .d(ds2[1]),
    .o(_al_u9093_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u9094 (
    .a(\exu/alu_au/sub_64 [1]),
    .b(rd_data_ds1),
    .c(rd_data_sub),
    .d(ds1[1]),
    .o(_al_u9094_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u9095 (
    .a(_al_u9093_o),
    .b(_al_u9094_o),
    .c(\exu/alu_au/add_64 [1]),
    .d(rd_data_add),
    .o(_al_u9095_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u9096 (
    .a(_al_u9095_o),
    .b(rd_data_xor),
    .c(ds1[1]),
    .d(ds2[1]),
    .o(_al_u9096_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u9097 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[1]),
    .d(ds2[1]),
    .o(\exu/alu_au/n33 [1]));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9098 (
    .a(_al_u9096_o),
    .b(_al_u2855_o),
    .c(\exu/alu_au/n33 [1]),
    .o(_al_u9098_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u9099 (
    .a(data_rd[1]),
    .b(data_rd[2]),
    .c(shift_r),
    .o(\exu/n57 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'ha088))
    _al_u9100 (
    .a(_al_u2855_o),
    .b(\exu/n57 [1]),
    .c(data_rd[0]),
    .d(shift_l),
    .o(_al_u9100_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u9101 (
    .a(_al_u9089_o),
    .b(_al_u9092_o),
    .c(_al_u9098_o),
    .d(_al_u9100_o),
    .o(\exu/n64 [1]));
  AL_MAP_LUT4 #(
    .EQN("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'hb080))
    _al_u9102 (
    .a(uncache_data[0]),
    .b(_al_u3224_o),
    .c(\exu/lsu/n0_lutinv ),
    .d(\biu/l1d_out [0]),
    .o(_al_u9102_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf5cf))
    _al_u9103 (
    .a(_al_u7933_o),
    .b(_al_u7935_o),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9103_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(D*C))"),
    .INIT(16'h0444))
    _al_u9104 (
    .a(_al_u9102_o),
    .b(_al_u9103_o),
    .c(_al_u7932_o),
    .d(\exu/lsu/n8_lutinv ),
    .o(_al_u9104_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9105 (
    .a(\exu/n60_lutinv ),
    .b(data_rd[0]),
    .o(_al_u9105_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(B*~A)))"),
    .INIT(16'h00f4))
    _al_u9106 (
    .a(_al_u9104_o),
    .b(_al_u7953_o),
    .c(_al_u9105_o),
    .d(\exu/n59_lutinv ),
    .o(_al_u9106_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf35f))
    _al_u9107 (
    .a(uncache_data[8]),
    .b(uncache_data[16]),
    .c(addr_ex[0]),
    .d(addr_ex[1]),
    .o(_al_u9107_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u9108 (
    .a(_al_u9107_o),
    .b(uncache_data[24]),
    .c(\exu/lsu/n8_lutinv ),
    .o(_al_u9108_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9109 (
    .a(uncache_data[0]),
    .b(\exu/lsu/n0_lutinv ),
    .o(\exu/lsu/n22 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(~B*A)))"),
    .INIT(16'h002f))
    _al_u9110 (
    .a(_al_u9108_o),
    .b(\exu/lsu/n22 [0]),
    .c(_al_u7956_o),
    .d(\exu/c_stb_lutinv ),
    .o(_al_u9110_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(~D*~C)))"),
    .INIT(16'h222a))
    _al_u9111 (
    .a(\exu/c_stb_lutinv ),
    .b(rd_data_or),
    .c(ds1[0]),
    .d(ds2[0]),
    .o(_al_u9111_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u9112 (
    .a(\exu/alu_au/add_64 [0]),
    .b(rd_data_add),
    .c(rd_data_ds1),
    .d(ds1[0]),
    .o(_al_u9112_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u9113 (
    .a(_al_u9111_o),
    .b(_al_u9112_o),
    .c(\exu/alu_au/sub_64 [0]),
    .d(rd_data_sub),
    .o(_al_u9113_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u9114 (
    .a(_al_u9113_o),
    .b(rd_data_xor),
    .c(ds1[0]),
    .d(ds2[0]),
    .o(_al_u9114_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9115 (
    .a(\exu/alu_au/ds1_light_than_ds2_lutinv ),
    .b(rd_data_slt),
    .o(\exu/alu_au/n39 [0]));
  AL_MAP_LUT4 #(
    .EQN("(C*B*(D@A))"),
    .INIT(16'h4080))
    _al_u9116 (
    .a(and_clr),
    .b(rd_data_and),
    .c(ds1[0]),
    .d(ds2[0]),
    .o(\exu/alu_au/n33 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~B*A))"),
    .INIT(16'h0f0d))
    _al_u9117 (
    .a(_al_u9114_o),
    .b(\exu/alu_au/n39 [0]),
    .c(_al_u2855_o),
    .d(\exu/alu_au/n33 [0]),
    .o(_al_u9117_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u9118 (
    .a(data_rd[0]),
    .b(data_rd[1]),
    .c(shift_r),
    .o(_al_u9118_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u9119 (
    .a(_al_u2855_o),
    .b(_al_u9118_o),
    .c(shift_l),
    .o(_al_u9119_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*~(B*~A)))"),
    .INIT(16'hffb0))
    _al_u9120 (
    .a(_al_u9106_o),
    .b(_al_u9110_o),
    .c(_al_u9117_o),
    .d(_al_u9119_o),
    .o(\exu/n64 [0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9121 (
    .a(cache_flush),
    .b(cache_reset),
    .o(_al_u9121_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u9122 (
    .a(_al_u2852_o),
    .b(_al_u9121_o),
    .c(amo),
    .o(_al_u9122_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u9123 (
    .a(ex_ill_ins),
    .b(ex_ins_acc_fault),
    .c(ex_ins_addr_mis),
    .d(ex_ins_page_fault),
    .o(\exu/n17_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u9124 (
    .a(\exu/c_stb_lutinv ),
    .b(\exu/n17_lutinv ),
    .c(ex_valid),
    .o(\exu/n19 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(~D*~A))"),
    .INIT(16'h0c08))
    _al_u9125 (
    .a(_al_u9122_o),
    .b(\exu/n19 ),
    .c(load),
    .d(store),
    .o(_al_u9125_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u9126 (
    .a(_al_u6309_o),
    .b(_al_u6320_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [7]),
    .d(\biu/cache_ctrl_logic/l1d_pte [7]),
    .o(_al_u9126_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(~D*B)))"),
    .INIT(16'h0a0e))
    _al_u9127 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u3222_o),
    .c(_al_u2848_o),
    .d(_al_u7150_o),
    .o(_al_u9127_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(B*A)))"),
    .INIT(16'h80f0))
    _al_u9128 (
    .a(_al_u6426_o),
    .b(_al_u9126_o),
    .c(_al_u9127_o),
    .d(\biu/cache_ctrl_logic/n55_lutinv ),
    .o(_al_u9128_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9129 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u3224_o),
    .o(_al_u9129_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u9130 (
    .a(ex_more_exception_neg_lutinv),
    .b(_al_u9128_o),
    .c(_al_u9129_o),
    .o(_al_u9130_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(B*C*~(D)+~(B)*~(C)*D))"),
    .INIT(16'h0140))
    _al_u9131 (
    .a(_al_u9130_o),
    .b(\exu/main_state [0]),
    .c(\exu/main_state [1]),
    .d(\exu/main_state [2]),
    .o(_al_u9131_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(~C*B))"),
    .INIT(8'hae))
    _al_u9132 (
    .a(_al_u9125_o),
    .b(\exu/main_state [2]),
    .c(_al_u9131_o),
    .o(\exu/n45 [2]));
  AL_MAP_LUT4 #(
    .EQN("~((D*~A)*~(B)*~(C)+(D*~A)*B*~(C)+~((D*~A))*B*C+(D*~A)*B*C)"),
    .INIT(16'h3a3f))
    _al_u9133 (
    .a(_al_u9131_o),
    .b(ex_more_exception_neg_lutinv),
    .c(_al_u2910_o),
    .d(\exu/main_state [3]),
    .o(_al_u9133_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u9134 (
    .a(\exu/n19 ),
    .b(load),
    .c(store),
    .o(_al_u9134_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u9135 (
    .a(_al_u9121_o),
    .b(load),
    .c(store),
    .o(_al_u9135_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u9136 (
    .a(_al_u9135_o),
    .b(_al_u2852_o),
    .c(amo),
    .o(\exu/n138_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u9137 (
    .a(_al_u9134_o),
    .b(_al_u2852_o),
    .c(\exu/n138_lutinv ),
    .o(_al_u9137_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u9138 (
    .a(_al_u9133_o),
    .b(_al_u9137_o),
    .o(\exu/n45 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u9139 (
    .a(\exu/main_state [0]),
    .b(\exu/main_state [1]),
    .c(\exu/main_state [2]),
    .d(\exu/main_state [3]),
    .o(_al_u9139_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u9140 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u3224_o),
    .c(_al_u9139_o),
    .o(\exu/n10 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u9141 (
    .a(\exu/shift_count [4]),
    .b(\exu/shift_count [5]),
    .c(\exu/shift_count [6]),
    .d(\exu/shift_count [7]),
    .o(_al_u9141_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u9142 (
    .a(\exu/shift_count [0]),
    .b(\exu/shift_count [1]),
    .c(\exu/shift_count [2]),
    .d(\exu/shift_count [3]),
    .o(_al_u9142_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u9143 (
    .a(_al_u2855_o),
    .b(_al_u9141_o),
    .c(_al_u9142_o),
    .o(\exu/shift_multi_ready ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u9144 (
    .a(\exu/n138_lutinv ),
    .b(\exu/shift_multi_ready ),
    .c(_al_u2852_o),
    .o(_al_u9144_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u9145 (
    .a(\exu/main_state [0]),
    .b(\exu/main_state [1]),
    .c(\exu/main_state [2]),
    .d(\exu/main_state [3]),
    .o(\exu/c_load_1_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(~C*~A)))"),
    .INIT(16'h04cc))
    _al_u9146 (
    .a(\exu/n10 ),
    .b(_al_u9144_o),
    .c(\exu/c_load_1_lutinv ),
    .d(load),
    .o(_al_u9146_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9147 (
    .a(\exu/c_fence_lutinv ),
    .b(_al_u9121_o),
    .o(_al_u9147_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u9148 (
    .a(_al_u6254_o),
    .b(_al_u6255_o),
    .c(amo),
    .d(store),
    .o(_al_u9148_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D*~C)))"),
    .INIT(16'h8c88))
    _al_u9149 (
    .a(_al_u9128_o),
    .b(_al_u9146_o),
    .c(_al_u9147_o),
    .d(_al_u9148_o),
    .o(_al_u9149_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u9150 (
    .a(_al_u9149_o),
    .b(ex_more_exception_neg_lutinv),
    .c(\exu/n17_lutinv ),
    .d(ex_valid),
    .o(\exu/n95 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9151 (
    .a(_al_u9130_o),
    .b(_al_u6255_o),
    .o(_al_u9151_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u9152 (
    .a(ex_more_exception_neg_lutinv),
    .b(_al_u9129_o),
    .c(_al_u2910_o),
    .o(_al_u9152_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9153 (
    .a(\exu/main_state [2]),
    .b(\exu/main_state [3]),
    .o(_al_u9153_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u9154 (
    .a(_al_u9153_o),
    .b(\exu/main_state [0]),
    .c(\exu/main_state [1]),
    .o(_al_u9154_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u9155 (
    .a(_al_u9151_o),
    .b(_al_u9152_o),
    .c(_al_u9154_o),
    .o(_al_u9155_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u9156 (
    .a(\exu/n10 ),
    .b(\exu/n19 ),
    .c(load),
    .o(_al_u9156_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u9157 (
    .a(_al_u9155_o),
    .b(_al_u9156_o),
    .c(\exu/n19 ),
    .o(\exu/n45 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hbc30))
    _al_u9158 (
    .a(_al_u9130_o),
    .b(_al_u9153_o),
    .c(\exu/main_state [0]),
    .d(\exu/main_state [1]),
    .o(_al_u9158_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9159 (
    .a(_al_u9158_o),
    .b(\exu/shift_multi_ready ),
    .o(_al_u9159_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u9160 (
    .a(ex_more_exception_neg_lutinv),
    .b(_al_u2910_o),
    .c(_al_u9139_o),
    .o(_al_u9160_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9161 (
    .a(_al_u9160_o),
    .b(_al_u9128_o),
    .o(_al_u9161_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9162 (
    .a(_al_u9134_o),
    .b(_al_u2852_o),
    .o(_al_u9162_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u9163 (
    .a(_al_u9159_o),
    .b(_al_u9161_o),
    .c(_al_u9162_o),
    .o(\exu/n45 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(~D*A))"),
    .INIT(16'hc341))
    _al_u9164 (
    .a(id_rs2_index[4]),
    .b(id_rs2_index[0]),
    .c(wb_rd_index[0]),
    .d(wb_rd_index[4]),
    .o(_al_u9164_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u9165 (
    .a(id_rs2_index[2]),
    .b(wb_rd_index[2]),
    .o(_al_u9165_o));
  AL_MAP_LUT4 #(
    .EQN("(D*B*~(C*~A))"),
    .INIT(16'h8c00))
    _al_u9166 (
    .a(id_rs2_index[4]),
    .b(_al_u5144_o),
    .c(wb_rd_index[4]),
    .d(id_valid),
    .o(_al_u9166_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u9167 (
    .a(id_rs2_index[3]),
    .b(id_rs2_index[1]),
    .c(wb_rd_index[1]),
    .d(wb_rd_index[3]),
    .o(_al_u9167_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9168 (
    .a(_al_u9164_o),
    .b(_al_u9165_o),
    .c(_al_u9166_o),
    .d(_al_u9167_o),
    .o(_al_u9168_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u9169 (
    .a(_al_u4872_o),
    .b(id_rs1_index[4]),
    .c(id_rs1_index[3]),
    .d(id_valid),
    .o(\pip_ctrl/n34 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(~D*A))"),
    .INIT(16'hcf45))
    _al_u9170 (
    .a(id_rs1_index[3]),
    .b(id_rs1_index[0]),
    .c(wb_rd_index[0]),
    .d(wb_rd_index[3]),
    .o(_al_u9170_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*~A))"),
    .INIT(16'ha2f3))
    _al_u9171 (
    .a(id_rs1_index[4]),
    .b(id_rs1_index[0]),
    .c(wb_rd_index[0]),
    .d(wb_rd_index[4]),
    .o(_al_u9171_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u9172 (
    .a(id_rs1_index[1]),
    .b(wb_rd_index[1]),
    .o(\pip_ctrl/eq2/xor_i0[1]_i1[1]_o_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9173 (
    .a(id_ins[19]),
    .b(wb_rd_index[4]),
    .o(_al_u9173_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9174 (
    .a(id_ins[18]),
    .b(wb_rd_index[3]),
    .o(_al_u9174_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D@A))"),
    .INIT(16'h0201))
    _al_u9175 (
    .a(id_rs1_index[2]),
    .b(_al_u9173_o),
    .c(_al_u9174_o),
    .d(wb_rd_index[2]),
    .o(_al_u9175_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u9176 (
    .a(_al_u9170_o),
    .b(_al_u9171_o),
    .c(\pip_ctrl/eq2/xor_i0[1]_i1[1]_o_lutinv ),
    .d(_al_u9175_o),
    .o(_al_u9176_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9177 (
    .a(_al_u9168_o),
    .b(\pip_ctrl/n34 ),
    .c(_al_u9176_o),
    .o(_al_u9177_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D@A))"),
    .INIT(16'ha251))
    _al_u9178 (
    .a(id_rs2_index[3]),
    .b(id_rs2_index[2]),
    .c(ex_rd_index[2]),
    .d(ex_rd_index[3]),
    .o(_al_u9178_o));
  AL_MAP_LUT4 #(
    .EQN("(D*B*~(C*~A))"),
    .INIT(16'h8c00))
    _al_u9179 (
    .a(id_rs2_index[4]),
    .b(_al_u5144_o),
    .c(ex_rd_index[4]),
    .d(id_valid),
    .o(_al_u9179_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(~D*A))"),
    .INIT(16'hcf45))
    _al_u9180 (
    .a(id_rs2_index[4]),
    .b(id_rs2_index[2]),
    .c(ex_rd_index[2]),
    .d(ex_rd_index[4]),
    .o(_al_u9180_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u9181 (
    .a(id_rs2_index[1]),
    .b(id_rs2_index[0]),
    .c(ex_rd_index[0]),
    .d(ex_rd_index[1]),
    .o(_al_u9181_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9182 (
    .a(_al_u9178_o),
    .b(_al_u9179_o),
    .c(_al_u9180_o),
    .d(_al_u9181_o),
    .o(_al_u9182_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u9183 (
    .a(id_rs1_index[4]),
    .b(id_rs1_index[1]),
    .c(ex_rd_index[1]),
    .d(ex_rd_index[4]),
    .o(_al_u9183_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u9184 (
    .a(id_rs1_index[3]),
    .b(id_rs1_index[0]),
    .c(ex_rd_index[0]),
    .d(ex_rd_index[3]),
    .o(_al_u9184_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u9185 (
    .a(_al_u9183_o),
    .b(_al_u9184_o),
    .c(id_rs1_index[2]),
    .d(ex_rd_index[2]),
    .o(\pip_ctrl/n36_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9186 (
    .a(ex_gpr_write),
    .b(ex_valid),
    .o(_al_u9186_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(C*A)))"),
    .INIT(16'hec00))
    _al_u9187 (
    .a(\pip_ctrl/n34 ),
    .b(_al_u9182_o),
    .c(\pip_ctrl/n36_lutinv ),
    .d(_al_u9186_o),
    .o(\pip_ctrl/id_ex_war_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9188 (
    .a(wb_gpr_write),
    .b(wb_valid),
    .o(_al_u9188_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*~B))"),
    .INIT(16'h0405))
    _al_u9189 (
    .a(_al_u9149_o),
    .b(_al_u9177_o),
    .c(\pip_ctrl/id_ex_war_lutinv ),
    .d(_al_u9188_o),
    .o(_al_u9189_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u9190 (
    .a(id_system),
    .b(_al_u2695_o),
    .c(id_int_acc),
    .o(_al_u9190_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    _al_u9191 (
    .a(id_ill_ins),
    .b(\ins_dec/n302 ),
    .c(_al_u9190_o),
    .d(id_valid),
    .o(\pip_ctrl/id_exception ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u9192 (
    .a(ex_ebreak),
    .b(ex_ecall),
    .c(ex_jmp),
    .d(ex_system),
    .o(_al_u9192_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u9193 (
    .a(_al_u9192_o),
    .b(ex_int_acc),
    .c(ex_m_ret),
    .d(ex_s_ret),
    .o(_al_u9193_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u9194 (
    .a(ex_more_exception_neg_lutinv),
    .b(_al_u9193_o),
    .c(\exu/n17_lutinv ),
    .d(ex_valid),
    .o(\pip_ctrl/ex_exception ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u9195 (
    .a(\pip_ctrl/id_exception ),
    .b(\pip_ctrl/ex_exception ),
    .c(ex_nop),
    .o(_al_u9195_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9196 (
    .a(_al_u9189_o),
    .b(_al_u9195_o),
    .o(if_hold));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9197 (
    .a(\pip_ctrl/ex_exception ),
    .b(ex_nop),
    .o(_al_u9197_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*~B))"),
    .INIT(16'h080a))
    _al_u9198 (
    .a(_al_u9197_o),
    .b(_al_u9177_o),
    .c(\pip_ctrl/id_ex_war_lutinv ),
    .d(_al_u9188_o),
    .o(id_nop_neg_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9199 (
    .a(id_nop_neg_lutinv),
    .b(_al_u9149_o),
    .o(id_hold));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9200 (
    .a(id_nop_neg_lutinv),
    .b(\ins_dec/n107 ),
    .o(\ins_dec/u478_sel_is_0_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9201 (
    .a(if_hold),
    .b(\ins_fetch/hold ),
    .o(\ins_fetch/n9 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9202 (
    .a(_al_u9189_o),
    .b(_al_u9197_o),
    .o(\ins_dec/u461_sel_is_0_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9203 (
    .a(id_hold),
    .b(\ins_dec/n107 ),
    .o(\ins_dec/mux13_b0_sel_is_0_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9204 (
    .a(_al_u9189_o),
    .b(_al_u9195_o),
    .o(_al_u9204_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u9205 (
    .a(\biu/cache_ctrl_logic/l1i_va [13]),
    .b(\biu/cache_ctrl_logic/l1i_va [58]),
    .c(addr_if[13]),
    .d(addr_if[58]),
    .o(_al_u9205_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u9206 (
    .a(\biu/cache_ctrl_logic/l1i_va [13]),
    .b(\biu/cache_ctrl_logic/l1i_va [49]),
    .c(addr_if[13]),
    .d(addr_if[49]),
    .o(_al_u9206_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u9207 (
    .a(\biu/cache_ctrl_logic/l1i_va [18]),
    .b(\biu/cache_ctrl_logic/l1i_va [24]),
    .c(addr_if[18]),
    .d(addr_if[24]),
    .o(_al_u9207_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u9208 (
    .a(\biu/cache_ctrl_logic/l1i_va [24]),
    .b(\biu/cache_ctrl_logic/l1i_va [58]),
    .c(addr_if[24]),
    .d(addr_if[58]),
    .o(_al_u9208_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9209 (
    .a(_al_u9205_o),
    .b(_al_u9206_o),
    .c(_al_u9207_o),
    .d(_al_u9208_o),
    .o(_al_u9209_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u9210 (
    .a(\biu/cache_ctrl_logic/l1i_va [39]),
    .b(\biu/cache_ctrl_logic/l1i_va [49]),
    .c(addr_if[39]),
    .d(addr_if[49]),
    .o(_al_u9210_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u9211 (
    .a(_al_u9209_o),
    .b(_al_u9210_o),
    .c(\biu/cache_ctrl_logic/l1i_va [37]),
    .d(addr_if[37]),
    .o(_al_u9211_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u9212 (
    .a(\biu/cache_ctrl_logic/l1i_va [29]),
    .b(\biu/cache_ctrl_logic/l1i_va [31]),
    .c(addr_if[29]),
    .d(addr_if[31]),
    .o(_al_u9212_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u9213 (
    .a(\biu/cache_ctrl_logic/l1i_va [48]),
    .b(\biu/cache_ctrl_logic/l1i_va [62]),
    .c(addr_if[48]),
    .d(addr_if[62]),
    .o(_al_u9213_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u9214 (
    .a(_al_u9212_o),
    .b(_al_u9213_o),
    .c(\biu/cache_ctrl_logic/l1i_va [35]),
    .d(addr_if[35]),
    .o(_al_u9214_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u9215 (
    .a(\biu/cache_ctrl_logic/l1i_va [43]),
    .b(\biu/cache_ctrl_logic/l1i_va [45]),
    .c(addr_if[43]),
    .d(addr_if[45]),
    .o(_al_u9215_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u9216 (
    .a(\biu/cache_ctrl_logic/l1i_va [23]),
    .b(\biu/cache_ctrl_logic/l1i_va [39]),
    .c(addr_if[23]),
    .d(addr_if[39]),
    .o(_al_u9216_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u9217 (
    .a(\biu/cache_ctrl_logic/l1i_va [23]),
    .b(\biu/cache_ctrl_logic/l1i_va [37]),
    .c(addr_if[23]),
    .d(addr_if[37]),
    .o(_al_u9217_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9218 (
    .a(_al_u9214_o),
    .b(_al_u9215_o),
    .c(_al_u9216_o),
    .d(_al_u9217_o),
    .o(_al_u9218_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u9219 (
    .a(\biu/cache_ctrl_logic/l1i_va [17]),
    .b(\biu/cache_ctrl_logic/l1i_va [21]),
    .c(addr_if[17]),
    .d(addr_if[21]),
    .o(_al_u9219_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u9220 (
    .a(\biu/cache_ctrl_logic/l1i_va [19]),
    .b(\biu/cache_ctrl_logic/l1i_va [21]),
    .c(addr_if[19]),
    .d(addr_if[21]),
    .o(_al_u9220_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u9221 (
    .a(\biu/cache_ctrl_logic/l1i_va [32]),
    .b(\biu/cache_ctrl_logic/l1i_va [44]),
    .c(addr_if[32]),
    .d(addr_if[44]),
    .o(_al_u9221_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u9222 (
    .a(\biu/cache_ctrl_logic/l1i_va [16]),
    .b(\biu/cache_ctrl_logic/l1i_va [30]),
    .c(addr_if[16]),
    .d(addr_if[30]),
    .o(_al_u9222_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9223 (
    .a(_al_u9219_o),
    .b(_al_u9220_o),
    .c(_al_u9221_o),
    .d(_al_u9222_o),
    .o(_al_u9223_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u9224 (
    .a(\biu/cache_ctrl_logic/l1i_va [14]),
    .b(\biu/cache_ctrl_logic/l1i_va [40]),
    .c(addr_if[14]),
    .d(addr_if[40]),
    .o(_al_u9224_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u9225 (
    .a(\biu/cache_ctrl_logic/l1i_va [22]),
    .b(\biu/cache_ctrl_logic/l1i_va [48]),
    .c(addr_if[22]),
    .d(addr_if[48]),
    .o(_al_u9225_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u9226 (
    .a(\biu/cache_ctrl_logic/l1i_va [19]),
    .b(\biu/cache_ctrl_logic/l1i_va [60]),
    .c(addr_if[19]),
    .d(addr_if[60]),
    .o(_al_u9226_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u9227 (
    .a(\biu/cache_ctrl_logic/l1i_va [36]),
    .b(\biu/cache_ctrl_logic/l1i_va [60]),
    .c(addr_if[36]),
    .d(addr_if[60]),
    .o(_al_u9227_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9228 (
    .a(_al_u9224_o),
    .b(_al_u9225_o),
    .c(_al_u9226_o),
    .d(_al_u9227_o),
    .o(_al_u9228_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9229 (
    .a(_al_u9211_o),
    .b(_al_u9218_o),
    .c(_al_u9223_o),
    .d(_al_u9228_o),
    .o(_al_u9229_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u9230 (
    .a(\biu/cache_ctrl_logic/l1i_va [61]),
    .b(\biu/cache_ctrl_logic/l1i_va [63]),
    .c(addr_if[61]),
    .d(addr_if[63]),
    .o(_al_u9230_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u9231 (
    .a(_al_u9230_o),
    .b(\biu/cache_ctrl_logic/l1i_va [15]),
    .c(addr_if[15]),
    .o(_al_u9231_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u9232 (
    .a(\biu/cache_ctrl_logic/l1i_va [59]),
    .b(\biu/cache_ctrl_logic/l1i_va [61]),
    .c(addr_if[59]),
    .d(addr_if[61]),
    .o(_al_u9232_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u9233 (
    .a(_al_u9231_o),
    .b(_al_u9232_o),
    .c(\biu/cache_ctrl_logic/l1i_va [27]),
    .d(addr_if[27]),
    .o(_al_u9233_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u9234 (
    .a(\biu/cache_ctrl_logic/l1i_va [51]),
    .b(\biu/cache_ctrl_logic/l1i_va [55]),
    .c(addr_if[51]),
    .d(addr_if[55]),
    .o(_al_u9234_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u9235 (
    .a(_al_u9234_o),
    .b(\biu/cache_ctrl_logic/l1i_va [25]),
    .c(addr_if[25]),
    .o(_al_u9235_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u9236 (
    .a(\biu/cache_ctrl_logic/l1i_va [20]),
    .b(\biu/cache_ctrl_logic/l1i_va [56]),
    .c(addr_if[20]),
    .d(addr_if[56]),
    .o(_al_u9236_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u9237 (
    .a(\biu/cache_ctrl_logic/l1i_va [53]),
    .b(\biu/cache_ctrl_logic/l1i_va [57]),
    .c(addr_if[53]),
    .d(addr_if[57]),
    .o(_al_u9237_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u9238 (
    .a(_al_u9235_o),
    .b(_al_u9236_o),
    .c(_al_u9237_o),
    .o(_al_u9238_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u9239 (
    .a(\biu/cache_ctrl_logic/l1i_value ),
    .b(\biu/cache_ctrl_logic/l1i_va [63]),
    .c(addr_if[63]),
    .o(_al_u9239_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u9240 (
    .a(\biu/cache_ctrl_logic/l1i_va [41]),
    .b(\biu/cache_ctrl_logic/l1i_va [47]),
    .c(addr_if[41]),
    .d(addr_if[47]),
    .o(_al_u9240_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u9241 (
    .a(_al_u9239_o),
    .b(_al_u9240_o),
    .c(\biu/cache_ctrl_logic/l1i_va [33]),
    .d(addr_if[33]),
    .o(_al_u9241_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u9242 (
    .a(_al_u9233_o),
    .b(_al_u9238_o),
    .c(_al_u9241_o),
    .o(_al_u9242_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9243 (
    .a(\biu/cache_ctrl_logic/l1i_va [18]),
    .b(addr_if[18]),
    .o(_al_u9243_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9244 (
    .a(\biu/cache_ctrl_logic/l1i_va [42]),
    .b(addr_if[42]),
    .o(_al_u9244_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(D@C))"),
    .INIT(16'h1001))
    _al_u9245 (
    .a(_al_u9243_o),
    .b(_al_u9244_o),
    .c(\biu/cache_ctrl_logic/l1i_va [12]),
    .d(addr_if[12]),
    .o(_al_u9245_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u9246 (
    .a(\biu/cache_ctrl_logic/l1i_va [14]),
    .b(\biu/cache_ctrl_logic/l1i_va [22]),
    .c(addr_if[14]),
    .d(addr_if[22]),
    .o(_al_u9246_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u9247 (
    .a(\biu/cache_ctrl_logic/l1i_va [34]),
    .b(\biu/cache_ctrl_logic/l1i_va [38]),
    .c(addr_if[34]),
    .d(addr_if[38]),
    .o(_al_u9247_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u9248 (
    .a(\biu/cache_ctrl_logic/l1i_va [16]),
    .b(\biu/cache_ctrl_logic/l1i_va [36]),
    .c(addr_if[16]),
    .d(addr_if[36]),
    .o(_al_u9248_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u9249 (
    .a(\biu/cache_ctrl_logic/l1i_va [26]),
    .b(\biu/cache_ctrl_logic/l1i_va [28]),
    .c(addr_if[26]),
    .d(addr_if[28]),
    .o(_al_u9249_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9250 (
    .a(_al_u9246_o),
    .b(_al_u9247_o),
    .c(_al_u9248_o),
    .d(_al_u9249_o),
    .o(_al_u9250_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u9251 (
    .a(\biu/cache_ctrl_logic/l1i_va [38]),
    .b(\biu/cache_ctrl_logic/l1i_va [40]),
    .c(addr_if[38]),
    .d(addr_if[40]),
    .o(_al_u9251_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u9252 (
    .a(\biu/cache_ctrl_logic/l1i_va [46]),
    .b(\biu/cache_ctrl_logic/l1i_va [50]),
    .c(addr_if[46]),
    .d(addr_if[50]),
    .o(_al_u9252_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9253 (
    .a(_al_u9245_o),
    .b(_al_u9250_o),
    .c(_al_u9251_o),
    .d(_al_u9252_o),
    .o(_al_u9253_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u9254 (
    .a(\biu/cache_ctrl_logic/l1i_va [44]),
    .b(\biu/cache_ctrl_logic/l1i_va [54]),
    .c(addr_if[44]),
    .d(addr_if[54]),
    .o(_al_u9254_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u9255 (
    .a(\biu/cache_ctrl_logic/l1i_va [32]),
    .b(\biu/cache_ctrl_logic/l1i_va [34]),
    .c(addr_if[32]),
    .d(addr_if[34]),
    .o(_al_u9255_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u9256 (
    .a(\biu/cache_ctrl_logic/l1i_va [17]),
    .b(\biu/cache_ctrl_logic/l1i_va [59]),
    .c(addr_if[17]),
    .d(addr_if[59]),
    .o(_al_u9256_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u9257 (
    .a(\biu/cache_ctrl_logic/l1i_va [54]),
    .b(\biu/cache_ctrl_logic/l1i_va [62]),
    .c(addr_if[54]),
    .d(addr_if[62]),
    .o(_al_u9257_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9258 (
    .a(_al_u9254_o),
    .b(_al_u9255_o),
    .c(_al_u9256_o),
    .d(_al_u9257_o),
    .o(_al_u9258_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u9259 (
    .a(\biu/cache_ctrl_logic/l1i_va [42]),
    .b(\biu/cache_ctrl_logic/l1i_va [50]),
    .c(addr_if[42]),
    .d(addr_if[50]),
    .o(_al_u9259_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u9260 (
    .a(_al_u9259_o),
    .b(\biu/cache_ctrl_logic/l1i_va [52]),
    .c(addr_if[52]),
    .o(_al_u9260_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u9261 (
    .a(\biu/cache_ctrl_logic/l1i_va [30]),
    .b(\biu/cache_ctrl_logic/l1i_va [46]),
    .c(addr_if[30]),
    .d(addr_if[46]),
    .o(_al_u9261_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u9262 (
    .a(\biu/cache_ctrl_logic/l1i_va [26]),
    .b(\biu/cache_ctrl_logic/l1i_va [28]),
    .c(addr_if[26]),
    .d(addr_if[28]),
    .o(_al_u9262_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9263 (
    .a(_al_u9258_o),
    .b(_al_u9260_o),
    .c(_al_u9261_o),
    .d(_al_u9262_o),
    .o(_al_u9263_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9264 (
    .a(_al_u9229_o),
    .b(_al_u9242_o),
    .c(_al_u9253_o),
    .d(_al_u9263_o),
    .o(_al_u9264_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(D*A))"),
    .INIT(16'h040c))
    _al_u9265 (
    .a(\biu/bus_unit/mmu/n7_lutinv ),
    .b(_al_u6319_o),
    .c(\biu/bus_unit/mmu/n8_lutinv ),
    .d(\biu/cache_ctrl_logic/l1i_pte [4]),
    .o(_al_u9265_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u9266 (
    .a(_al_u2838_o),
    .b(\biu/cache_ctrl_logic/statu [0]),
    .c(\biu/cache_ctrl_logic/statu [1]),
    .o(_al_u9266_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(C*B*A))"),
    .INIT(16'hff80))
    _al_u9267 (
    .a(_al_u9204_o),
    .b(_al_u9264_o),
    .c(_al_u9265_o),
    .d(_al_u9266_o),
    .o(ins_page_fault));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u9268 (
    .a(_al_u6704_o),
    .b(_al_u9265_o),
    .c(\biu/cache_ctrl_logic/n55_lutinv ),
    .o(_al_u9268_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u9269 (
    .a(_al_u9189_o),
    .b(_al_u9195_o),
    .c(_al_u9268_o),
    .d(_al_u9264_o),
    .o(\ins_fetch/n27 ));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u9270 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u7149_o),
    .c(_al_u4399_o),
    .d(\biu/cache_ctrl_logic/l1i_pte [7]),
    .o(_al_u9270_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9271 (
    .a(_al_u9270_o),
    .b(_al_u3224_o),
    .o(_al_u9271_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u9272 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .c(\biu/cache_ctrl_logic/l1d_pte [7]),
    .o(_al_u9272_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~C*~(D*B)))"),
    .INIT(16'ha8a0))
    _al_u9273 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u7149_o),
    .c(_al_u3945_o),
    .d(_al_u7150_o),
    .o(_al_u9273_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u9274 (
    .a(_al_u3945_o),
    .b(_al_u7150_o),
    .c(_al_u7151_o),
    .o(_al_u9274_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9275 (
    .a(_al_u9273_o),
    .b(_al_u9274_o),
    .c(\biu/cache_ctrl_logic/statu [3]),
    .o(_al_u9275_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*~B)))"),
    .INIT(16'haa20))
    _al_u9276 (
    .a(_al_u9271_o),
    .b(_al_u9272_o),
    .c(_al_u9275_o),
    .d(_al_u4399_o),
    .o(_al_u9276_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u9277 (
    .a(_al_u7163_o),
    .b(_al_u3224_o),
    .c(_al_u4834_o),
    .o(_al_u9277_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*~A))"),
    .INIT(16'h80c0))
    _al_u9278 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u7149_o),
    .c(_al_u4834_o),
    .d(\biu/cache_ctrl_logic/pte_temp [7]),
    .o(_al_u9278_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u9279 (
    .a(_al_u9276_o),
    .b(_al_u9277_o),
    .c(_al_u9278_o),
    .o(_al_u9279_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u9280 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u7158_o),
    .c(\biu/cacheable ),
    .d(_al_u6257_o),
    .o(_al_u9280_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~B*~A))"),
    .INIT(16'h0e0f))
    _al_u9281 (
    .a(_al_u9279_o),
    .b(\biu/cache_ctrl_logic/n149 ),
    .c(_al_u9280_o),
    .d(_al_u7159_o),
    .o(_al_u9281_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9282 (
    .a(_al_u9281_o),
    .b(_al_u7193_o),
    .c(_al_u7162_o),
    .o(\biu/cache_ctrl_logic/n128 [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u9283 (
    .a(_al_u6309_o),
    .b(_al_u6257_o),
    .c(\biu/cache_ctrl_logic/n55_lutinv ),
    .o(_al_u9283_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*A))"),
    .INIT(16'h3133))
    _al_u9284 (
    .a(_al_u9204_o),
    .b(_al_u9283_o),
    .c(_al_u9264_o),
    .d(\biu/cache_ctrl_logic/n55_lutinv ),
    .o(_al_u9284_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9285 (
    .a(_al_u7193_o),
    .b(\biu/cache_ctrl_logic/l1d_pte [7]),
    .o(_al_u9285_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9286 (
    .a(_al_u7162_o),
    .b(\biu/cache_ctrl_logic/l1i_pte [7]),
    .o(_al_u9286_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9287 (
    .a(_al_u9285_o),
    .b(_al_u9286_o),
    .o(_al_u9287_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u9288 (
    .a(\biu/cache_ctrl_logic/n128 [3]),
    .b(_al_u9284_o),
    .c(_al_u9287_o),
    .o(\biu/cache_ctrl_logic/n132 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9289 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [9]),
    .d(addr_if[11]),
    .o(_al_u9289_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u9290 (
    .a(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .b(\cu_ru/trap_target_m ),
    .c(\cu_ru/stvec [0]),
    .d(\cu_ru/mtvec [0]),
    .o(_al_u9290_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9291 (
    .a(_al_u9290_o),
    .b(_al_u4138_o),
    .o(\cu_ru/mux34_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9292 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [13]),
    .c(\cu_ru/n43 [9]),
    .o(_al_u9292_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9293 (
    .a(_al_u9292_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[11]),
    .o(_al_u9293_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9294 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [11]),
    .d(\cu_ru/mepc [11]),
    .o(_al_u9294_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9295 (
    .a(_al_u9289_o),
    .b(_al_u9293_o),
    .c(pip_flush),
    .d(_al_u9294_o),
    .o(\ins_fetch/n4 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9296 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [8]),
    .d(addr_if[10]),
    .o(_al_u9296_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9297 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [12]),
    .c(\cu_ru/n43 [8]),
    .o(_al_u9297_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9298 (
    .a(_al_u9297_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[10]),
    .o(_al_u9298_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9299 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [10]),
    .d(\cu_ru/mepc [10]),
    .o(_al_u9299_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9300 (
    .a(_al_u9296_o),
    .b(_al_u9298_o),
    .c(pip_flush),
    .d(_al_u9299_o),
    .o(\ins_fetch/n4 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9301 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [7]),
    .d(addr_if[9]),
    .o(_al_u9301_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9302 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [11]),
    .c(\cu_ru/n43 [7]),
    .o(_al_u9302_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9303 (
    .a(_al_u9302_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[9]),
    .o(_al_u9303_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9304 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [9]),
    .d(\cu_ru/mepc [9]),
    .o(_al_u9304_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9305 (
    .a(_al_u9301_o),
    .b(_al_u9303_o),
    .c(pip_flush),
    .d(_al_u9304_o),
    .o(\ins_fetch/n4 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9306 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [6]),
    .d(addr_if[8]),
    .o(_al_u9306_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9307 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [10]),
    .c(\cu_ru/n43 [6]),
    .o(_al_u9307_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9308 (
    .a(_al_u9307_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[8]),
    .o(_al_u9308_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9309 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [8]),
    .d(\cu_ru/mepc [8]),
    .o(_al_u9309_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9310 (
    .a(_al_u9306_o),
    .b(_al_u9308_o),
    .c(pip_flush),
    .d(_al_u9309_o),
    .o(\ins_fetch/n4 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9311 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [61]),
    .d(addr_if[63]),
    .o(_al_u9311_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .INIT(16'h1d3f))
    _al_u9312 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [63]),
    .d(new_pc[63]),
    .o(_al_u9312_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C))"),
    .INIT(16'h08a8))
    _al_u9313 (
    .a(pip_flush),
    .b(_al_u9312_o),
    .c(\cu_ru/m_s_status/n2 ),
    .d(\cu_ru/mepc [63]),
    .o(_al_u9313_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9314 (
    .a(_al_u9311_o),
    .b(_al_u9313_o),
    .o(\ins_fetch/n4 [63]));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u9315 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(_al_u6055_o),
    .c(\cu_ru/add0_2_co ),
    .d(new_pc[62]),
    .o(_al_u9315_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C))"),
    .INIT(16'h0232))
    _al_u9316 (
    .a(_al_u9315_o),
    .b(\cu_ru/m_s_status/n2 ),
    .c(_al_u2844_o),
    .d(\cu_ru/sepc [62]),
    .o(_al_u9316_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h3120))
    _al_u9317 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [60]),
    .d(addr_if[62]),
    .o(_al_u9317_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u9318 (
    .a(pip_flush),
    .b(\cu_ru/m_s_status/n2 ),
    .c(\cu_ru/mepc [62]),
    .o(_al_u9318_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*~A))"),
    .INIT(8'hdc))
    _al_u9319 (
    .a(_al_u9316_o),
    .b(_al_u9317_o),
    .c(_al_u9318_o),
    .o(\ins_fetch/n4 [62]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9320 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [5]),
    .d(addr_if[7]),
    .o(_al_u9320_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9321 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [9]),
    .c(\cu_ru/n43 [5]),
    .o(_al_u9321_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9322 (
    .a(_al_u9321_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[7]),
    .o(_al_u9322_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9323 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [7]),
    .d(\cu_ru/mepc [7]),
    .o(_al_u9323_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9324 (
    .a(_al_u9320_o),
    .b(_al_u9322_o),
    .c(pip_flush),
    .d(_al_u9323_o),
    .o(\ins_fetch/n4 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9325 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [59]),
    .d(addr_if[61]),
    .o(_al_u9325_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9326 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [63]),
    .c(\cu_ru/n43 [59]),
    .o(_al_u9326_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9327 (
    .a(_al_u9326_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[61]),
    .o(_al_u9327_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9328 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [61]),
    .d(\cu_ru/mepc [61]),
    .o(_al_u9328_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9329 (
    .a(_al_u9325_o),
    .b(_al_u9327_o),
    .c(pip_flush),
    .d(_al_u9328_o),
    .o(\ins_fetch/n4 [61]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9330 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [58]),
    .d(addr_if[60]),
    .o(_al_u9330_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9331 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [62]),
    .c(\cu_ru/n43 [58]),
    .o(_al_u9331_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9332 (
    .a(_al_u9331_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[60]),
    .o(_al_u9332_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9333 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [60]),
    .d(\cu_ru/mepc [60]),
    .o(_al_u9333_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9334 (
    .a(_al_u9330_o),
    .b(_al_u9332_o),
    .c(pip_flush),
    .d(_al_u9333_o),
    .o(\ins_fetch/n4 [60]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9335 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [57]),
    .d(addr_if[59]),
    .o(_al_u9335_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9336 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [61]),
    .c(\cu_ru/n43 [57]),
    .o(_al_u9336_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9337 (
    .a(_al_u9336_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[59]),
    .o(_al_u9337_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9338 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [59]),
    .d(\cu_ru/mepc [59]),
    .o(_al_u9338_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9339 (
    .a(_al_u9335_o),
    .b(_al_u9337_o),
    .c(pip_flush),
    .d(_al_u9338_o),
    .o(\ins_fetch/n4 [59]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9340 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [56]),
    .d(addr_if[58]),
    .o(_al_u9340_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9341 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [60]),
    .c(\cu_ru/n43 [56]),
    .o(_al_u9341_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9342 (
    .a(_al_u9341_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[58]),
    .o(_al_u9342_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9343 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [58]),
    .d(\cu_ru/mepc [58]),
    .o(_al_u9343_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9344 (
    .a(_al_u9340_o),
    .b(_al_u9342_o),
    .c(pip_flush),
    .d(_al_u9343_o),
    .o(\ins_fetch/n4 [58]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9345 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [55]),
    .d(addr_if[57]),
    .o(_al_u9345_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9346 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [59]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [55]),
    .o(_al_u9346_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9347 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[57]),
    .o(_al_u9347_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9348 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [57]),
    .o(_al_u9348_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9349 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [57]),
    .o(_al_u9349_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9350 (
    .a(_al_u9346_o),
    .b(_al_u9347_o),
    .c(_al_u9348_o),
    .d(_al_u9349_o),
    .o(_al_u9350_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9351 (
    .a(_al_u9345_o),
    .b(_al_u9350_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [57]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9352 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [54]),
    .d(addr_if[56]),
    .o(_al_u9352_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9353 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [58]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [54]),
    .o(_al_u9353_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9354 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[56]),
    .o(_al_u9354_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9355 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [56]),
    .o(_al_u9355_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9356 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [56]),
    .o(_al_u9356_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9357 (
    .a(_al_u9353_o),
    .b(_al_u9354_o),
    .c(_al_u9355_o),
    .d(_al_u9356_o),
    .o(_al_u9357_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9358 (
    .a(_al_u9352_o),
    .b(_al_u9357_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [56]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9359 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [53]),
    .d(addr_if[55]),
    .o(_al_u9359_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9360 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [57]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [53]),
    .o(_al_u9360_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9361 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[55]),
    .o(_al_u9361_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9362 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [55]),
    .o(_al_u9362_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9363 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [55]),
    .o(_al_u9363_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9364 (
    .a(_al_u9360_o),
    .b(_al_u9361_o),
    .c(_al_u9362_o),
    .d(_al_u9363_o),
    .o(_al_u9364_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9365 (
    .a(_al_u9359_o),
    .b(_al_u9364_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [55]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9366 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [52]),
    .d(addr_if[54]),
    .o(_al_u9366_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9367 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [56]),
    .c(\cu_ru/n43 [52]),
    .o(_al_u9367_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9368 (
    .a(_al_u9367_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[54]),
    .o(_al_u9368_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9369 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [54]),
    .d(\cu_ru/mepc [54]),
    .o(_al_u9369_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9370 (
    .a(_al_u9366_o),
    .b(_al_u9368_o),
    .c(pip_flush),
    .d(_al_u9369_o),
    .o(\ins_fetch/n4 [54]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9371 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [51]),
    .d(addr_if[53]),
    .o(_al_u9371_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9372 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [55]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [51]),
    .o(_al_u9372_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9373 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[53]),
    .o(_al_u9373_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9374 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [53]),
    .o(_al_u9374_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9375 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [53]),
    .o(_al_u9375_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9376 (
    .a(_al_u9372_o),
    .b(_al_u9373_o),
    .c(_al_u9374_o),
    .d(_al_u9375_o),
    .o(_al_u9376_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9377 (
    .a(_al_u9371_o),
    .b(_al_u9376_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [53]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9378 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [50]),
    .d(addr_if[52]),
    .o(_al_u9378_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9379 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [54]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [50]),
    .o(_al_u9379_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9380 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[52]),
    .o(_al_u9380_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9381 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [52]),
    .o(_al_u9381_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9382 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [52]),
    .o(_al_u9382_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9383 (
    .a(_al_u9379_o),
    .b(_al_u9380_o),
    .c(_al_u9381_o),
    .d(_al_u9382_o),
    .o(_al_u9383_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9384 (
    .a(_al_u9378_o),
    .b(_al_u9383_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [52]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9385 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [4]),
    .d(addr_if[6]),
    .o(_al_u9385_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9386 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [8]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [4]),
    .o(_al_u9386_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9387 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[6]),
    .o(_al_u9387_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9388 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [6]),
    .o(_al_u9388_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9389 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [6]),
    .o(_al_u9389_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9390 (
    .a(_al_u9386_o),
    .b(_al_u9387_o),
    .c(_al_u9388_o),
    .d(_al_u9389_o),
    .o(_al_u9390_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9391 (
    .a(_al_u9385_o),
    .b(_al_u9390_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9392 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [49]),
    .d(addr_if[51]),
    .o(_al_u9392_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9393 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [53]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [49]),
    .o(_al_u9393_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9394 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[51]),
    .o(_al_u9394_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9395 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [51]),
    .o(_al_u9395_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9396 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [51]),
    .o(_al_u9396_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9397 (
    .a(_al_u9393_o),
    .b(_al_u9394_o),
    .c(_al_u9395_o),
    .d(_al_u9396_o),
    .o(_al_u9397_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9398 (
    .a(_al_u9392_o),
    .b(_al_u9397_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [51]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9399 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [48]),
    .d(addr_if[50]),
    .o(_al_u9399_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9400 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [52]),
    .c(\cu_ru/n43 [48]),
    .o(_al_u9400_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9401 (
    .a(_al_u9400_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[50]),
    .o(_al_u9401_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9402 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [50]),
    .d(\cu_ru/mepc [50]),
    .o(_al_u9402_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9403 (
    .a(_al_u9399_o),
    .b(_al_u9401_o),
    .c(pip_flush),
    .d(_al_u9402_o),
    .o(\ins_fetch/n4 [50]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9404 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [47]),
    .d(addr_if[49]),
    .o(_al_u9404_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9405 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [51]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [47]),
    .o(_al_u9405_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9406 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[49]),
    .o(_al_u9406_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9407 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [49]),
    .o(_al_u9407_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9408 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [49]),
    .o(_al_u9408_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9409 (
    .a(_al_u9405_o),
    .b(_al_u9406_o),
    .c(_al_u9407_o),
    .d(_al_u9408_o),
    .o(_al_u9409_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9410 (
    .a(_al_u9404_o),
    .b(_al_u9409_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [49]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9411 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [46]),
    .d(addr_if[48]),
    .o(_al_u9411_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9412 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [50]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [46]),
    .o(_al_u9412_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9413 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[48]),
    .o(_al_u9413_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9414 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [48]),
    .o(_al_u9414_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9415 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [48]),
    .o(_al_u9415_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9416 (
    .a(_al_u9412_o),
    .b(_al_u9413_o),
    .c(_al_u9414_o),
    .d(_al_u9415_o),
    .o(_al_u9416_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9417 (
    .a(_al_u9411_o),
    .b(_al_u9416_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [48]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9418 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [45]),
    .d(addr_if[47]),
    .o(_al_u9418_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9419 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [49]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [45]),
    .o(_al_u9419_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9420 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[47]),
    .o(_al_u9420_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9421 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [47]),
    .o(_al_u9421_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9422 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [47]),
    .o(_al_u9422_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9423 (
    .a(_al_u9419_o),
    .b(_al_u9420_o),
    .c(_al_u9421_o),
    .d(_al_u9422_o),
    .o(_al_u9423_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9424 (
    .a(_al_u9418_o),
    .b(_al_u9423_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [47]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9425 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [44]),
    .d(addr_if[46]),
    .o(_al_u9425_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9426 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [48]),
    .c(\cu_ru/n43 [44]),
    .o(_al_u9426_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9427 (
    .a(_al_u9426_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[46]),
    .o(_al_u9427_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9428 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [46]),
    .d(\cu_ru/mepc [46]),
    .o(_al_u9428_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9429 (
    .a(_al_u9425_o),
    .b(_al_u9427_o),
    .c(pip_flush),
    .d(_al_u9428_o),
    .o(\ins_fetch/n4 [46]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9430 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [43]),
    .d(addr_if[45]),
    .o(_al_u9430_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9431 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [47]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [43]),
    .o(_al_u9431_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9432 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[45]),
    .o(_al_u9432_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9433 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [45]),
    .o(_al_u9433_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9434 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [45]),
    .o(_al_u9434_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9435 (
    .a(_al_u9431_o),
    .b(_al_u9432_o),
    .c(_al_u9433_o),
    .d(_al_u9434_o),
    .o(_al_u9435_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9436 (
    .a(_al_u9430_o),
    .b(_al_u9435_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [45]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9437 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [42]),
    .d(addr_if[44]),
    .o(_al_u9437_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9438 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [46]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [42]),
    .o(_al_u9438_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9439 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[44]),
    .o(_al_u9439_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9440 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [44]),
    .o(_al_u9440_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9441 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [44]),
    .o(_al_u9441_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9442 (
    .a(_al_u9438_o),
    .b(_al_u9439_o),
    .c(_al_u9440_o),
    .d(_al_u9441_o),
    .o(_al_u9442_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9443 (
    .a(_al_u9437_o),
    .b(_al_u9442_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [44]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9444 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [41]),
    .d(addr_if[43]),
    .o(_al_u9444_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9445 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [45]),
    .c(\cu_ru/n43 [41]),
    .o(_al_u9445_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9446 (
    .a(_al_u9445_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[43]),
    .o(_al_u9446_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9447 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [43]),
    .d(\cu_ru/mepc [43]),
    .o(_al_u9447_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9448 (
    .a(_al_u9444_o),
    .b(_al_u9446_o),
    .c(pip_flush),
    .d(_al_u9447_o),
    .o(\ins_fetch/n4 [43]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9449 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [40]),
    .d(addr_if[42]),
    .o(_al_u9449_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9450 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [44]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [40]),
    .o(_al_u9450_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9451 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[42]),
    .o(_al_u9451_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9452 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [42]),
    .o(_al_u9452_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9453 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [42]),
    .o(_al_u9453_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9454 (
    .a(_al_u9450_o),
    .b(_al_u9451_o),
    .c(_al_u9452_o),
    .d(_al_u9453_o),
    .o(_al_u9454_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9455 (
    .a(_al_u9449_o),
    .b(_al_u9454_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [42]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9456 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [3]),
    .d(addr_if[5]),
    .o(_al_u9456_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9457 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [7]),
    .c(\cu_ru/n43 [3]),
    .o(_al_u9457_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9458 (
    .a(_al_u9457_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[5]),
    .o(_al_u9458_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9459 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [5]),
    .d(\cu_ru/mepc [5]),
    .o(_al_u9459_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9460 (
    .a(_al_u9456_o),
    .b(_al_u9458_o),
    .c(pip_flush),
    .d(_al_u9459_o),
    .o(\ins_fetch/n4 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9461 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [39]),
    .d(addr_if[41]),
    .o(_al_u9461_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9462 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [43]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [39]),
    .o(_al_u9462_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9463 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[41]),
    .o(_al_u9463_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9464 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [41]),
    .o(_al_u9464_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9465 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [41]),
    .o(_al_u9465_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9466 (
    .a(_al_u9462_o),
    .b(_al_u9463_o),
    .c(_al_u9464_o),
    .d(_al_u9465_o),
    .o(_al_u9466_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9467 (
    .a(_al_u9461_o),
    .b(_al_u9466_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [41]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9468 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [38]),
    .d(addr_if[40]),
    .o(_al_u9468_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9469 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [42]),
    .c(\cu_ru/n43 [38]),
    .o(_al_u9469_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9470 (
    .a(_al_u9469_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[40]),
    .o(_al_u9470_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9471 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [40]),
    .d(\cu_ru/mepc [40]),
    .o(_al_u9471_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9472 (
    .a(_al_u9468_o),
    .b(_al_u9470_o),
    .c(pip_flush),
    .d(_al_u9471_o),
    .o(\ins_fetch/n4 [40]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9473 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [37]),
    .d(addr_if[39]),
    .o(_al_u9473_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9474 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [41]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [37]),
    .o(_al_u9474_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9475 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[39]),
    .o(_al_u9475_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9476 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [39]),
    .o(_al_u9476_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9477 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [39]),
    .o(_al_u9477_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9478 (
    .a(_al_u9474_o),
    .b(_al_u9475_o),
    .c(_al_u9476_o),
    .d(_al_u9477_o),
    .o(_al_u9478_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9479 (
    .a(_al_u9473_o),
    .b(_al_u9478_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [39]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9480 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [36]),
    .d(addr_if[38]),
    .o(_al_u9480_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9481 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [40]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [36]),
    .o(_al_u9481_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9482 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[38]),
    .o(_al_u9482_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9483 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [38]),
    .o(_al_u9483_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9484 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [38]),
    .o(_al_u9484_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9485 (
    .a(_al_u9481_o),
    .b(_al_u9482_o),
    .c(_al_u9483_o),
    .d(_al_u9484_o),
    .o(_al_u9485_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9486 (
    .a(_al_u9480_o),
    .b(_al_u9485_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [38]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9487 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [35]),
    .d(addr_if[37]),
    .o(_al_u9487_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9488 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [39]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [35]),
    .o(_al_u9488_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9489 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[37]),
    .o(_al_u9489_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9490 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [37]),
    .o(_al_u9490_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9491 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [37]),
    .o(_al_u9491_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9492 (
    .a(_al_u9488_o),
    .b(_al_u9489_o),
    .c(_al_u9490_o),
    .d(_al_u9491_o),
    .o(_al_u9492_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9493 (
    .a(_al_u9487_o),
    .b(_al_u9492_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [37]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9494 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [34]),
    .d(addr_if[36]),
    .o(_al_u9494_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9495 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [38]),
    .c(\cu_ru/n43 [34]),
    .o(_al_u9495_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9496 (
    .a(_al_u9495_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[36]),
    .o(_al_u9496_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9497 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [36]),
    .d(\cu_ru/mepc [36]),
    .o(_al_u9497_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9498 (
    .a(_al_u9494_o),
    .b(_al_u9496_o),
    .c(pip_flush),
    .d(_al_u9497_o),
    .o(\ins_fetch/n4 [36]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9499 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [33]),
    .d(addr_if[35]),
    .o(_al_u9499_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9500 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [37]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [33]),
    .o(_al_u9500_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9501 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[35]),
    .o(_al_u9501_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9502 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [35]),
    .o(_al_u9502_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9503 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [35]),
    .o(_al_u9503_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9504 (
    .a(_al_u9500_o),
    .b(_al_u9501_o),
    .c(_al_u9502_o),
    .d(_al_u9503_o),
    .o(_al_u9504_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9505 (
    .a(_al_u9499_o),
    .b(_al_u9504_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [35]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9506 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [32]),
    .d(addr_if[34]),
    .o(_al_u9506_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9507 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [36]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [32]),
    .o(_al_u9507_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9508 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[34]),
    .o(_al_u9508_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9509 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [34]),
    .o(_al_u9509_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9510 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [34]),
    .o(_al_u9510_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9511 (
    .a(_al_u9507_o),
    .b(_al_u9508_o),
    .c(_al_u9509_o),
    .d(_al_u9510_o),
    .o(_al_u9511_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9512 (
    .a(_al_u9506_o),
    .b(_al_u9511_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [34]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9513 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [31]),
    .d(addr_if[33]),
    .o(_al_u9513_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9514 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [35]),
    .c(\cu_ru/n43 [31]),
    .o(_al_u9514_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9515 (
    .a(_al_u9514_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[33]),
    .o(_al_u9515_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9516 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [33]),
    .d(\cu_ru/mepc [33]),
    .o(_al_u9516_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9517 (
    .a(_al_u9513_o),
    .b(_al_u9515_o),
    .c(pip_flush),
    .d(_al_u9516_o),
    .o(\ins_fetch/n4 [33]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9518 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [30]),
    .d(addr_if[32]),
    .o(_al_u9518_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9519 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [34]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [30]),
    .o(_al_u9519_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9520 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[32]),
    .o(_al_u9520_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9521 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [32]),
    .o(_al_u9521_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9522 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [32]),
    .o(_al_u9522_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9523 (
    .a(_al_u9519_o),
    .b(_al_u9520_o),
    .c(_al_u9521_o),
    .d(_al_u9522_o),
    .o(_al_u9523_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9524 (
    .a(_al_u9518_o),
    .b(_al_u9523_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [32]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9525 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [2]),
    .d(addr_if[4]),
    .o(_al_u9525_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9526 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [6]),
    .c(\cu_ru/n43 [2]),
    .o(_al_u9526_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9527 (
    .a(_al_u9526_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[4]),
    .o(_al_u9527_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9528 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [4]),
    .d(\cu_ru/mepc [4]),
    .o(_al_u9528_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9529 (
    .a(_al_u9525_o),
    .b(_al_u9527_o),
    .c(pip_flush),
    .d(_al_u9528_o),
    .o(\ins_fetch/n4 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9530 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [29]),
    .d(addr_if[31]),
    .o(_al_u9530_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9531 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [33]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [29]),
    .o(_al_u9531_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9532 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[31]),
    .o(_al_u9532_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9533 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [31]),
    .o(_al_u9533_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9534 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [31]),
    .o(_al_u9534_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9535 (
    .a(_al_u9531_o),
    .b(_al_u9532_o),
    .c(_al_u9533_o),
    .d(_al_u9534_o),
    .o(_al_u9535_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9536 (
    .a(_al_u9530_o),
    .b(_al_u9535_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9537 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [28]),
    .d(addr_if[30]),
    .o(_al_u9537_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9538 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [32]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [28]),
    .o(_al_u9538_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9539 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[30]),
    .o(_al_u9539_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9540 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [30]),
    .o(_al_u9540_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9541 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [30]),
    .o(_al_u9541_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9542 (
    .a(_al_u9538_o),
    .b(_al_u9539_o),
    .c(_al_u9540_o),
    .d(_al_u9541_o),
    .o(_al_u9542_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9543 (
    .a(_al_u9537_o),
    .b(_al_u9542_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9544 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [27]),
    .d(addr_if[29]),
    .o(_al_u9544_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9545 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [31]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [27]),
    .o(_al_u9545_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9546 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[29]),
    .o(_al_u9546_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9547 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [29]),
    .o(_al_u9547_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9548 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [29]),
    .o(_al_u9548_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9549 (
    .a(_al_u9545_o),
    .b(_al_u9546_o),
    .c(_al_u9547_o),
    .d(_al_u9548_o),
    .o(_al_u9549_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9550 (
    .a(_al_u9544_o),
    .b(_al_u9549_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9551 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [26]),
    .d(addr_if[28]),
    .o(_al_u9551_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9552 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [30]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [26]),
    .o(_al_u9552_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9553 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[28]),
    .o(_al_u9553_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9554 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [28]),
    .o(_al_u9554_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9555 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [28]),
    .o(_al_u9555_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9556 (
    .a(_al_u9552_o),
    .b(_al_u9553_o),
    .c(_al_u9554_o),
    .d(_al_u9555_o),
    .o(_al_u9556_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9557 (
    .a(_al_u9551_o),
    .b(_al_u9556_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9558 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [25]),
    .d(addr_if[27]),
    .o(_al_u9558_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9559 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [29]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [25]),
    .o(_al_u9559_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9560 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[27]),
    .o(_al_u9560_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9561 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [27]),
    .o(_al_u9561_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9562 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [27]),
    .o(_al_u9562_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9563 (
    .a(_al_u9559_o),
    .b(_al_u9560_o),
    .c(_al_u9561_o),
    .d(_al_u9562_o),
    .o(_al_u9563_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9564 (
    .a(_al_u9558_o),
    .b(_al_u9563_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9565 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [24]),
    .d(addr_if[26]),
    .o(_al_u9565_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9566 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [28]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [24]),
    .o(_al_u9566_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9567 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[26]),
    .o(_al_u9567_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9568 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [26]),
    .o(_al_u9568_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9569 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [26]),
    .o(_al_u9569_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9570 (
    .a(_al_u9566_o),
    .b(_al_u9567_o),
    .c(_al_u9568_o),
    .d(_al_u9569_o),
    .o(_al_u9570_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9571 (
    .a(_al_u9565_o),
    .b(_al_u9570_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9572 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [23]),
    .d(addr_if[25]),
    .o(_al_u9572_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9573 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [27]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [23]),
    .o(_al_u9573_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9574 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[25]),
    .o(_al_u9574_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9575 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [25]),
    .o(_al_u9575_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9576 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [25]),
    .o(_al_u9576_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9577 (
    .a(_al_u9573_o),
    .b(_al_u9574_o),
    .c(_al_u9575_o),
    .d(_al_u9576_o),
    .o(_al_u9577_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9578 (
    .a(_al_u9572_o),
    .b(_al_u9577_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9579 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [22]),
    .d(addr_if[24]),
    .o(_al_u9579_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9580 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [26]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [22]),
    .o(_al_u9580_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9581 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[24]),
    .o(_al_u9581_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9582 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [24]),
    .o(_al_u9582_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9583 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [24]),
    .o(_al_u9583_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9584 (
    .a(_al_u9580_o),
    .b(_al_u9581_o),
    .c(_al_u9582_o),
    .d(_al_u9583_o),
    .o(_al_u9584_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9585 (
    .a(_al_u9579_o),
    .b(_al_u9584_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9586 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [21]),
    .d(addr_if[23]),
    .o(_al_u9586_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9587 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [25]),
    .c(\cu_ru/n43 [21]),
    .o(_al_u9587_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9588 (
    .a(_al_u9587_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[23]),
    .o(_al_u9588_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9589 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [23]),
    .d(\cu_ru/mepc [23]),
    .o(_al_u9589_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9590 (
    .a(_al_u9586_o),
    .b(_al_u9588_o),
    .c(pip_flush),
    .d(_al_u9589_o),
    .o(\ins_fetch/n4 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9591 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [20]),
    .d(addr_if[22]),
    .o(_al_u9591_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9592 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [24]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [20]),
    .o(_al_u9592_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9593 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[22]),
    .o(_al_u9593_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9594 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [22]),
    .o(_al_u9594_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9595 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [22]),
    .o(_al_u9595_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9596 (
    .a(_al_u9592_o),
    .b(_al_u9593_o),
    .c(_al_u9594_o),
    .d(_al_u9595_o),
    .o(_al_u9596_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9597 (
    .a(_al_u9591_o),
    .b(_al_u9596_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9598 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [1]),
    .d(addr_if[3]),
    .o(_al_u9598_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9599 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [5]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [1]),
    .o(_al_u9599_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9600 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[3]),
    .o(_al_u9600_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9601 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [3]),
    .o(_al_u9601_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9602 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [3]),
    .o(_al_u9602_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9603 (
    .a(_al_u9599_o),
    .b(_al_u9600_o),
    .c(_al_u9601_o),
    .d(_al_u9602_o),
    .o(_al_u9603_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9604 (
    .a(_al_u9598_o),
    .b(_al_u9603_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9605 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [19]),
    .d(addr_if[21]),
    .o(_al_u9605_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9606 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [23]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [19]),
    .o(_al_u9606_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9607 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[21]),
    .o(_al_u9607_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9608 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [21]),
    .o(_al_u9608_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9609 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [21]),
    .o(_al_u9609_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9610 (
    .a(_al_u9606_o),
    .b(_al_u9607_o),
    .c(_al_u9608_o),
    .d(_al_u9609_o),
    .o(_al_u9610_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9611 (
    .a(_al_u9605_o),
    .b(_al_u9610_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9612 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [18]),
    .d(addr_if[20]),
    .o(_al_u9612_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9613 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [22]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [18]),
    .o(_al_u9613_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9614 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[20]),
    .o(_al_u9614_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9615 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [20]),
    .o(_al_u9615_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9616 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [20]),
    .o(_al_u9616_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9617 (
    .a(_al_u9613_o),
    .b(_al_u9614_o),
    .c(_al_u9615_o),
    .d(_al_u9616_o),
    .o(_al_u9617_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9618 (
    .a(_al_u9612_o),
    .b(_al_u9617_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [20]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9619 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [17]),
    .d(addr_if[19]),
    .o(_al_u9619_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9620 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [21]),
    .c(\cu_ru/n43 [17]),
    .o(_al_u9620_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9621 (
    .a(_al_u9620_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[19]),
    .o(_al_u9621_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9622 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [19]),
    .d(\cu_ru/mepc [19]),
    .o(_al_u9622_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9623 (
    .a(_al_u9619_o),
    .b(_al_u9621_o),
    .c(pip_flush),
    .d(_al_u9622_o),
    .o(\ins_fetch/n4 [19]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9624 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [16]),
    .d(addr_if[18]),
    .o(_al_u9624_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9625 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [20]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [16]),
    .o(_al_u9625_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9626 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[18]),
    .o(_al_u9626_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9627 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [18]),
    .o(_al_u9627_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9628 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [18]),
    .o(_al_u9628_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9629 (
    .a(_al_u9625_o),
    .b(_al_u9626_o),
    .c(_al_u9627_o),
    .d(_al_u9628_o),
    .o(_al_u9629_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9630 (
    .a(_al_u9624_o),
    .b(_al_u9629_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9631 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [15]),
    .d(addr_if[17]),
    .o(_al_u9631_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9632 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [19]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [15]),
    .o(_al_u9632_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9633 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[17]),
    .o(_al_u9633_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9634 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [17]),
    .o(_al_u9634_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9635 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [17]),
    .o(_al_u9635_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9636 (
    .a(_al_u9632_o),
    .b(_al_u9633_o),
    .c(_al_u9634_o),
    .d(_al_u9635_o),
    .o(_al_u9636_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9637 (
    .a(_al_u9631_o),
    .b(_al_u9636_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9638 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [14]),
    .d(addr_if[16]),
    .o(_al_u9638_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9639 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [18]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [14]),
    .o(_al_u9639_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9640 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[16]),
    .o(_al_u9640_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9641 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [16]),
    .o(_al_u9641_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9642 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [16]),
    .o(_al_u9642_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9643 (
    .a(_al_u9639_o),
    .b(_al_u9640_o),
    .c(_al_u9641_o),
    .d(_al_u9642_o),
    .o(_al_u9643_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9644 (
    .a(_al_u9638_o),
    .b(_al_u9643_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9645 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [13]),
    .d(addr_if[15]),
    .o(_al_u9645_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9646 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [17]),
    .c(\cu_ru/n43 [13]),
    .o(_al_u9646_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9647 (
    .a(_al_u9646_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[15]),
    .o(_al_u9647_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9648 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [15]),
    .d(\cu_ru/mepc [15]),
    .o(_al_u9648_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9649 (
    .a(_al_u9645_o),
    .b(_al_u9647_o),
    .c(pip_flush),
    .d(_al_u9648_o),
    .o(\ins_fetch/n4 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9650 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [12]),
    .d(addr_if[14]),
    .o(_al_u9650_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9651 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [16]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [12]),
    .o(_al_u9651_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9652 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[14]),
    .o(_al_u9652_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9653 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [14]),
    .o(_al_u9653_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9654 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [14]),
    .o(_al_u9654_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9655 (
    .a(_al_u9651_o),
    .b(_al_u9652_o),
    .c(_al_u9653_o),
    .d(_al_u9654_o),
    .o(_al_u9655_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9656 (
    .a(_al_u9650_o),
    .b(_al_u9655_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9657 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [11]),
    .d(addr_if[13]),
    .o(_al_u9657_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9658 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [15]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [11]),
    .o(_al_u9658_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9659 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[13]),
    .o(_al_u9659_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9660 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [13]),
    .o(_al_u9660_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9661 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [13]),
    .o(_al_u9661_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9662 (
    .a(_al_u9658_o),
    .b(_al_u9659_o),
    .c(_al_u9660_o),
    .d(_al_u9661_o),
    .o(_al_u9662_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9663 (
    .a(_al_u9657_o),
    .b(_al_u9662_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9664 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [10]),
    .d(addr_if[12]),
    .o(_al_u9664_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u9665 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [14]),
    .c(\cu_ru/n43 [10]),
    .o(_al_u9665_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u9666 (
    .a(_al_u9665_o),
    .b(_al_u6055_o),
    .c(_al_u2842_o),
    .d(new_pc[12]),
    .o(_al_u9666_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(D)*~(A)+(C*B)*D*~(A)+~((C*B))*D*A+(C*B)*D*A)"),
    .INIT(16'h15bf))
    _al_u9667 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [12]),
    .d(\cu_ru/mepc [12]),
    .o(_al_u9667_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u9668 (
    .a(_al_u9664_o),
    .b(_al_u9666_o),
    .c(pip_flush),
    .d(_al_u9667_o),
    .o(\ins_fetch/n4 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u9669 (
    .a(\ins_fetch/n27 ),
    .b(pip_flush),
    .c(\ins_fetch/n1 [0]),
    .d(addr_if[2]),
    .o(_al_u9669_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .INIT(16'h010b))
    _al_u9670 (
    .a(\cu_ru/mux34_b0_sel_is_2_o ),
    .b(\cu_ru/tvec [4]),
    .c(_al_u6055_o),
    .d(\cu_ru/n43 [0]),
    .o(_al_u9670_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*A))"),
    .INIT(8'h31))
    _al_u9671 (
    .a(_al_u6055_o),
    .b(_al_u2844_o),
    .c(new_pc[2]),
    .o(_al_u9671_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9672 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(\cu_ru/mepc [2]),
    .o(_al_u9672_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9673 (
    .a(\cu_ru/m_s_status/n2 ),
    .b(_al_u2844_o),
    .c(\cu_ru/sepc [2]),
    .o(_al_u9673_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B*~A)))"),
    .INIT(16'h040f))
    _al_u9674 (
    .a(_al_u9670_o),
    .b(_al_u9671_o),
    .c(_al_u9672_o),
    .d(_al_u9673_o),
    .o(_al_u9674_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u9675 (
    .a(_al_u9669_o),
    .b(_al_u9674_o),
    .c(pip_flush),
    .o(\ins_fetch/n4 [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u9676 (
    .a(_al_u9204_o),
    .b(_al_u9264_o),
    .c(\biu/cache_ctrl_logic/n55_lutinv ),
    .o(_al_u9676_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9677 (
    .a(_al_u7149_o),
    .b(_al_u3950_o),
    .o(_al_u9677_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~C*~A))"),
    .INIT(16'h3233))
    _al_u9678 (
    .a(_al_u3947_o),
    .b(_al_u3950_o),
    .c(_al_u7151_o),
    .d(\biu/cache_ctrl_logic/statu [0]),
    .o(_al_u9678_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D*A)))"),
    .INIT(16'h2303))
    _al_u9679 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u9677_o),
    .c(_al_u9678_o),
    .d(_al_u3947_o),
    .o(_al_u9679_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u9680 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/n204_lutinv ),
    .o(_al_u9680_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9681 (
    .a(_al_u7149_o),
    .b(\biu/cache_ctrl_logic/n97_lutinv ),
    .o(_al_u9681_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*~A))"),
    .INIT(16'hf0e0))
    _al_u9682 (
    .a(_al_u9272_o),
    .b(_al_u9679_o),
    .c(_al_u9680_o),
    .d(_al_u9681_o),
    .o(_al_u9682_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9683 (
    .a(_al_u9682_o),
    .b(\biu/cache_ctrl_logic/n100 [4]),
    .c(_al_u4834_o),
    .o(_al_u9683_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u9684 (
    .a(_al_u7190_o),
    .b(read),
    .c(\biu/cache_ctrl_logic/n100 [4]),
    .o(\biu/cache_ctrl_logic/n83 [0]));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u9685 (
    .a(\biu/cache_ctrl_logic/n83 [0]),
    .b(_al_u7157_o),
    .c(\biu/cache_ctrl_logic/n75_lutinv ),
    .d(write),
    .o(_al_u9685_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9686 (
    .a(_al_u7149_o),
    .b(write),
    .o(_al_u9686_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(D*~A)))"),
    .INIT(16'h0703))
    _al_u9687 (
    .a(_al_u9686_o),
    .b(\biu/cache_ctrl_logic/l1d_wr_sel_lutinv ),
    .c(\biu/cache_ctrl_logic/n75_lutinv ),
    .d(\biu/cache_ctrl_logic/n100 [4]),
    .o(_al_u9687_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*C*~A))"),
    .INIT(16'h3323))
    _al_u9688 (
    .a(_al_u9683_o),
    .b(_al_u9685_o),
    .c(_al_u9687_o),
    .d(_al_u2848_o),
    .o(_al_u9688_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9689 (
    .a(_al_u7190_o),
    .b(_al_u7191_o),
    .o(_al_u9689_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd0d5))
    _al_u9690 (
    .a(_al_u9689_o),
    .b(\biu/cache_ctrl_logic/n100 [4]),
    .c(_al_u7149_o),
    .d(_al_u2886_o),
    .o(_al_u9690_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9691 (
    .a(_al_u9690_o),
    .b(_al_u7162_o),
    .o(_al_u9691_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*A))"),
    .INIT(16'h0007))
    _al_u9692 (
    .a(_al_u9688_o),
    .b(_al_u9691_o),
    .c(_al_u9286_o),
    .d(_al_u7193_o),
    .o(_al_u9692_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u9693 (
    .a(_al_u9283_o),
    .b(\exu/c_fence_lutinv ),
    .c(\biu/cache_ctrl_logic/n55_lutinv ),
    .d(cache_flush),
    .o(_al_u9693_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(~A*~(~C*~B)))"),
    .INIT(16'h54ff))
    _al_u9694 (
    .a(_al_u9676_o),
    .b(_al_u9692_o),
    .c(_al_u9285_o),
    .d(_al_u9693_o),
    .o(\biu/cache_ctrl_logic/n132[0]_d ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u9695 (
    .a(_al_u9273_o),
    .b(_al_u9274_o),
    .c(\biu/cache_ctrl_logic/statu [2]),
    .o(_al_u9695_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(C*~B)))"),
    .INIT(16'haa20))
    _al_u9696 (
    .a(_al_u9271_o),
    .b(_al_u9272_o),
    .c(_al_u9695_o),
    .d(_al_u4399_o),
    .o(_al_u9696_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u9697 (
    .a(_al_u9278_o),
    .b(\biu/cache_ctrl_logic/n100 [4]),
    .o(_al_u9697_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9698 (
    .a(_al_u7149_o),
    .b(_al_u3224_o),
    .o(_al_u9698_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u9699 (
    .a(_al_u9696_o),
    .b(_al_u9697_o),
    .c(_al_u9698_o),
    .o(_al_u9699_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u9700 (
    .a(_al_u9699_o),
    .b(_al_u9280_o),
    .c(_al_u7159_o),
    .d(_al_u2886_o),
    .o(_al_u9700_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u9701 (
    .a(_al_u7163_o),
    .b(_al_u2885_o),
    .o(_al_u9701_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(~C*~A)))"),
    .INIT(16'hcc04))
    _al_u9702 (
    .a(_al_u9700_o),
    .b(_al_u7192_o),
    .c(_al_u9701_o),
    .d(\biu/bus_unit/mmu/n19_lutinv ),
    .o(_al_u9702_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*A*~(~D*~B))"),
    .INIT(16'h5f7f))
    _al_u9703 (
    .a(_al_u9284_o),
    .b(_al_u9702_o),
    .c(_al_u9287_o),
    .d(_al_u7193_o),
    .o(\biu/cache_ctrl_logic/n132 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9704 (
    .a(_al_u7151_o),
    .b(\biu/cache_ctrl_logic/statu [1]),
    .o(_al_u9704_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u9705 (
    .a(_al_u7149_o),
    .b(_al_u9704_o),
    .c(_al_u3947_o),
    .o(_al_u9705_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u9706 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u9705_o),
    .c(_al_u3950_o),
    .o(_al_u9706_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u9707 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(_al_u4399_o),
    .c(\biu/cache_ctrl_logic/l1i_pte [7]),
    .o(_al_u9707_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u9708 (
    .a(\biu/cache_ctrl_logic/n100 [4]),
    .b(\biu/cache_ctrl_logic/n75_lutinv ),
    .c(\biu/cache_ctrl_logic/n204_lutinv ),
    .o(_al_u9708_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(~D*~A))"),
    .INIT(16'h3020))
    _al_u9709 (
    .a(_al_u9706_o),
    .b(_al_u9707_o),
    .c(_al_u9708_o),
    .d(_al_u9681_o),
    .o(_al_u9709_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u9710 (
    .a(_al_u7163_o),
    .b(_al_u2885_o),
    .o(_al_u9710_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(~C*~A)))"),
    .INIT(16'h00cd))
    _al_u9711 (
    .a(_al_u9709_o),
    .b(_al_u9710_o),
    .c(_al_u7158_o),
    .d(\biu/bus_unit/mmu/n19_lutinv ),
    .o(_al_u9711_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~C*~A))"),
    .INIT(16'h3332))
    _al_u9712 (
    .a(_al_u9711_o),
    .b(_al_u7162_o),
    .c(_al_u9689_o),
    .d(_al_u2848_o),
    .o(_al_u9712_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcd0d))
    _al_u9713 (
    .a(_al_u9712_o),
    .b(_al_u9286_o),
    .c(_al_u7193_o),
    .d(\biu/cache_ctrl_logic/l1d_pte [7]),
    .o(_al_u9713_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B*~A))"),
    .INIT(8'h4f))
    _al_u9714 (
    .a(_al_u9676_o),
    .b(_al_u9713_o),
    .c(_al_u9693_o),
    .o(\biu/cache_ctrl_logic/n131[1]_d ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u9715 (
    .a(_al_u9284_o),
    .b(_al_u9287_o),
    .c(\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/mux44_b4_sel_is_2_o ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u9716 (
    .a(\biu/bus_unit/mmu/i [0]),
    .o(\biu/bus_unit/mmu/n59 [0]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u9717 (
    .a(if_hold),
    .o(_al_n0_en));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add0/u0  (
    .a(\biu/bus_unit/addr_counter [0]),
    .b(1'b1),
    .c(\biu/bus_unit/add0/c0 ),
    .o({\biu/bus_unit/add0/c1 ,\biu/bus_unit/n39 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add0/u1  (
    .a(\biu/bus_unit/addr_counter [1]),
    .b(1'b0),
    .c(\biu/bus_unit/add0/c1 ),
    .o({\biu/bus_unit/add0/c2 ,\biu/bus_unit/n39 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add0/u2  (
    .a(\biu/bus_unit/addr_counter [2]),
    .b(1'b0),
    .c(\biu/bus_unit/add0/c2 ),
    .o({\biu/bus_unit/add0/c3 ,\biu/bus_unit/n39 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add0/u3  (
    .a(\biu/bus_unit/addr_counter [3]),
    .b(1'b0),
    .c(\biu/bus_unit/add0/c3 ),
    .o({\biu/bus_unit/add0/c4 ,\biu/bus_unit/n39 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add0/u4  (
    .a(\biu/bus_unit/addr_counter [4]),
    .b(1'b0),
    .c(\biu/bus_unit/add0/c4 ),
    .o({\biu/bus_unit/add0/c5 ,\biu/bus_unit/n39 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add0/u5  (
    .a(\biu/bus_unit/addr_counter [5]),
    .b(1'b0),
    .c(\biu/bus_unit/add0/c5 ),
    .o({\biu/bus_unit/add0/c6 ,\biu/bus_unit/n39 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add0/u6  (
    .a(\biu/bus_unit/addr_counter [6]),
    .b(1'b0),
    .c(\biu/bus_unit/add0/c6 ),
    .o({\biu/bus_unit/add0/c7 ,\biu/bus_unit/n39 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add0/u7  (
    .a(\biu/bus_unit/addr_counter [7]),
    .b(1'b0),
    .c(\biu/bus_unit/add0/c7 ),
    .o({\biu/bus_unit/add0/c8 ,\biu/bus_unit/n39 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add0/u8  (
    .a(\biu/bus_unit/addr_counter [8]),
    .b(1'b0),
    .c(\biu/bus_unit/add0/c8 ),
    .o({open_n5237,\biu/bus_unit/n39 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \biu/bus_unit/add0/ucin  (
    .a(1'b0),
    .o({\biu/bus_unit/add0/c0 ,open_n5240}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u0  (
    .a(\biu/bus_unit/addr_counter [0]),
    .b(\biu/maddress [3]),
    .c(\biu/bus_unit/add1/c0 ),
    .o({\biu/bus_unit/add1/c1 ,\biu/bus_unit/n49 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u1  (
    .a(\biu/bus_unit/addr_counter [1]),
    .b(\biu/maddress [4]),
    .c(\biu/bus_unit/add1/c1 ),
    .o({\biu/bus_unit/add1/c2 ,\biu/bus_unit/n49 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u10  (
    .a(1'b0),
    .b(\biu/maddress [13]),
    .c(\biu/bus_unit/add1/c10 ),
    .o({\biu/bus_unit/add1/c11 ,\biu/bus_unit/n49 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u11  (
    .a(1'b0),
    .b(\biu/maddress [14]),
    .c(\biu/bus_unit/add1/c11 ),
    .o({\biu/bus_unit/add1/c12 ,\biu/bus_unit/n49 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u12  (
    .a(1'b0),
    .b(\biu/maddress [15]),
    .c(\biu/bus_unit/add1/c12 ),
    .o({\biu/bus_unit/add1/c13 ,\biu/bus_unit/n49 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u13  (
    .a(1'b0),
    .b(\biu/maddress [16]),
    .c(\biu/bus_unit/add1/c13 ),
    .o({\biu/bus_unit/add1/c14 ,\biu/bus_unit/n49 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u14  (
    .a(1'b0),
    .b(\biu/maddress [17]),
    .c(\biu/bus_unit/add1/c14 ),
    .o({\biu/bus_unit/add1/c15 ,\biu/bus_unit/n49 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u15  (
    .a(1'b0),
    .b(\biu/maddress [18]),
    .c(\biu/bus_unit/add1/c15 ),
    .o({\biu/bus_unit/add1/c16 ,\biu/bus_unit/n49 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u16  (
    .a(1'b0),
    .b(\biu/maddress [19]),
    .c(\biu/bus_unit/add1/c16 ),
    .o({\biu/bus_unit/add1/c17 ,\biu/bus_unit/n49 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u17  (
    .a(1'b0),
    .b(\biu/maddress [20]),
    .c(\biu/bus_unit/add1/c17 ),
    .o({\biu/bus_unit/add1/c18 ,\biu/bus_unit/n49 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u18  (
    .a(1'b0),
    .b(\biu/maddress [21]),
    .c(\biu/bus_unit/add1/c18 ),
    .o({\biu/bus_unit/add1/c19 ,\biu/bus_unit/n49 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u19  (
    .a(1'b0),
    .b(\biu/maddress [22]),
    .c(\biu/bus_unit/add1/c19 ),
    .o({\biu/bus_unit/add1/c20 ,\biu/bus_unit/n49 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u2  (
    .a(\biu/bus_unit/addr_counter [2]),
    .b(\biu/maddress [5]),
    .c(\biu/bus_unit/add1/c2 ),
    .o({\biu/bus_unit/add1/c3 ,\biu/bus_unit/n49 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u20  (
    .a(1'b0),
    .b(\biu/maddress [23]),
    .c(\biu/bus_unit/add1/c20 ),
    .o({\biu/bus_unit/add1/c21 ,\biu/bus_unit/n49 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u21  (
    .a(1'b0),
    .b(\biu/maddress [24]),
    .c(\biu/bus_unit/add1/c21 ),
    .o({\biu/bus_unit/add1/c22 ,\biu/bus_unit/n49 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u22  (
    .a(1'b0),
    .b(\biu/maddress [25]),
    .c(\biu/bus_unit/add1/c22 ),
    .o({\biu/bus_unit/add1/c23 ,\biu/bus_unit/n49 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u23  (
    .a(1'b0),
    .b(\biu/maddress [26]),
    .c(\biu/bus_unit/add1/c23 ),
    .o({\biu/bus_unit/add1/c24 ,\biu/bus_unit/n49 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u24  (
    .a(1'b0),
    .b(\biu/maddress [27]),
    .c(\biu/bus_unit/add1/c24 ),
    .o({\biu/bus_unit/add1/c25 ,\biu/bus_unit/n49 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u25  (
    .a(1'b0),
    .b(\biu/maddress [28]),
    .c(\biu/bus_unit/add1/c25 ),
    .o({\biu/bus_unit/add1/c26 ,\biu/bus_unit/n49 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u26  (
    .a(1'b0),
    .b(\biu/maddress [29]),
    .c(\biu/bus_unit/add1/c26 ),
    .o({\biu/bus_unit/add1/c27 ,\biu/bus_unit/n49 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u27  (
    .a(1'b0),
    .b(\biu/maddress [30]),
    .c(\biu/bus_unit/add1/c27 ),
    .o({\biu/bus_unit/add1/c28 ,\biu/bus_unit/n49 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u28  (
    .a(1'b0),
    .b(\biu/maddress [31]),
    .c(\biu/bus_unit/add1/c28 ),
    .o({\biu/bus_unit/add1/c29 ,\biu/bus_unit/n49 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u29  (
    .a(1'b0),
    .b(\biu/maddress [32]),
    .c(\biu/bus_unit/add1/c29 ),
    .o({\biu/bus_unit/add1/c30 ,\biu/bus_unit/n49 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u3  (
    .a(\biu/bus_unit/addr_counter [3]),
    .b(\biu/maddress [6]),
    .c(\biu/bus_unit/add1/c3 ),
    .o({\biu/bus_unit/add1/c4 ,\biu/bus_unit/n49 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u30  (
    .a(1'b0),
    .b(\biu/maddress [33]),
    .c(\biu/bus_unit/add1/c30 ),
    .o({\biu/bus_unit/add1/c31 ,\biu/bus_unit/n49 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u31  (
    .a(1'b0),
    .b(\biu/maddress [34]),
    .c(\biu/bus_unit/add1/c31 ),
    .o({\biu/bus_unit/add1/c32 ,\biu/bus_unit/n49 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u32  (
    .a(1'b0),
    .b(\biu/maddress [35]),
    .c(\biu/bus_unit/add1/c32 ),
    .o({\biu/bus_unit/add1/c33 ,\biu/bus_unit/n49 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u33  (
    .a(1'b0),
    .b(\biu/maddress [36]),
    .c(\biu/bus_unit/add1/c33 ),
    .o({\biu/bus_unit/add1/c34 ,\biu/bus_unit/n49 [33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u34  (
    .a(1'b0),
    .b(\biu/maddress [37]),
    .c(\biu/bus_unit/add1/c34 ),
    .o({\biu/bus_unit/add1/c35 ,\biu/bus_unit/n49 [34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u35  (
    .a(1'b0),
    .b(\biu/maddress [38]),
    .c(\biu/bus_unit/add1/c35 ),
    .o({\biu/bus_unit/add1/c36 ,\biu/bus_unit/n49 [35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u36  (
    .a(1'b0),
    .b(\biu/maddress [39]),
    .c(\biu/bus_unit/add1/c36 ),
    .o({\biu/bus_unit/add1/c37 ,\biu/bus_unit/n49 [36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u37  (
    .a(1'b0),
    .b(\biu/maddress [40]),
    .c(\biu/bus_unit/add1/c37 ),
    .o({\biu/bus_unit/add1/c38 ,\biu/bus_unit/n49 [37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u38  (
    .a(1'b0),
    .b(\biu/maddress [41]),
    .c(\biu/bus_unit/add1/c38 ),
    .o({\biu/bus_unit/add1/c39 ,\biu/bus_unit/n49 [38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u39  (
    .a(1'b0),
    .b(\biu/maddress [42]),
    .c(\biu/bus_unit/add1/c39 ),
    .o({\biu/bus_unit/add1/c40 ,\biu/bus_unit/n49 [39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u4  (
    .a(\biu/bus_unit/addr_counter [4]),
    .b(\biu/maddress [7]),
    .c(\biu/bus_unit/add1/c4 ),
    .o({\biu/bus_unit/add1/c5 ,\biu/bus_unit/n49 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u40  (
    .a(1'b0),
    .b(\biu/maddress [43]),
    .c(\biu/bus_unit/add1/c40 ),
    .o({\biu/bus_unit/add1/c41 ,\biu/bus_unit/n49 [40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u41  (
    .a(1'b0),
    .b(\biu/maddress [44]),
    .c(\biu/bus_unit/add1/c41 ),
    .o({\biu/bus_unit/add1/c42 ,\biu/bus_unit/n49 [41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u42  (
    .a(1'b0),
    .b(\biu/maddress [45]),
    .c(\biu/bus_unit/add1/c42 ),
    .o({\biu/bus_unit/add1/c43 ,\biu/bus_unit/n49 [42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u43  (
    .a(1'b0),
    .b(\biu/maddress [46]),
    .c(\biu/bus_unit/add1/c43 ),
    .o({\biu/bus_unit/add1/c44 ,\biu/bus_unit/n49 [43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u44  (
    .a(1'b0),
    .b(\biu/maddress [47]),
    .c(\biu/bus_unit/add1/c44 ),
    .o({\biu/bus_unit/add1/c45 ,\biu/bus_unit/n49 [44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u45  (
    .a(1'b0),
    .b(\biu/maddress [48]),
    .c(\biu/bus_unit/add1/c45 ),
    .o({\biu/bus_unit/add1/c46 ,\biu/bus_unit/n49 [45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u46  (
    .a(1'b0),
    .b(\biu/maddress [49]),
    .c(\biu/bus_unit/add1/c46 ),
    .o({\biu/bus_unit/add1/c47 ,\biu/bus_unit/n49 [46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u47  (
    .a(1'b0),
    .b(\biu/maddress [50]),
    .c(\biu/bus_unit/add1/c47 ),
    .o({\biu/bus_unit/add1/c48 ,\biu/bus_unit/n49 [47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u48  (
    .a(1'b0),
    .b(\biu/maddress [51]),
    .c(\biu/bus_unit/add1/c48 ),
    .o({\biu/bus_unit/add1/c49 ,\biu/bus_unit/n49 [48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u49  (
    .a(1'b0),
    .b(\biu/maddress [52]),
    .c(\biu/bus_unit/add1/c49 ),
    .o({\biu/bus_unit/add1/c50 ,\biu/bus_unit/n49 [49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u5  (
    .a(\biu/bus_unit/addr_counter [5]),
    .b(\biu/maddress [8]),
    .c(\biu/bus_unit/add1/c5 ),
    .o({\biu/bus_unit/add1/c6 ,\biu/bus_unit/n49 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u50  (
    .a(1'b0),
    .b(\biu/maddress [53]),
    .c(\biu/bus_unit/add1/c50 ),
    .o({\biu/bus_unit/add1/c51 ,\biu/bus_unit/n49 [50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u51  (
    .a(1'b0),
    .b(\biu/maddress [54]),
    .c(\biu/bus_unit/add1/c51 ),
    .o({\biu/bus_unit/add1/c52 ,\biu/bus_unit/n49 [51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u52  (
    .a(1'b0),
    .b(\biu/maddress [55]),
    .c(\biu/bus_unit/add1/c52 ),
    .o({\biu/bus_unit/add1/c53 ,\biu/bus_unit/n49 [52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u53  (
    .a(1'b0),
    .b(\biu/maddress [56]),
    .c(\biu/bus_unit/add1/c53 ),
    .o({\biu/bus_unit/add1/c54 ,\biu/bus_unit/n49 [53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u54  (
    .a(1'b0),
    .b(\biu/maddress [57]),
    .c(\biu/bus_unit/add1/c54 ),
    .o({\biu/bus_unit/add1/c55 ,\biu/bus_unit/n49 [54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u55  (
    .a(1'b0),
    .b(\biu/maddress [58]),
    .c(\biu/bus_unit/add1/c55 ),
    .o({\biu/bus_unit/add1/c56 ,\biu/bus_unit/n49 [55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u56  (
    .a(1'b0),
    .b(\biu/maddress [59]),
    .c(\biu/bus_unit/add1/c56 ),
    .o({\biu/bus_unit/add1/c57 ,\biu/bus_unit/n49 [56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u57  (
    .a(1'b0),
    .b(\biu/maddress [60]),
    .c(\biu/bus_unit/add1/c57 ),
    .o({\biu/bus_unit/add1/c58 ,\biu/bus_unit/n49 [57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u58  (
    .a(1'b0),
    .b(\biu/maddress [61]),
    .c(\biu/bus_unit/add1/c58 ),
    .o({\biu/bus_unit/add1/c59 ,\biu/bus_unit/n49 [58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u59  (
    .a(1'b0),
    .b(\biu/maddress [62]),
    .c(\biu/bus_unit/add1/c59 ),
    .o({\biu/bus_unit/add1/c60 ,\biu/bus_unit/n49 [59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u6  (
    .a(\biu/bus_unit/addr_counter [6]),
    .b(\biu/maddress [9]),
    .c(\biu/bus_unit/add1/c6 ),
    .o({\biu/bus_unit/add1/c7 ,\biu/bus_unit/n49 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u60  (
    .a(1'b0),
    .b(\biu/maddress [63]),
    .c(\biu/bus_unit/add1/c60 ),
    .o({open_n5241,\biu/bus_unit/n49 [60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u7  (
    .a(\biu/bus_unit/addr_counter [7]),
    .b(\biu/maddress [10]),
    .c(\biu/bus_unit/add1/c7 ),
    .o({\biu/bus_unit/add1/c8 ,\biu/bus_unit/n49 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u8  (
    .a(\biu/bus_unit/addr_counter [8]),
    .b(\biu/maddress [11]),
    .c(\biu/bus_unit/add1/c8 ),
    .o({\biu/bus_unit/add1/c9 ,\biu/bus_unit/n49 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/bus_unit/add1/u9  (
    .a(1'b0),
    .b(\biu/maddress [12]),
    .c(\biu/bus_unit/add1/c9 ),
    .o({\biu/bus_unit/add1/c10 ,\biu/bus_unit/n49 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \biu/bus_unit/add1/ucin  (
    .a(1'b0),
    .o({\biu/bus_unit/add1/c0 ,open_n5244}));
  reg_sr_as_w1 \biu/bus_unit/mmu/reg0_b0  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n59 [0]),
    .en(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/mmu/n58 ),
    .set(1'b0),
    .q(\biu/bus_unit/mmu/i [0]));  // ../../RTL/CPU/BIU/mmu.v(166)
  reg_ar_ss_w1 \biu/bus_unit/mmu/reg0_b1  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n59 [1]),
    .en(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(\biu/bus_unit/mmu/n58 ),
    .q(\biu/bus_unit/mmu/i [1]));  // ../../RTL/CPU/BIU/mmu.v(166)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b0  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [0]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b1  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [1]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b10  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [10]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b11  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [11]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b12  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [12]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b13  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [13]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b14  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [14]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b15  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [15]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b16  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [16]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b17  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [17]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b18  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [18]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b19  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [19]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b2  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [2]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b20  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [20]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b21  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [21]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b22  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [22]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b23  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [23]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b24  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [24]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b25  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [25]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b26  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [26]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b27  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [27]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b28  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [28]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b29  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [29]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b3  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [3]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b30  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [30]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b31  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [31]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b32  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [32]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b33  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [33]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b34  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [34]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b35  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [35]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b36  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [36]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b37  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [37]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b38  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [38]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b39  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [39]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b4  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [4]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b40  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [40]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b41  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [41]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b42  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [42]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b43  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [43]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b44  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [44]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b45  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [45]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b46  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [46]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b47  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [47]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b48  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [48]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b49  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [49]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b5  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [5]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b50  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [50]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b51  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [51]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b52  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [52]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b53  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [53]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b54  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [54]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b55  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [55]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b56  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [56]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b57  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [57]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b58  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [58]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b59  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [59]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b6  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [6]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b60  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [60]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b61  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [61]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b62  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [62]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b63  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [63]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b7  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [7]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b8  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [8]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b9  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n66 [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [9]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b0  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [64]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b1  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [65]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b10  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [74]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b11  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [75]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b12  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [76]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b13  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [77]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b14  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [78]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b15  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [79]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b16  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [80]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b17  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [81]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b18  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [82]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b19  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [83]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b2  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [66]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b20  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [84]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b21  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [85]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b22  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [86]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b23  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [87]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b24  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [88]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b25  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [89]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b26  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [90]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b27  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [91]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b28  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [92]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b29  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [93]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b3  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [67]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b30  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [94]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b31  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [95]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b32  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [96]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b33  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [97]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b34  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [98]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b35  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [99]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b36  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [100]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b37  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [101]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b38  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [102]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b39  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [103]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b4  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [68]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b40  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [104]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b41  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [105]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b42  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [106]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b43  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [107]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b44  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [108]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b45  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [109]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b46  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [110]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b47  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [111]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b48  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [112]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b49  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [113]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b5  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [69]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b50  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [114]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b51  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [115]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b52  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [116]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b53  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [117]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b54  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [118]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b55  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [119]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b56  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [120]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b57  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [121]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b58  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [122]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b59  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [123]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b6  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [70]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b60  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [124]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b61  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [125]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b62  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [126]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b63  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [127]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b7  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [71]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b8  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [72]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b9  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n71 [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/paddress [73]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b0  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [0]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b1  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [1]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b10  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [10]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b11  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [11]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b12  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [12]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b13  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [13]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b14  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [14]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b15  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [15]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b16  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [16]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b17  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [17]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b18  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [18]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b19  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [19]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b2  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [2]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b20  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [20]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b21  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [21]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b22  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [22]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b23  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [23]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b24  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [24]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b25  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [25]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b26  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [26]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b27  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [27]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b28  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [28]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b29  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [29]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b3  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [3]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b30  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [30]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b31  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [31]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b32  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [32]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b33  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [33]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b34  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [34]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b35  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [35]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b36  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [36]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b37  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [37]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b38  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [38]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b39  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [39]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b4  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [4]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b40  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [40]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b41  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [41]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b42  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [42]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b43  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [43]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b44  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [44]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b45  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [45]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b46  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [46]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b47  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [47]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b48  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [48]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b49  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [49]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b5  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [5]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b50  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [50]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b51  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [51]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b52  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [52]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b53  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [53]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b54  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [54]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b55  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [55]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b56  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [56]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b57  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [57]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b58  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [58]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b59  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [59]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b6  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [6]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b60  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [60]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b61  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [61]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b62  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [62]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b63  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [63]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b7  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [7]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b8  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [8]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b9  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n79 [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [9]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg4_b0  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n56 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu/statu [0]));  // ../../RTL/CPU/BIU/mmu.v(154)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg4_b1  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n56 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu/statu [1]));  // ../../RTL/CPU/BIU/mmu.v(154)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg4_b2  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n56 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/mmu/statu [2]));  // ../../RTL/CPU/BIU/mmu.v(154)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg4_b3  (
    .clk(clk_pad),
    .d(\biu/bus_unit/mmu/n54 [3]),
    .en(1'b1),
    .reset(~\biu/bus_unit/mmu/mux18_b3_sel_is_2_o ),
    .set(1'b0),
    .q(\biu/bus_unit/mmu/statu [3]));  // ../../RTL/CPU/BIU/mmu.v(154)
  reg_sr_as_w1 \biu/bus_unit/reg0_b0  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n39[0]_d ),
    .en(\biu/bus_unit/n39[0]_en ),
    .reset(\biu/bus_unit/n37 ),
    .set(1'b0),
    .q(\biu/bus_unit/addr_counter [0]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_as_w1 \biu/bus_unit/reg0_b1  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n39[1]_d ),
    .en(\biu/bus_unit/n39[0]_en ),
    .reset(\biu/bus_unit/n37 ),
    .set(1'b0),
    .q(\biu/bus_unit/addr_counter [1]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_as_w1 \biu/bus_unit/reg0_b2  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n39[2]_d ),
    .en(\biu/bus_unit/n39[0]_en ),
    .reset(\biu/bus_unit/n37 ),
    .set(1'b0),
    .q(\biu/bus_unit/addr_counter [2]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_as_w1 \biu/bus_unit/reg0_b3  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n39[3]_d ),
    .en(\biu/bus_unit/n39[0]_en ),
    .reset(\biu/bus_unit/n37 ),
    .set(1'b0),
    .q(\biu/bus_unit/addr_counter [3]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_as_w1 \biu/bus_unit/reg0_b4  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n39[4]_d ),
    .en(\biu/bus_unit/n39[0]_en ),
    .reset(\biu/bus_unit/n37 ),
    .set(1'b0),
    .q(\biu/bus_unit/addr_counter [4]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_as_w1 \biu/bus_unit/reg0_b5  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n39[5]_d ),
    .en(\biu/bus_unit/n39[0]_en ),
    .reset(\biu/bus_unit/n37 ),
    .set(1'b0),
    .q(\biu/bus_unit/addr_counter [5]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_as_w1 \biu/bus_unit/reg0_b6  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n39[6]_d ),
    .en(\biu/bus_unit/n39[0]_en ),
    .reset(\biu/bus_unit/n37 ),
    .set(1'b0),
    .q(\biu/bus_unit/addr_counter [6]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_as_w1 \biu/bus_unit/reg0_b7  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n39[7]_d ),
    .en(\biu/bus_unit/n39[0]_en ),
    .reset(\biu/bus_unit/n37 ),
    .set(1'b0),
    .q(\biu/bus_unit/addr_counter [7]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_as_w1 \biu/bus_unit/reg0_b8  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n39[8]_d ),
    .en(\biu/bus_unit/n39[0]_en ),
    .reset(\biu/bus_unit/n37 ),
    .set(1'b0),
    .q(\biu/bus_unit/addr_counter [8]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_as_w1 \biu/bus_unit/reg1_b0  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n35 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/statu [0]));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  reg_sr_as_w1 \biu/bus_unit/reg1_b1  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n35 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/statu [1]));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  reg_sr_as_w1 \biu/bus_unit/reg1_b2  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n35 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/statu [2]));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  reg_sr_as_w1 \biu/bus_unit/reg1_b3  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n35 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/bus_unit/statu [3]));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  reg_sr_as_w1 \biu/bus_unit/reg1_b4  (
    .clk(clk_pad),
    .d(\biu/bus_unit/n30 [4]),
    .en(1'b1),
    .reset(~\biu/bus_unit/mux17_b4_sel_is_2_o ),
    .set(1'b0),
    .q(\biu/bus_unit/statu [4]));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \biu/bus_unit/sub0/u0  (
    .a(\biu/bus_unit/addr_counter [0]),
    .b(1'b1),
    .c(\biu/bus_unit/sub0/c0 ),
    .o({\biu/bus_unit/sub0/c1 ,\biu/bus_unit/last_addr [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \biu/bus_unit/sub0/u1  (
    .a(\biu/bus_unit/addr_counter [1]),
    .b(1'b0),
    .c(\biu/bus_unit/sub0/c1 ),
    .o({\biu/bus_unit/sub0/c2 ,\biu/bus_unit/last_addr [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \biu/bus_unit/sub0/u2  (
    .a(\biu/bus_unit/addr_counter [2]),
    .b(1'b0),
    .c(\biu/bus_unit/sub0/c2 ),
    .o({\biu/bus_unit/sub0/c3 ,\biu/bus_unit/last_addr [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \biu/bus_unit/sub0/u3  (
    .a(\biu/bus_unit/addr_counter [3]),
    .b(1'b0),
    .c(\biu/bus_unit/sub0/c3 ),
    .o({\biu/bus_unit/sub0/c4 ,\biu/bus_unit/last_addr [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \biu/bus_unit/sub0/u4  (
    .a(\biu/bus_unit/addr_counter [4]),
    .b(1'b0),
    .c(\biu/bus_unit/sub0/c4 ),
    .o({\biu/bus_unit/sub0/c5 ,\biu/bus_unit/last_addr [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \biu/bus_unit/sub0/u5  (
    .a(\biu/bus_unit/addr_counter [5]),
    .b(1'b0),
    .c(\biu/bus_unit/sub0/c5 ),
    .o({\biu/bus_unit/sub0/c6 ,\biu/bus_unit/last_addr [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \biu/bus_unit/sub0/u6  (
    .a(\biu/bus_unit/addr_counter [6]),
    .b(1'b0),
    .c(\biu/bus_unit/sub0/c6 ),
    .o({\biu/bus_unit/sub0/c7 ,\biu/bus_unit/last_addr [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \biu/bus_unit/sub0/u7  (
    .a(\biu/bus_unit/addr_counter [7]),
    .b(1'b0),
    .c(\biu/bus_unit/sub0/c7 ),
    .o({\biu/bus_unit/sub0/c8 ,\biu/bus_unit/last_addr [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \biu/bus_unit/sub0/u8  (
    .a(\biu/bus_unit/addr_counter [8]),
    .b(1'b0),
    .c(\biu/bus_unit/sub0/c8 ),
    .o({open_n5245,\biu/bus_unit/last_addr [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \biu/bus_unit/sub0/ucin  (
    .a(1'b0),
    .o({\biu/bus_unit/sub0/c0 ,open_n5248}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d00_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5271,\biu/l1i_in [7:0]}),
    .wea(\biu/cache/n1 ),
    .doa({open_n5286,\biu/l1d_out [7:0]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d10_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5318,\biu/l1i_in [15:8]}),
    .wea(\biu/cache/n3 ),
    .doa({open_n5333,\biu/l1d_out [15:8]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d20_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5365,\biu/l1i_in [23:16]}),
    .wea(\biu/cache/n5 ),
    .doa({open_n5380,\biu/l1d_out [23:16]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d30_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5412,\biu/l1i_in [31:24]}),
    .wea(\biu/cache/n7 ),
    .doa({open_n5427,\biu/l1d_out [31:24]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d40_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5459,\biu/l1i_in [39:32]}),
    .wea(\biu/cache/n9 ),
    .doa({open_n5474,\biu/l1d_out [39:32]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d50_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5506,\biu/l1i_in [47:40]}),
    .wea(\biu/cache/n11 ),
    .doa({open_n5521,\biu/l1d_out [47:40]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d60_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5553,\biu/l1i_in [55:48]}),
    .wea(\biu/cache/n13 ),
    .doa({open_n5568,\biu/l1d_out [55:48]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d70_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1d_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5600,\biu/l1i_in [63:56]}),
    .wea(\biu/cache/n15 ),
    .doa({open_n5615,\biu/l1d_out [63:56]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i00_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5647,\biu/l1i_in [7:0]}),
    .wea(\biu/cache/n17 ),
    .doa({open_n5662,ins_read[7:0]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i10_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5694,\biu/l1i_in [15:8]}),
    .wea(\biu/cache/n19 ),
    .doa({open_n5709,ins_read[15:8]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i20_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5741,\biu/l1i_in [23:16]}),
    .wea(\biu/cache/n21 ),
    .doa({open_n5756,ins_read[23:16]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i30_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5788,\biu/l1i_in [31:24]}),
    .wea(\biu/cache/n23 ),
    .doa({open_n5803,ins_read[31:24]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i40_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5835,\biu/l1i_in [39:32]}),
    .wea(\biu/cache/n25 ),
    .doa({open_n5850,ins_read[39:32]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i50_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5882,\biu/l1i_in [47:40]}),
    .wea(\biu/cache/n27 ),
    .doa({open_n5897,ins_read[47:40]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i60_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5929,\biu/l1i_in [55:48]}),
    .wea(\biu/cache/n29 ),
    .doa({open_n5944,ins_read[55:48]}));
  // address_offset=0;data_offset=0;depth=512;width=8;num_section=1;width_per_section=8;section_size=8;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i70_512x8_sub_000000_000  (
    .addra({1'b0,\biu/l1i_addr ,3'b111}),
    .clka(clk_pad),
    .dia({open_n5976,\biu/l1i_in [63:56]}),
    .wea(\biu/cache/n31 ),
    .doa({open_n5991,ins_read[63:56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u0  (
    .a(\biu/cache_ctrl_logic/pa_temp [0]),
    .b(\biu/cache_ctrl_logic/off [0]),
    .c(\biu/cache_ctrl_logic/add0/c0 ),
    .o({\biu/cache_ctrl_logic/add0/c1 ,\biu/cache_ctrl_logic/n207 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u1  (
    .a(\biu/cache_ctrl_logic/pa_temp [1]),
    .b(\biu/cache_ctrl_logic/off [1]),
    .c(\biu/cache_ctrl_logic/add0/c1 ),
    .o({\biu/cache_ctrl_logic/add0/c2 ,\biu/cache_ctrl_logic/n207 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u10  (
    .a(\biu/cache_ctrl_logic/pa_temp [10]),
    .b(\biu/cache_ctrl_logic/off [10]),
    .c(\biu/cache_ctrl_logic/add0/c10 ),
    .o({\biu/cache_ctrl_logic/add0/c11 ,\biu/cache_ctrl_logic/n207 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u11  (
    .a(\biu/cache_ctrl_logic/pa_temp [11]),
    .b(\biu/cache_ctrl_logic/off [11]),
    .c(\biu/cache_ctrl_logic/add0/c11 ),
    .o({\biu/cache_ctrl_logic/add0/c12 ,\biu/cache_ctrl_logic/n207 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u12  (
    .a(\biu/cache_ctrl_logic/pa_temp [12]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c12 ),
    .o({\biu/cache_ctrl_logic/add0/c13 ,\biu/cache_ctrl_logic/n207 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u13  (
    .a(\biu/cache_ctrl_logic/pa_temp [13]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c13 ),
    .o({\biu/cache_ctrl_logic/add0/c14 ,\biu/cache_ctrl_logic/n207 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u14  (
    .a(\biu/cache_ctrl_logic/pa_temp [14]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c14 ),
    .o({\biu/cache_ctrl_logic/add0/c15 ,\biu/cache_ctrl_logic/n207 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u15  (
    .a(\biu/cache_ctrl_logic/pa_temp [15]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c15 ),
    .o({\biu/cache_ctrl_logic/add0/c16 ,\biu/cache_ctrl_logic/n207 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u16  (
    .a(\biu/cache_ctrl_logic/pa_temp [16]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c16 ),
    .o({\biu/cache_ctrl_logic/add0/c17 ,\biu/cache_ctrl_logic/n207 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u17  (
    .a(\biu/cache_ctrl_logic/pa_temp [17]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c17 ),
    .o({\biu/cache_ctrl_logic/add0/c18 ,\biu/cache_ctrl_logic/n207 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u18  (
    .a(\biu/cache_ctrl_logic/pa_temp [18]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c18 ),
    .o({\biu/cache_ctrl_logic/add0/c19 ,\biu/cache_ctrl_logic/n207 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u19  (
    .a(\biu/cache_ctrl_logic/pa_temp [19]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c19 ),
    .o({\biu/cache_ctrl_logic/add0/c20 ,\biu/cache_ctrl_logic/n207 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u2  (
    .a(\biu/cache_ctrl_logic/pa_temp [2]),
    .b(\biu/cache_ctrl_logic/off [2]),
    .c(\biu/cache_ctrl_logic/add0/c2 ),
    .o({\biu/cache_ctrl_logic/add0/c3 ,\biu/cache_ctrl_logic/n207 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u20  (
    .a(\biu/cache_ctrl_logic/pa_temp [20]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c20 ),
    .o({\biu/cache_ctrl_logic/add0/c21 ,\biu/cache_ctrl_logic/n207 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u21  (
    .a(\biu/cache_ctrl_logic/pa_temp [21]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c21 ),
    .o({\biu/cache_ctrl_logic/add0/c22 ,\biu/cache_ctrl_logic/n207 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u22  (
    .a(\biu/cache_ctrl_logic/pa_temp [22]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c22 ),
    .o({\biu/cache_ctrl_logic/add0/c23 ,\biu/cache_ctrl_logic/n207 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u23  (
    .a(\biu/cache_ctrl_logic/pa_temp [23]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c23 ),
    .o({\biu/cache_ctrl_logic/add0/c24 ,\biu/cache_ctrl_logic/n207 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u24  (
    .a(\biu/cache_ctrl_logic/pa_temp [24]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c24 ),
    .o({\biu/cache_ctrl_logic/add0/c25 ,\biu/cache_ctrl_logic/n207 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u25  (
    .a(\biu/cache_ctrl_logic/pa_temp [25]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c25 ),
    .o({\biu/cache_ctrl_logic/add0/c26 ,\biu/cache_ctrl_logic/n207 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u26  (
    .a(\biu/cache_ctrl_logic/pa_temp [26]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c26 ),
    .o({\biu/cache_ctrl_logic/add0/c27 ,\biu/cache_ctrl_logic/n207 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u27  (
    .a(\biu/cache_ctrl_logic/pa_temp [27]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c27 ),
    .o({\biu/cache_ctrl_logic/add0/c28 ,\biu/cache_ctrl_logic/n207 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u28  (
    .a(\biu/cache_ctrl_logic/pa_temp [28]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c28 ),
    .o({\biu/cache_ctrl_logic/add0/c29 ,\biu/cache_ctrl_logic/n207 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u29  (
    .a(\biu/cache_ctrl_logic/pa_temp [29]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c29 ),
    .o({\biu/cache_ctrl_logic/add0/c30 ,\biu/cache_ctrl_logic/n207 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u3  (
    .a(\biu/cache_ctrl_logic/pa_temp [3]),
    .b(\biu/cache_ctrl_logic/off [3]),
    .c(\biu/cache_ctrl_logic/add0/c3 ),
    .o({\biu/cache_ctrl_logic/add0/c4 ,\biu/cache_ctrl_logic/n207 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u30  (
    .a(\biu/cache_ctrl_logic/pa_temp [30]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c30 ),
    .o({\biu/cache_ctrl_logic/add0/c31 ,\biu/cache_ctrl_logic/n207 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u31  (
    .a(\biu/cache_ctrl_logic/pa_temp [31]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c31 ),
    .o({\biu/cache_ctrl_logic/add0/c32 ,\biu/cache_ctrl_logic/n207 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u32  (
    .a(\biu/cache_ctrl_logic/pa_temp [32]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c32 ),
    .o({\biu/cache_ctrl_logic/add0/c33 ,\biu/cache_ctrl_logic/n207 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u33  (
    .a(\biu/cache_ctrl_logic/pa_temp [33]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c33 ),
    .o({\biu/cache_ctrl_logic/add0/c34 ,\biu/cache_ctrl_logic/n207 [33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u34  (
    .a(\biu/cache_ctrl_logic/pa_temp [34]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c34 ),
    .o({\biu/cache_ctrl_logic/add0/c35 ,\biu/cache_ctrl_logic/n207 [34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u35  (
    .a(\biu/cache_ctrl_logic/pa_temp [35]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c35 ),
    .o({\biu/cache_ctrl_logic/add0/c36 ,\biu/cache_ctrl_logic/n207 [35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u36  (
    .a(\biu/cache_ctrl_logic/pa_temp [36]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c36 ),
    .o({\biu/cache_ctrl_logic/add0/c37 ,\biu/cache_ctrl_logic/n207 [36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u37  (
    .a(\biu/cache_ctrl_logic/pa_temp [37]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c37 ),
    .o({\biu/cache_ctrl_logic/add0/c38 ,\biu/cache_ctrl_logic/n207 [37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u38  (
    .a(\biu/cache_ctrl_logic/pa_temp [38]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c38 ),
    .o({\biu/cache_ctrl_logic/add0/c39 ,\biu/cache_ctrl_logic/n207 [38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u39  (
    .a(\biu/cache_ctrl_logic/pa_temp [39]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c39 ),
    .o({\biu/cache_ctrl_logic/add0/c40 ,\biu/cache_ctrl_logic/n207 [39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u4  (
    .a(\biu/cache_ctrl_logic/pa_temp [4]),
    .b(\biu/cache_ctrl_logic/off [4]),
    .c(\biu/cache_ctrl_logic/add0/c4 ),
    .o({\biu/cache_ctrl_logic/add0/c5 ,\biu/cache_ctrl_logic/n207 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u40  (
    .a(\biu/cache_ctrl_logic/pa_temp [40]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c40 ),
    .o({\biu/cache_ctrl_logic/add0/c41 ,\biu/cache_ctrl_logic/n207 [40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u41  (
    .a(\biu/cache_ctrl_logic/pa_temp [41]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c41 ),
    .o({\biu/cache_ctrl_logic/add0/c42 ,\biu/cache_ctrl_logic/n207 [41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u42  (
    .a(\biu/cache_ctrl_logic/pa_temp [42]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c42 ),
    .o({\biu/cache_ctrl_logic/add0/c43 ,\biu/cache_ctrl_logic/n207 [42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u43  (
    .a(\biu/cache_ctrl_logic/pa_temp [43]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c43 ),
    .o({\biu/cache_ctrl_logic/add0/c44 ,\biu/cache_ctrl_logic/n207 [43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u44  (
    .a(\biu/cache_ctrl_logic/pa_temp [44]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c44 ),
    .o({\biu/cache_ctrl_logic/add0/c45 ,\biu/cache_ctrl_logic/n207 [44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u45  (
    .a(\biu/cache_ctrl_logic/pa_temp [45]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c45 ),
    .o({\biu/cache_ctrl_logic/add0/c46 ,\biu/cache_ctrl_logic/n207 [45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u46  (
    .a(\biu/cache_ctrl_logic/pa_temp [46]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c46 ),
    .o({\biu/cache_ctrl_logic/add0/c47 ,\biu/cache_ctrl_logic/n207 [46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u47  (
    .a(\biu/cache_ctrl_logic/pa_temp [47]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c47 ),
    .o({\biu/cache_ctrl_logic/add0/c48 ,\biu/cache_ctrl_logic/n207 [47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u48  (
    .a(\biu/cache_ctrl_logic/pa_temp [48]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c48 ),
    .o({\biu/cache_ctrl_logic/add0/c49 ,\biu/cache_ctrl_logic/n207 [48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u49  (
    .a(\biu/cache_ctrl_logic/pa_temp [49]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c49 ),
    .o({\biu/cache_ctrl_logic/add0/c50 ,\biu/cache_ctrl_logic/n207 [49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u5  (
    .a(\biu/cache_ctrl_logic/pa_temp [5]),
    .b(\biu/cache_ctrl_logic/off [5]),
    .c(\biu/cache_ctrl_logic/add0/c5 ),
    .o({\biu/cache_ctrl_logic/add0/c6 ,\biu/cache_ctrl_logic/n207 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u50  (
    .a(\biu/cache_ctrl_logic/pa_temp [50]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c50 ),
    .o({\biu/cache_ctrl_logic/add0/c51 ,\biu/cache_ctrl_logic/n207 [50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u51  (
    .a(\biu/cache_ctrl_logic/pa_temp [51]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c51 ),
    .o({\biu/cache_ctrl_logic/add0/c52 ,\biu/cache_ctrl_logic/n207 [51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u52  (
    .a(\biu/cache_ctrl_logic/pa_temp [52]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c52 ),
    .o({\biu/cache_ctrl_logic/add0/c53 ,\biu/cache_ctrl_logic/n207 [52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u53  (
    .a(\biu/cache_ctrl_logic/pa_temp [53]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c53 ),
    .o({\biu/cache_ctrl_logic/add0/c54 ,\biu/cache_ctrl_logic/n207 [53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u54  (
    .a(\biu/cache_ctrl_logic/pa_temp [54]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c54 ),
    .o({\biu/cache_ctrl_logic/add0/c55 ,\biu/cache_ctrl_logic/n207 [54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u55  (
    .a(\biu/cache_ctrl_logic/pa_temp [55]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c55 ),
    .o({\biu/cache_ctrl_logic/add0/c56 ,\biu/cache_ctrl_logic/n207 [55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u56  (
    .a(\biu/cache_ctrl_logic/pa_temp [56]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c56 ),
    .o({\biu/cache_ctrl_logic/add0/c57 ,\biu/cache_ctrl_logic/n207 [56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u57  (
    .a(\biu/cache_ctrl_logic/pa_temp [57]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c57 ),
    .o({\biu/cache_ctrl_logic/add0/c58 ,\biu/cache_ctrl_logic/n207 [57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u58  (
    .a(\biu/cache_ctrl_logic/pa_temp [58]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c58 ),
    .o({\biu/cache_ctrl_logic/add0/c59 ,\biu/cache_ctrl_logic/n207 [58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u59  (
    .a(\biu/cache_ctrl_logic/pa_temp [59]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c59 ),
    .o({\biu/cache_ctrl_logic/add0/c60 ,\biu/cache_ctrl_logic/n207 [59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u6  (
    .a(\biu/cache_ctrl_logic/pa_temp [6]),
    .b(\biu/cache_ctrl_logic/off [6]),
    .c(\biu/cache_ctrl_logic/add0/c6 ),
    .o({\biu/cache_ctrl_logic/add0/c7 ,\biu/cache_ctrl_logic/n207 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u60  (
    .a(\biu/cache_ctrl_logic/pa_temp [60]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c60 ),
    .o({\biu/cache_ctrl_logic/add0/c61 ,\biu/cache_ctrl_logic/n207 [60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u61  (
    .a(\biu/cache_ctrl_logic/pa_temp [61]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c61 ),
    .o({\biu/cache_ctrl_logic/add0/c62 ,\biu/cache_ctrl_logic/n207 [61]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u62  (
    .a(\biu/cache_ctrl_logic/pa_temp [62]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c62 ),
    .o({\biu/cache_ctrl_logic/add0/c63 ,\biu/cache_ctrl_logic/n207 [62]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u63  (
    .a(\biu/cache_ctrl_logic/pa_temp [63]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add0/c63 ),
    .o({open_n6001,\biu/cache_ctrl_logic/n207 [63]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u7  (
    .a(\biu/cache_ctrl_logic/pa_temp [7]),
    .b(\biu/cache_ctrl_logic/off [7]),
    .c(\biu/cache_ctrl_logic/add0/c7 ),
    .o({\biu/cache_ctrl_logic/add0/c8 ,\biu/cache_ctrl_logic/n207 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u8  (
    .a(\biu/cache_ctrl_logic/pa_temp [8]),
    .b(\biu/cache_ctrl_logic/off [8]),
    .c(\biu/cache_ctrl_logic/add0/c8 ),
    .o({\biu/cache_ctrl_logic/add0/c9 ,\biu/cache_ctrl_logic/n207 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add0/u9  (
    .a(\biu/cache_ctrl_logic/pa_temp [9]),
    .b(\biu/cache_ctrl_logic/off [9]),
    .c(\biu/cache_ctrl_logic/add0/c9 ),
    .o({\biu/cache_ctrl_logic/add0/c10 ,\biu/cache_ctrl_logic/n207 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \biu/cache_ctrl_logic/add0/ucin  (
    .a(1'b0),
    .o({\biu/cache_ctrl_logic/add0/c0 ,open_n6004}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u0  (
    .a(\biu/cache_ctrl_logic/l1i_pa [0]),
    .b(\biu/cache_ctrl_logic/off [0]),
    .c(\biu/cache_ctrl_logic/add1/c0 ),
    .o({\biu/cache_ctrl_logic/add1/c1 ,\biu/cache_ctrl_logic/n209 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u1  (
    .a(\biu/cache_ctrl_logic/l1i_pa [1]),
    .b(\biu/cache_ctrl_logic/off [1]),
    .c(\biu/cache_ctrl_logic/add1/c1 ),
    .o({\biu/cache_ctrl_logic/add1/c2 ,\biu/cache_ctrl_logic/n209 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u10  (
    .a(\biu/cache_ctrl_logic/l1i_pa [10]),
    .b(\biu/cache_ctrl_logic/off [10]),
    .c(\biu/cache_ctrl_logic/add1/c10 ),
    .o({\biu/cache_ctrl_logic/add1/c11 ,\biu/cache_ctrl_logic/n209 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u11  (
    .a(\biu/cache_ctrl_logic/l1i_pa [11]),
    .b(\biu/cache_ctrl_logic/off [11]),
    .c(\biu/cache_ctrl_logic/add1/c11 ),
    .o({\biu/cache_ctrl_logic/add1/c12 ,\biu/cache_ctrl_logic/n209 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u12  (
    .a(\biu/cache_ctrl_logic/l1i_pa [12]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c12 ),
    .o({\biu/cache_ctrl_logic/add1/c13 ,\biu/cache_ctrl_logic/n209 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u13  (
    .a(\biu/cache_ctrl_logic/l1i_pa [13]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c13 ),
    .o({\biu/cache_ctrl_logic/add1/c14 ,\biu/cache_ctrl_logic/n209 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u14  (
    .a(\biu/cache_ctrl_logic/l1i_pa [14]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c14 ),
    .o({\biu/cache_ctrl_logic/add1/c15 ,\biu/cache_ctrl_logic/n209 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u15  (
    .a(\biu/cache_ctrl_logic/l1i_pa [15]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c15 ),
    .o({\biu/cache_ctrl_logic/add1/c16 ,\biu/cache_ctrl_logic/n209 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u16  (
    .a(\biu/cache_ctrl_logic/l1i_pa [16]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c16 ),
    .o({\biu/cache_ctrl_logic/add1/c17 ,\biu/cache_ctrl_logic/n209 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u17  (
    .a(\biu/cache_ctrl_logic/l1i_pa [17]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c17 ),
    .o({\biu/cache_ctrl_logic/add1/c18 ,\biu/cache_ctrl_logic/n209 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u18  (
    .a(\biu/cache_ctrl_logic/l1i_pa [18]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c18 ),
    .o({\biu/cache_ctrl_logic/add1/c19 ,\biu/cache_ctrl_logic/n209 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u19  (
    .a(\biu/cache_ctrl_logic/l1i_pa [19]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c19 ),
    .o({\biu/cache_ctrl_logic/add1/c20 ,\biu/cache_ctrl_logic/n209 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u2  (
    .a(\biu/cache_ctrl_logic/l1i_pa [2]),
    .b(\biu/cache_ctrl_logic/off [2]),
    .c(\biu/cache_ctrl_logic/add1/c2 ),
    .o({\biu/cache_ctrl_logic/add1/c3 ,\biu/cache_ctrl_logic/n209 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u20  (
    .a(\biu/cache_ctrl_logic/l1i_pa [20]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c20 ),
    .o({\biu/cache_ctrl_logic/add1/c21 ,\biu/cache_ctrl_logic/n209 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u21  (
    .a(\biu/cache_ctrl_logic/l1i_pa [21]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c21 ),
    .o({\biu/cache_ctrl_logic/add1/c22 ,\biu/cache_ctrl_logic/n209 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u22  (
    .a(\biu/cache_ctrl_logic/l1i_pa [22]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c22 ),
    .o({\biu/cache_ctrl_logic/add1/c23 ,\biu/cache_ctrl_logic/n209 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u23  (
    .a(\biu/cache_ctrl_logic/l1i_pa [23]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c23 ),
    .o({\biu/cache_ctrl_logic/add1/c24 ,\biu/cache_ctrl_logic/n209 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u24  (
    .a(\biu/cache_ctrl_logic/l1i_pa [24]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c24 ),
    .o({\biu/cache_ctrl_logic/add1/c25 ,\biu/cache_ctrl_logic/n209 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u25  (
    .a(\biu/cache_ctrl_logic/l1i_pa [25]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c25 ),
    .o({\biu/cache_ctrl_logic/add1/c26 ,\biu/cache_ctrl_logic/n209 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u26  (
    .a(\biu/cache_ctrl_logic/l1i_pa [26]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c26 ),
    .o({\biu/cache_ctrl_logic/add1/c27 ,\biu/cache_ctrl_logic/n209 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u27  (
    .a(\biu/cache_ctrl_logic/l1i_pa [27]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c27 ),
    .o({\biu/cache_ctrl_logic/add1/c28 ,\biu/cache_ctrl_logic/n209 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u28  (
    .a(\biu/cache_ctrl_logic/l1i_pa [28]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c28 ),
    .o({\biu/cache_ctrl_logic/add1/c29 ,\biu/cache_ctrl_logic/n209 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u29  (
    .a(\biu/cache_ctrl_logic/l1i_pa [29]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c29 ),
    .o({\biu/cache_ctrl_logic/add1/c30 ,\biu/cache_ctrl_logic/n209 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u3  (
    .a(\biu/cache_ctrl_logic/l1i_pa [3]),
    .b(\biu/cache_ctrl_logic/off [3]),
    .c(\biu/cache_ctrl_logic/add1/c3 ),
    .o({\biu/cache_ctrl_logic/add1/c4 ,\biu/cache_ctrl_logic/n209 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u30  (
    .a(\biu/cache_ctrl_logic/l1i_pa [30]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c30 ),
    .o({\biu/cache_ctrl_logic/add1/c31 ,\biu/cache_ctrl_logic/n209 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u31  (
    .a(\biu/cache_ctrl_logic/l1i_pa [31]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c31 ),
    .o({\biu/cache_ctrl_logic/add1/c32 ,\biu/cache_ctrl_logic/n209 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u32  (
    .a(\biu/cache_ctrl_logic/l1i_pa [32]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c32 ),
    .o({\biu/cache_ctrl_logic/add1/c33 ,\biu/cache_ctrl_logic/n209 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u33  (
    .a(\biu/cache_ctrl_logic/l1i_pa [33]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c33 ),
    .o({\biu/cache_ctrl_logic/add1/c34 ,\biu/cache_ctrl_logic/n209 [33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u34  (
    .a(\biu/cache_ctrl_logic/l1i_pa [34]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c34 ),
    .o({\biu/cache_ctrl_logic/add1/c35 ,\biu/cache_ctrl_logic/n209 [34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u35  (
    .a(\biu/cache_ctrl_logic/l1i_pa [35]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c35 ),
    .o({\biu/cache_ctrl_logic/add1/c36 ,\biu/cache_ctrl_logic/n209 [35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u36  (
    .a(\biu/cache_ctrl_logic/l1i_pa [36]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c36 ),
    .o({\biu/cache_ctrl_logic/add1/c37 ,\biu/cache_ctrl_logic/n209 [36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u37  (
    .a(\biu/cache_ctrl_logic/l1i_pa [37]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c37 ),
    .o({\biu/cache_ctrl_logic/add1/c38 ,\biu/cache_ctrl_logic/n209 [37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u38  (
    .a(\biu/cache_ctrl_logic/l1i_pa [38]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c38 ),
    .o({\biu/cache_ctrl_logic/add1/c39 ,\biu/cache_ctrl_logic/n209 [38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u39  (
    .a(\biu/cache_ctrl_logic/l1i_pa [39]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c39 ),
    .o({\biu/cache_ctrl_logic/add1/c40 ,\biu/cache_ctrl_logic/n209 [39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u4  (
    .a(\biu/cache_ctrl_logic/l1i_pa [4]),
    .b(\biu/cache_ctrl_logic/off [4]),
    .c(\biu/cache_ctrl_logic/add1/c4 ),
    .o({\biu/cache_ctrl_logic/add1/c5 ,\biu/cache_ctrl_logic/n209 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u40  (
    .a(\biu/cache_ctrl_logic/l1i_pa [40]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c40 ),
    .o({\biu/cache_ctrl_logic/add1/c41 ,\biu/cache_ctrl_logic/n209 [40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u41  (
    .a(\biu/cache_ctrl_logic/l1i_pa [41]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c41 ),
    .o({\biu/cache_ctrl_logic/add1/c42 ,\biu/cache_ctrl_logic/n209 [41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u42  (
    .a(\biu/cache_ctrl_logic/l1i_pa [42]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c42 ),
    .o({\biu/cache_ctrl_logic/add1/c43 ,\biu/cache_ctrl_logic/n209 [42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u43  (
    .a(\biu/cache_ctrl_logic/l1i_pa [43]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c43 ),
    .o({\biu/cache_ctrl_logic/add1/c44 ,\biu/cache_ctrl_logic/n209 [43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u44  (
    .a(\biu/cache_ctrl_logic/l1i_pa [44]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c44 ),
    .o({\biu/cache_ctrl_logic/add1/c45 ,\biu/cache_ctrl_logic/n209 [44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u45  (
    .a(\biu/cache_ctrl_logic/l1i_pa [45]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c45 ),
    .o({\biu/cache_ctrl_logic/add1/c46 ,\biu/cache_ctrl_logic/n209 [45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u46  (
    .a(\biu/cache_ctrl_logic/l1i_pa [46]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c46 ),
    .o({\biu/cache_ctrl_logic/add1/c47 ,\biu/cache_ctrl_logic/n209 [46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u47  (
    .a(\biu/cache_ctrl_logic/l1i_pa [47]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c47 ),
    .o({\biu/cache_ctrl_logic/add1/c48 ,\biu/cache_ctrl_logic/n209 [47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u48  (
    .a(\biu/cache_ctrl_logic/l1i_pa [48]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c48 ),
    .o({\biu/cache_ctrl_logic/add1/c49 ,\biu/cache_ctrl_logic/n209 [48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u49  (
    .a(\biu/cache_ctrl_logic/l1i_pa [49]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c49 ),
    .o({\biu/cache_ctrl_logic/add1/c50 ,\biu/cache_ctrl_logic/n209 [49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u5  (
    .a(\biu/cache_ctrl_logic/l1i_pa [5]),
    .b(\biu/cache_ctrl_logic/off [5]),
    .c(\biu/cache_ctrl_logic/add1/c5 ),
    .o({\biu/cache_ctrl_logic/add1/c6 ,\biu/cache_ctrl_logic/n209 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u50  (
    .a(\biu/cache_ctrl_logic/l1i_pa [50]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c50 ),
    .o({\biu/cache_ctrl_logic/add1/c51 ,\biu/cache_ctrl_logic/n209 [50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u51  (
    .a(\biu/cache_ctrl_logic/l1i_pa [51]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c51 ),
    .o({\biu/cache_ctrl_logic/add1/c52 ,\biu/cache_ctrl_logic/n209 [51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u52  (
    .a(\biu/cache_ctrl_logic/l1i_pa [52]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c52 ),
    .o({\biu/cache_ctrl_logic/add1/c53 ,\biu/cache_ctrl_logic/n209 [52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u53  (
    .a(\biu/cache_ctrl_logic/l1i_pa [53]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c53 ),
    .o({\biu/cache_ctrl_logic/add1/c54 ,\biu/cache_ctrl_logic/n209 [53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u54  (
    .a(\biu/cache_ctrl_logic/l1i_pa [54]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c54 ),
    .o({\biu/cache_ctrl_logic/add1/c55 ,\biu/cache_ctrl_logic/n209 [54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u55  (
    .a(\biu/cache_ctrl_logic/l1i_pa [55]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c55 ),
    .o({\biu/cache_ctrl_logic/add1/c56 ,\biu/cache_ctrl_logic/n209 [55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u56  (
    .a(\biu/cache_ctrl_logic/l1i_pa [56]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c56 ),
    .o({\biu/cache_ctrl_logic/add1/c57 ,\biu/cache_ctrl_logic/n209 [56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u57  (
    .a(\biu/cache_ctrl_logic/l1i_pa [57]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c57 ),
    .o({\biu/cache_ctrl_logic/add1/c58 ,\biu/cache_ctrl_logic/n209 [57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u58  (
    .a(\biu/cache_ctrl_logic/l1i_pa [58]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c58 ),
    .o({\biu/cache_ctrl_logic/add1/c59 ,\biu/cache_ctrl_logic/n209 [58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u59  (
    .a(\biu/cache_ctrl_logic/l1i_pa [59]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c59 ),
    .o({\biu/cache_ctrl_logic/add1/c60 ,\biu/cache_ctrl_logic/n209 [59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u6  (
    .a(\biu/cache_ctrl_logic/l1i_pa [6]),
    .b(\biu/cache_ctrl_logic/off [6]),
    .c(\biu/cache_ctrl_logic/add1/c6 ),
    .o({\biu/cache_ctrl_logic/add1/c7 ,\biu/cache_ctrl_logic/n209 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u60  (
    .a(\biu/cache_ctrl_logic/l1i_pa [60]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c60 ),
    .o({\biu/cache_ctrl_logic/add1/c61 ,\biu/cache_ctrl_logic/n209 [60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u61  (
    .a(\biu/cache_ctrl_logic/l1i_pa [61]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c61 ),
    .o({\biu/cache_ctrl_logic/add1/c62 ,\biu/cache_ctrl_logic/n209 [61]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u62  (
    .a(\biu/cache_ctrl_logic/l1i_pa [62]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c62 ),
    .o({\biu/cache_ctrl_logic/add1/c63 ,\biu/cache_ctrl_logic/n209 [62]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u63  (
    .a(\biu/cache_ctrl_logic/l1i_pa [63]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add1/c63 ),
    .o({open_n6005,\biu/cache_ctrl_logic/n209 [63]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u7  (
    .a(\biu/cache_ctrl_logic/l1i_pa [7]),
    .b(\biu/cache_ctrl_logic/off [7]),
    .c(\biu/cache_ctrl_logic/add1/c7 ),
    .o({\biu/cache_ctrl_logic/add1/c8 ,\biu/cache_ctrl_logic/n209 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u8  (
    .a(\biu/cache_ctrl_logic/l1i_pa [8]),
    .b(\biu/cache_ctrl_logic/off [8]),
    .c(\biu/cache_ctrl_logic/add1/c8 ),
    .o({\biu/cache_ctrl_logic/add1/c9 ,\biu/cache_ctrl_logic/n209 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add1/u9  (
    .a(\biu/cache_ctrl_logic/l1i_pa [9]),
    .b(\biu/cache_ctrl_logic/off [9]),
    .c(\biu/cache_ctrl_logic/add1/c9 ),
    .o({\biu/cache_ctrl_logic/add1/c10 ,\biu/cache_ctrl_logic/n209 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \biu/cache_ctrl_logic/add1/ucin  (
    .a(1'b0),
    .o({\biu/cache_ctrl_logic/add1/c0 ,open_n6008}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u0  (
    .a(\biu/cache_ctrl_logic/l1d_pa [0]),
    .b(\biu/cache_ctrl_logic/off [0]),
    .c(\biu/cache_ctrl_logic/add2/c0 ),
    .o({\biu/cache_ctrl_logic/add2/c1 ,\biu/cache_ctrl_logic/n212 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u1  (
    .a(\biu/cache_ctrl_logic/l1d_pa [1]),
    .b(\biu/cache_ctrl_logic/off [1]),
    .c(\biu/cache_ctrl_logic/add2/c1 ),
    .o({\biu/cache_ctrl_logic/add2/c2 ,\biu/cache_ctrl_logic/n212 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u10  (
    .a(\biu/cache_ctrl_logic/l1d_pa [10]),
    .b(\biu/cache_ctrl_logic/off [10]),
    .c(\biu/cache_ctrl_logic/add2/c10 ),
    .o({\biu/cache_ctrl_logic/add2/c11 ,\biu/cache_ctrl_logic/n212 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u11  (
    .a(\biu/cache_ctrl_logic/l1d_pa [11]),
    .b(\biu/cache_ctrl_logic/off [11]),
    .c(\biu/cache_ctrl_logic/add2/c11 ),
    .o({\biu/cache_ctrl_logic/add2/c12 ,\biu/cache_ctrl_logic/n212 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u12  (
    .a(\biu/cache_ctrl_logic/l1d_pa [12]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c12 ),
    .o({\biu/cache_ctrl_logic/add2/c13 ,\biu/cache_ctrl_logic/n212 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u13  (
    .a(\biu/cache_ctrl_logic/l1d_pa [13]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c13 ),
    .o({\biu/cache_ctrl_logic/add2/c14 ,\biu/cache_ctrl_logic/n212 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u14  (
    .a(\biu/cache_ctrl_logic/l1d_pa [14]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c14 ),
    .o({\biu/cache_ctrl_logic/add2/c15 ,\biu/cache_ctrl_logic/n212 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u15  (
    .a(\biu/cache_ctrl_logic/l1d_pa [15]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c15 ),
    .o({\biu/cache_ctrl_logic/add2/c16 ,\biu/cache_ctrl_logic/n212 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u16  (
    .a(\biu/cache_ctrl_logic/l1d_pa [16]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c16 ),
    .o({\biu/cache_ctrl_logic/add2/c17 ,\biu/cache_ctrl_logic/n212 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u17  (
    .a(\biu/cache_ctrl_logic/l1d_pa [17]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c17 ),
    .o({\biu/cache_ctrl_logic/add2/c18 ,\biu/cache_ctrl_logic/n212 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u18  (
    .a(\biu/cache_ctrl_logic/l1d_pa [18]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c18 ),
    .o({\biu/cache_ctrl_logic/add2/c19 ,\biu/cache_ctrl_logic/n212 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u19  (
    .a(\biu/cache_ctrl_logic/l1d_pa [19]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c19 ),
    .o({\biu/cache_ctrl_logic/add2/c20 ,\biu/cache_ctrl_logic/n212 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u2  (
    .a(\biu/cache_ctrl_logic/l1d_pa [2]),
    .b(\biu/cache_ctrl_logic/off [2]),
    .c(\biu/cache_ctrl_logic/add2/c2 ),
    .o({\biu/cache_ctrl_logic/add2/c3 ,\biu/cache_ctrl_logic/n212 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u20  (
    .a(\biu/cache_ctrl_logic/l1d_pa [20]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c20 ),
    .o({\biu/cache_ctrl_logic/add2/c21 ,\biu/cache_ctrl_logic/n212 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u21  (
    .a(\biu/cache_ctrl_logic/l1d_pa [21]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c21 ),
    .o({\biu/cache_ctrl_logic/add2/c22 ,\biu/cache_ctrl_logic/n212 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u22  (
    .a(\biu/cache_ctrl_logic/l1d_pa [22]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c22 ),
    .o({\biu/cache_ctrl_logic/add2/c23 ,\biu/cache_ctrl_logic/n212 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u23  (
    .a(\biu/cache_ctrl_logic/l1d_pa [23]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c23 ),
    .o({\biu/cache_ctrl_logic/add2/c24 ,\biu/cache_ctrl_logic/n212 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u24  (
    .a(\biu/cache_ctrl_logic/l1d_pa [24]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c24 ),
    .o({\biu/cache_ctrl_logic/add2/c25 ,\biu/cache_ctrl_logic/n212 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u25  (
    .a(\biu/cache_ctrl_logic/l1d_pa [25]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c25 ),
    .o({\biu/cache_ctrl_logic/add2/c26 ,\biu/cache_ctrl_logic/n212 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u26  (
    .a(\biu/cache_ctrl_logic/l1d_pa [26]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c26 ),
    .o({\biu/cache_ctrl_logic/add2/c27 ,\biu/cache_ctrl_logic/n212 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u27  (
    .a(\biu/cache_ctrl_logic/l1d_pa [27]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c27 ),
    .o({\biu/cache_ctrl_logic/add2/c28 ,\biu/cache_ctrl_logic/n212 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u28  (
    .a(\biu/cache_ctrl_logic/l1d_pa [28]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c28 ),
    .o({\biu/cache_ctrl_logic/add2/c29 ,\biu/cache_ctrl_logic/n212 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u29  (
    .a(\biu/cache_ctrl_logic/l1d_pa [29]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c29 ),
    .o({\biu/cache_ctrl_logic/add2/c30 ,\biu/cache_ctrl_logic/n212 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u3  (
    .a(\biu/cache_ctrl_logic/l1d_pa [3]),
    .b(\biu/cache_ctrl_logic/off [3]),
    .c(\biu/cache_ctrl_logic/add2/c3 ),
    .o({\biu/cache_ctrl_logic/add2/c4 ,\biu/cache_ctrl_logic/n212 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u30  (
    .a(\biu/cache_ctrl_logic/l1d_pa [30]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c30 ),
    .o({\biu/cache_ctrl_logic/add2/c31 ,\biu/cache_ctrl_logic/n212 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u31  (
    .a(\biu/cache_ctrl_logic/l1d_pa [31]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c31 ),
    .o({\biu/cache_ctrl_logic/add2/c32 ,\biu/cache_ctrl_logic/n212 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u32  (
    .a(\biu/cache_ctrl_logic/l1d_pa [32]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c32 ),
    .o({\biu/cache_ctrl_logic/add2/c33 ,\biu/cache_ctrl_logic/n212 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u33  (
    .a(\biu/cache_ctrl_logic/l1d_pa [33]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c33 ),
    .o({\biu/cache_ctrl_logic/add2/c34 ,\biu/cache_ctrl_logic/n212 [33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u34  (
    .a(\biu/cache_ctrl_logic/l1d_pa [34]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c34 ),
    .o({\biu/cache_ctrl_logic/add2/c35 ,\biu/cache_ctrl_logic/n212 [34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u35  (
    .a(\biu/cache_ctrl_logic/l1d_pa [35]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c35 ),
    .o({\biu/cache_ctrl_logic/add2/c36 ,\biu/cache_ctrl_logic/n212 [35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u36  (
    .a(\biu/cache_ctrl_logic/l1d_pa [36]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c36 ),
    .o({\biu/cache_ctrl_logic/add2/c37 ,\biu/cache_ctrl_logic/n212 [36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u37  (
    .a(\biu/cache_ctrl_logic/l1d_pa [37]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c37 ),
    .o({\biu/cache_ctrl_logic/add2/c38 ,\biu/cache_ctrl_logic/n212 [37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u38  (
    .a(\biu/cache_ctrl_logic/l1d_pa [38]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c38 ),
    .o({\biu/cache_ctrl_logic/add2/c39 ,\biu/cache_ctrl_logic/n212 [38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u39  (
    .a(\biu/cache_ctrl_logic/l1d_pa [39]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c39 ),
    .o({\biu/cache_ctrl_logic/add2/c40 ,\biu/cache_ctrl_logic/n212 [39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u4  (
    .a(\biu/cache_ctrl_logic/l1d_pa [4]),
    .b(\biu/cache_ctrl_logic/off [4]),
    .c(\biu/cache_ctrl_logic/add2/c4 ),
    .o({\biu/cache_ctrl_logic/add2/c5 ,\biu/cache_ctrl_logic/n212 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u40  (
    .a(\biu/cache_ctrl_logic/l1d_pa [40]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c40 ),
    .o({\biu/cache_ctrl_logic/add2/c41 ,\biu/cache_ctrl_logic/n212 [40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u41  (
    .a(\biu/cache_ctrl_logic/l1d_pa [41]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c41 ),
    .o({\biu/cache_ctrl_logic/add2/c42 ,\biu/cache_ctrl_logic/n212 [41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u42  (
    .a(\biu/cache_ctrl_logic/l1d_pa [42]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c42 ),
    .o({\biu/cache_ctrl_logic/add2/c43 ,\biu/cache_ctrl_logic/n212 [42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u43  (
    .a(\biu/cache_ctrl_logic/l1d_pa [43]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c43 ),
    .o({\biu/cache_ctrl_logic/add2/c44 ,\biu/cache_ctrl_logic/n212 [43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u44  (
    .a(\biu/cache_ctrl_logic/l1d_pa [44]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c44 ),
    .o({\biu/cache_ctrl_logic/add2/c45 ,\biu/cache_ctrl_logic/n212 [44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u45  (
    .a(\biu/cache_ctrl_logic/l1d_pa [45]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c45 ),
    .o({\biu/cache_ctrl_logic/add2/c46 ,\biu/cache_ctrl_logic/n212 [45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u46  (
    .a(\biu/cache_ctrl_logic/l1d_pa [46]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c46 ),
    .o({\biu/cache_ctrl_logic/add2/c47 ,\biu/cache_ctrl_logic/n212 [46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u47  (
    .a(\biu/cache_ctrl_logic/l1d_pa [47]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c47 ),
    .o({\biu/cache_ctrl_logic/add2/c48 ,\biu/cache_ctrl_logic/n212 [47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u48  (
    .a(\biu/cache_ctrl_logic/l1d_pa [48]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c48 ),
    .o({\biu/cache_ctrl_logic/add2/c49 ,\biu/cache_ctrl_logic/n212 [48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u49  (
    .a(\biu/cache_ctrl_logic/l1d_pa [49]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c49 ),
    .o({\biu/cache_ctrl_logic/add2/c50 ,\biu/cache_ctrl_logic/n212 [49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u5  (
    .a(\biu/cache_ctrl_logic/l1d_pa [5]),
    .b(\biu/cache_ctrl_logic/off [5]),
    .c(\biu/cache_ctrl_logic/add2/c5 ),
    .o({\biu/cache_ctrl_logic/add2/c6 ,\biu/cache_ctrl_logic/n212 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u50  (
    .a(\biu/cache_ctrl_logic/l1d_pa [50]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c50 ),
    .o({\biu/cache_ctrl_logic/add2/c51 ,\biu/cache_ctrl_logic/n212 [50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u51  (
    .a(\biu/cache_ctrl_logic/l1d_pa [51]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c51 ),
    .o({\biu/cache_ctrl_logic/add2/c52 ,\biu/cache_ctrl_logic/n212 [51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u52  (
    .a(\biu/cache_ctrl_logic/l1d_pa [52]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c52 ),
    .o({\biu/cache_ctrl_logic/add2/c53 ,\biu/cache_ctrl_logic/n212 [52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u53  (
    .a(\biu/cache_ctrl_logic/l1d_pa [53]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c53 ),
    .o({\biu/cache_ctrl_logic/add2/c54 ,\biu/cache_ctrl_logic/n212 [53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u54  (
    .a(\biu/cache_ctrl_logic/l1d_pa [54]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c54 ),
    .o({\biu/cache_ctrl_logic/add2/c55 ,\biu/cache_ctrl_logic/n212 [54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u55  (
    .a(\biu/cache_ctrl_logic/l1d_pa [55]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c55 ),
    .o({\biu/cache_ctrl_logic/add2/c56 ,\biu/cache_ctrl_logic/n212 [55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u56  (
    .a(\biu/cache_ctrl_logic/l1d_pa [56]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c56 ),
    .o({\biu/cache_ctrl_logic/add2/c57 ,\biu/cache_ctrl_logic/n212 [56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u57  (
    .a(\biu/cache_ctrl_logic/l1d_pa [57]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c57 ),
    .o({\biu/cache_ctrl_logic/add2/c58 ,\biu/cache_ctrl_logic/n212 [57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u58  (
    .a(\biu/cache_ctrl_logic/l1d_pa [58]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c58 ),
    .o({\biu/cache_ctrl_logic/add2/c59 ,\biu/cache_ctrl_logic/n212 [58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u59  (
    .a(\biu/cache_ctrl_logic/l1d_pa [59]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c59 ),
    .o({\biu/cache_ctrl_logic/add2/c60 ,\biu/cache_ctrl_logic/n212 [59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u6  (
    .a(\biu/cache_ctrl_logic/l1d_pa [6]),
    .b(\biu/cache_ctrl_logic/off [6]),
    .c(\biu/cache_ctrl_logic/add2/c6 ),
    .o({\biu/cache_ctrl_logic/add2/c7 ,\biu/cache_ctrl_logic/n212 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u60  (
    .a(\biu/cache_ctrl_logic/l1d_pa [60]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c60 ),
    .o({\biu/cache_ctrl_logic/add2/c61 ,\biu/cache_ctrl_logic/n212 [60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u61  (
    .a(\biu/cache_ctrl_logic/l1d_pa [61]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c61 ),
    .o({\biu/cache_ctrl_logic/add2/c62 ,\biu/cache_ctrl_logic/n212 [61]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u62  (
    .a(\biu/cache_ctrl_logic/l1d_pa [62]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c62 ),
    .o({\biu/cache_ctrl_logic/add2/c63 ,\biu/cache_ctrl_logic/n212 [62]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u63  (
    .a(\biu/cache_ctrl_logic/l1d_pa [63]),
    .b(1'b0),
    .c(\biu/cache_ctrl_logic/add2/c63 ),
    .o({open_n6009,\biu/cache_ctrl_logic/n212 [63]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u7  (
    .a(\biu/cache_ctrl_logic/l1d_pa [7]),
    .b(\biu/cache_ctrl_logic/off [7]),
    .c(\biu/cache_ctrl_logic/add2/c7 ),
    .o({\biu/cache_ctrl_logic/add2/c8 ,\biu/cache_ctrl_logic/n212 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u8  (
    .a(\biu/cache_ctrl_logic/l1d_pa [8]),
    .b(\biu/cache_ctrl_logic/off [8]),
    .c(\biu/cache_ctrl_logic/add2/c8 ),
    .o({\biu/cache_ctrl_logic/add2/c9 ,\biu/cache_ctrl_logic/n212 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \biu/cache_ctrl_logic/add2/u9  (
    .a(\biu/cache_ctrl_logic/l1d_pa [9]),
    .b(\biu/cache_ctrl_logic/off [9]),
    .c(\biu/cache_ctrl_logic/add2/c9 ),
    .o({\biu/cache_ctrl_logic/add2/c10 ,\biu/cache_ctrl_logic/n212 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \biu/cache_ctrl_logic/add2/ucin  (
    .a(1'b0),
    .o({\biu/cache_ctrl_logic/add2/c0 ,open_n6012}));
  reg_sr_as_w1 \biu/cache_ctrl_logic/l1d_value_reg  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/l1d_value_d ),
    .en(1'b1),
    .reset(~\biu/cache_ctrl_logic/u128_sel_is_0_o ),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_value ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(394)
  reg_sr_as_w1 \biu/cache_ctrl_logic/l1i_value_reg  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/l1i_value_d ),
    .en(1'b1),
    .reset(~\biu/cache_ctrl_logic/u128_sel_is_0_o ),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_value ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(347)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b12  (
    .clk(clk_pad),
    .d(addr_if[12]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b13  (
    .clk(clk_pad),
    .d(addr_if[13]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b14  (
    .clk(clk_pad),
    .d(addr_if[14]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b15  (
    .clk(clk_pad),
    .d(addr_if[15]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b16  (
    .clk(clk_pad),
    .d(addr_if[16]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b17  (
    .clk(clk_pad),
    .d(addr_if[17]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b18  (
    .clk(clk_pad),
    .d(addr_if[18]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b19  (
    .clk(clk_pad),
    .d(addr_if[19]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b20  (
    .clk(clk_pad),
    .d(addr_if[20]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b21  (
    .clk(clk_pad),
    .d(addr_if[21]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b22  (
    .clk(clk_pad),
    .d(addr_if[22]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b23  (
    .clk(clk_pad),
    .d(addr_if[23]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b24  (
    .clk(clk_pad),
    .d(addr_if[24]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b25  (
    .clk(clk_pad),
    .d(addr_if[25]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b26  (
    .clk(clk_pad),
    .d(addr_if[26]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b27  (
    .clk(clk_pad),
    .d(addr_if[27]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b28  (
    .clk(clk_pad),
    .d(addr_if[28]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b29  (
    .clk(clk_pad),
    .d(addr_if[29]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b30  (
    .clk(clk_pad),
    .d(addr_if[30]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b31  (
    .clk(clk_pad),
    .d(addr_if[31]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b32  (
    .clk(clk_pad),
    .d(addr_if[32]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b33  (
    .clk(clk_pad),
    .d(addr_if[33]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b34  (
    .clk(clk_pad),
    .d(addr_if[34]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b35  (
    .clk(clk_pad),
    .d(addr_if[35]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b36  (
    .clk(clk_pad),
    .d(addr_if[36]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b37  (
    .clk(clk_pad),
    .d(addr_if[37]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b38  (
    .clk(clk_pad),
    .d(addr_if[38]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b39  (
    .clk(clk_pad),
    .d(addr_if[39]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b40  (
    .clk(clk_pad),
    .d(addr_if[40]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b41  (
    .clk(clk_pad),
    .d(addr_if[41]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b42  (
    .clk(clk_pad),
    .d(addr_if[42]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b43  (
    .clk(clk_pad),
    .d(addr_if[43]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b44  (
    .clk(clk_pad),
    .d(addr_if[44]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b45  (
    .clk(clk_pad),
    .d(addr_if[45]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b46  (
    .clk(clk_pad),
    .d(addr_if[46]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b47  (
    .clk(clk_pad),
    .d(addr_if[47]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b48  (
    .clk(clk_pad),
    .d(addr_if[48]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b49  (
    .clk(clk_pad),
    .d(addr_if[49]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b50  (
    .clk(clk_pad),
    .d(addr_if[50]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b51  (
    .clk(clk_pad),
    .d(addr_if[51]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b52  (
    .clk(clk_pad),
    .d(addr_if[52]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b53  (
    .clk(clk_pad),
    .d(addr_if[53]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b54  (
    .clk(clk_pad),
    .d(addr_if[54]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b55  (
    .clk(clk_pad),
    .d(addr_if[55]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b56  (
    .clk(clk_pad),
    .d(addr_if[56]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b57  (
    .clk(clk_pad),
    .d(addr_if[57]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b58  (
    .clk(clk_pad),
    .d(addr_if[58]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b59  (
    .clk(clk_pad),
    .d(addr_if[59]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b60  (
    .clk(clk_pad),
    .d(addr_if[60]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b61  (
    .clk(clk_pad),
    .d(addr_if[61]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b62  (
    .clk(clk_pad),
    .d(addr_if[62]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b63  (
    .clk(clk_pad),
    .d(addr_if[63]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b0  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [0]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b1  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [1]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b10  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [10]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b100  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [100]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [100]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b101  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [101]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [101]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b102  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [102]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [102]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b103  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [103]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [103]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b104  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [104]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [104]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b105  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [105]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [105]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b106  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [106]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [106]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b107  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [107]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [107]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b108  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [108]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [108]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b109  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [109]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [109]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b11  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [11]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b110  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [110]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [110]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b111  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [111]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [111]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b112  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [112]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [112]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b113  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [113]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [113]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b114  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [114]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [114]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b115  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [115]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [115]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b116  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [116]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [116]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b117  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [117]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [117]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b118  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [118]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [118]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b119  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [119]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [119]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b12  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [12]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b120  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [120]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [120]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b121  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [121]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [121]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b122  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [122]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [122]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b123  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [123]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [123]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b124  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [124]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [124]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b125  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [125]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [125]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b126  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [126]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [126]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b127  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [127]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [127]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b13  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [13]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b14  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [14]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b15  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [15]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b16  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [16]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b17  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [17]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b18  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [18]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b19  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [19]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b2  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [2]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b20  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [20]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b21  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [21]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b22  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [22]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b23  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [23]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b24  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [24]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b25  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [25]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b26  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [26]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b27  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [27]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b28  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [28]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b29  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [29]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b3  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [3]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b30  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [30]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b31  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [31]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b32  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [32]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b33  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [33]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b34  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [34]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b35  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [35]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b36  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [36]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b37  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [37]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b38  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [38]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b39  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [39]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b4  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [4]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b40  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [40]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b41  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [41]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b42  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [42]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b43  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [43]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b44  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [44]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b45  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [45]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b46  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [46]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b47  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [47]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b48  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [48]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b49  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [49]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b5  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [5]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b50  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [50]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b51  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [51]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b52  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [52]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b53  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [53]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b54  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [54]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b55  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [55]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b56  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [56]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b57  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [57]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b58  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [58]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b59  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [59]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b6  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [6]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b60  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [60]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b61  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [61]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b62  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [62]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b63  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [63]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b64  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [64]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [64]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b65  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [65]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [65]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b66  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [66]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [66]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b67  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [67]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [67]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b68  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [68]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [68]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b69  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [69]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [69]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b7  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [7]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b70  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [70]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [70]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b71  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [71]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [71]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b72  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [72]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [72]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b73  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [73]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [73]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b74  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [74]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [74]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b75  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [75]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [75]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b76  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [76]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [76]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b77  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [77]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [77]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b78  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [78]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [78]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b79  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [79]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [79]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b8  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [8]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b80  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [80]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [80]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b81  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [81]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [81]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b82  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [82]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [82]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b83  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [83]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [83]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b84  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [84]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [84]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b85  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [85]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [85]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b86  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [86]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [86]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b87  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [87]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [87]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b88  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [88]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [88]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b89  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [89]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [89]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b9  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [9]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b90  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [90]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [90]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b91  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [91]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [91]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b92  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [92]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [92]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b93  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [93]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [93]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b94  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [94]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [94]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b95  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [95]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [95]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b96  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [96]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [96]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b97  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [97]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [97]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b98  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [98]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [98]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b99  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [99]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [99]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b0  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [0]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b1  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [1]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b10  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [10]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b11  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [11]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b12  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [12]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b13  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [13]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b14  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [14]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b15  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [15]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b16  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [16]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b17  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [17]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b18  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [18]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b19  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [19]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b2  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [2]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b20  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [20]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b21  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [21]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b22  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [22]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b23  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [23]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b24  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [24]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b25  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [25]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b26  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [26]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b27  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [27]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b28  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [28]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b29  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [29]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b3  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [3]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b30  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [30]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b31  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [31]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b32  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [32]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b33  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [33]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b34  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [34]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b35  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [35]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b36  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [36]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b37  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [37]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b38  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [38]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b39  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [39]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b4  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [4]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b40  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [40]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b41  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [41]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b42  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [42]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b43  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [43]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b44  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [44]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b45  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [45]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b46  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [46]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b47  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [47]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b48  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [48]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b49  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [49]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b5  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [5]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b50  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [50]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b51  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [51]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b52  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [52]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b53  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [53]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b54  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [54]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b55  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [55]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b56  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [56]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b57  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [57]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b58  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [58]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b59  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [59]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b6  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [6]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b60  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [60]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b61  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [61]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b62  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [62]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b63  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [63]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b7  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n147 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b8  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [8]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b9  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [9]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b12  (
    .clk(clk_pad),
    .d(addr_ex[12]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b13  (
    .clk(clk_pad),
    .d(addr_ex[13]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b14  (
    .clk(clk_pad),
    .d(addr_ex[14]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b15  (
    .clk(clk_pad),
    .d(addr_ex[15]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b16  (
    .clk(clk_pad),
    .d(addr_ex[16]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b17  (
    .clk(clk_pad),
    .d(addr_ex[17]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b18  (
    .clk(clk_pad),
    .d(addr_ex[18]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b19  (
    .clk(clk_pad),
    .d(addr_ex[19]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b20  (
    .clk(clk_pad),
    .d(addr_ex[20]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b21  (
    .clk(clk_pad),
    .d(addr_ex[21]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b22  (
    .clk(clk_pad),
    .d(addr_ex[22]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b23  (
    .clk(clk_pad),
    .d(addr_ex[23]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b24  (
    .clk(clk_pad),
    .d(addr_ex[24]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b25  (
    .clk(clk_pad),
    .d(addr_ex[25]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b26  (
    .clk(clk_pad),
    .d(addr_ex[26]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b27  (
    .clk(clk_pad),
    .d(addr_ex[27]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b28  (
    .clk(clk_pad),
    .d(addr_ex[28]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b29  (
    .clk(clk_pad),
    .d(addr_ex[29]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b30  (
    .clk(clk_pad),
    .d(addr_ex[30]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b31  (
    .clk(clk_pad),
    .d(addr_ex[31]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b32  (
    .clk(clk_pad),
    .d(addr_ex[32]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b33  (
    .clk(clk_pad),
    .d(addr_ex[33]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b34  (
    .clk(clk_pad),
    .d(addr_ex[34]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b35  (
    .clk(clk_pad),
    .d(addr_ex[35]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b36  (
    .clk(clk_pad),
    .d(addr_ex[36]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b37  (
    .clk(clk_pad),
    .d(addr_ex[37]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b38  (
    .clk(clk_pad),
    .d(addr_ex[38]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b39  (
    .clk(clk_pad),
    .d(addr_ex[39]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b40  (
    .clk(clk_pad),
    .d(addr_ex[40]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b41  (
    .clk(clk_pad),
    .d(addr_ex[41]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b42  (
    .clk(clk_pad),
    .d(addr_ex[42]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b43  (
    .clk(clk_pad),
    .d(addr_ex[43]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b44  (
    .clk(clk_pad),
    .d(addr_ex[44]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b45  (
    .clk(clk_pad),
    .d(addr_ex[45]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b46  (
    .clk(clk_pad),
    .d(addr_ex[46]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b47  (
    .clk(clk_pad),
    .d(addr_ex[47]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b48  (
    .clk(clk_pad),
    .d(addr_ex[48]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b49  (
    .clk(clk_pad),
    .d(addr_ex[49]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b50  (
    .clk(clk_pad),
    .d(addr_ex[50]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b51  (
    .clk(clk_pad),
    .d(addr_ex[51]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b52  (
    .clk(clk_pad),
    .d(addr_ex[52]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b53  (
    .clk(clk_pad),
    .d(addr_ex[53]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b54  (
    .clk(clk_pad),
    .d(addr_ex[54]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b55  (
    .clk(clk_pad),
    .d(addr_ex[55]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b56  (
    .clk(clk_pad),
    .d(addr_ex[56]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b57  (
    .clk(clk_pad),
    .d(addr_ex[57]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b58  (
    .clk(clk_pad),
    .d(addr_ex[58]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b59  (
    .clk(clk_pad),
    .d(addr_ex[59]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b60  (
    .clk(clk_pad),
    .d(addr_ex[60]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b61  (
    .clk(clk_pad),
    .d(addr_ex[61]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b62  (
    .clk(clk_pad),
    .d(addr_ex[62]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b63  (
    .clk(clk_pad),
    .d(addr_ex[63]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b0  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [0]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b1  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [1]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b10  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [10]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b100  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [100]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [100]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b101  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [101]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [101]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b102  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [102]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [102]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b103  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [103]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [103]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b104  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [104]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [104]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b105  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [105]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [105]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b106  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [106]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [106]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b107  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [107]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [107]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b108  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [108]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [108]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b109  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [109]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [109]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b11  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [11]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b110  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [110]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [110]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b111  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [111]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [111]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b112  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [112]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [112]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b113  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [113]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [113]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b114  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [114]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [114]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b115  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [115]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [115]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b116  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [116]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [116]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b117  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [117]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [117]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b118  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [118]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [118]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b119  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [119]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [119]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b12  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [12]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b120  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [120]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [120]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b121  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [121]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [121]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b122  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [122]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [122]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b123  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [123]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [123]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b124  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [124]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [124]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b125  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [125]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [125]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b126  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [126]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [126]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b127  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [127]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [127]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b13  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [13]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b14  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [14]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b15  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [15]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b16  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [16]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b17  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [17]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b18  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [18]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b19  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [19]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b2  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [2]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b20  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [20]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b21  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [21]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b22  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [22]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b23  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [23]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b24  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [24]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b25  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [25]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b26  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [26]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b27  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [27]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b28  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [28]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b29  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [29]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b3  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [3]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b30  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [30]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b31  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [31]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b32  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [32]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b33  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [33]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b34  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [34]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b35  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [35]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b36  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [36]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b37  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [37]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b38  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [38]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b39  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [39]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b4  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [4]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b40  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [40]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b41  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [41]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b42  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [42]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b43  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [43]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b44  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [44]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b45  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [45]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b46  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [46]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b47  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [47]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b48  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [48]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b49  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [49]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b5  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [5]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b50  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [50]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b51  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [51]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b52  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [52]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b53  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [53]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b54  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [54]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b55  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [55]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b56  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [56]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b57  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [57]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b58  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [58]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b59  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [59]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b6  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [6]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b60  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [60]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b61  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [61]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b62  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [62]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b63  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [63]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b64  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [64]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [64]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b65  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [65]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [65]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b66  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [66]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [66]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b67  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [67]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [67]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b68  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [68]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [68]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b69  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [69]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [69]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b7  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [7]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b70  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [70]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [70]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b71  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [71]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [71]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b72  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [72]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [72]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b73  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [73]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [73]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b74  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [74]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [74]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b75  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [75]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [75]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b76  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [76]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [76]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b77  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [77]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [77]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b78  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [78]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [78]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b79  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [79]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [79]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b8  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [8]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b80  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [80]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [80]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b81  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [81]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [81]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b82  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [82]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [82]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b83  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [83]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [83]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b84  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [84]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [84]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b85  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [85]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [85]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b86  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [86]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [86]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b87  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [87]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [87]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b88  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [88]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [88]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b89  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [89]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [89]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b9  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [9]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b90  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [90]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [90]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b91  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [91]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [91]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b92  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [92]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [92]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b93  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [93]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [93]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b94  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [94]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [94]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b95  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [95]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [95]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b96  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [96]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [96]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b97  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [97]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [97]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b98  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [98]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [98]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b99  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pa_temp [99]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [99]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b0  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [0]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b1  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [1]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b10  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [10]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b11  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [11]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b12  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [12]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b13  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [13]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b14  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [14]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b15  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [15]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b16  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [16]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b17  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [17]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b18  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [18]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b19  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [19]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b2  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [2]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b20  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [20]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b21  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [21]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b22  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [22]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b23  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [23]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b24  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [24]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b25  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [25]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b26  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [26]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b27  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [27]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b28  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [28]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b29  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [29]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b3  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [3]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b30  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [30]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b31  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [31]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b32  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [32]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b33  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [33]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b34  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [34]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b35  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [35]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b36  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [36]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b37  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [37]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b38  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [38]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b39  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [39]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b4  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [4]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b40  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [40]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b41  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [41]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b42  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [42]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b43  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [43]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b44  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [44]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b45  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [45]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b46  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [46]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b47  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [47]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b48  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [48]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b49  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [49]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b5  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [5]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b50  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [50]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b51  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [51]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b52  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [52]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b53  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [53]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b54  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [54]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b55  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [55]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b56  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [56]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b57  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [57]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b58  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [58]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b59  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [59]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b6  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [6]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b60  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [60]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b61  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [61]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b62  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [62]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b63  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [63]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b7  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n158 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b8  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [8]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b9  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/pte_temp [9]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b0  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b1  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b10  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b100  (
    .clk(clk_pad),
    .d(\biu/paddress [100]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [100]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b101  (
    .clk(clk_pad),
    .d(\biu/paddress [101]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [101]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b102  (
    .clk(clk_pad),
    .d(\biu/paddress [102]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [102]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b103  (
    .clk(clk_pad),
    .d(\biu/paddress [103]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [103]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b104  (
    .clk(clk_pad),
    .d(\biu/paddress [104]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [104]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b105  (
    .clk(clk_pad),
    .d(\biu/paddress [105]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [105]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b106  (
    .clk(clk_pad),
    .d(\biu/paddress [106]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [106]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b107  (
    .clk(clk_pad),
    .d(\biu/paddress [107]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [107]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b108  (
    .clk(clk_pad),
    .d(\biu/paddress [108]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [108]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b109  (
    .clk(clk_pad),
    .d(\biu/paddress [109]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [109]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b11  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b110  (
    .clk(clk_pad),
    .d(\biu/paddress [110]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [110]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b111  (
    .clk(clk_pad),
    .d(\biu/paddress [111]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [111]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b112  (
    .clk(clk_pad),
    .d(\biu/paddress [112]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [112]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b113  (
    .clk(clk_pad),
    .d(\biu/paddress [113]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [113]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b114  (
    .clk(clk_pad),
    .d(\biu/paddress [114]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [114]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b115  (
    .clk(clk_pad),
    .d(\biu/paddress [115]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [115]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b116  (
    .clk(clk_pad),
    .d(\biu/paddress [116]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [116]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b117  (
    .clk(clk_pad),
    .d(\biu/paddress [117]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [117]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b118  (
    .clk(clk_pad),
    .d(\biu/paddress [118]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [118]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b119  (
    .clk(clk_pad),
    .d(\biu/paddress [119]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [119]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b12  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b120  (
    .clk(clk_pad),
    .d(\biu/paddress [120]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [120]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b121  (
    .clk(clk_pad),
    .d(\biu/paddress [121]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [121]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b122  (
    .clk(clk_pad),
    .d(\biu/paddress [122]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [122]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b123  (
    .clk(clk_pad),
    .d(\biu/paddress [123]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [123]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b124  (
    .clk(clk_pad),
    .d(\biu/paddress [124]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [124]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b125  (
    .clk(clk_pad),
    .d(\biu/paddress [125]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [125]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b126  (
    .clk(clk_pad),
    .d(\biu/paddress [126]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [126]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b127  (
    .clk(clk_pad),
    .d(\biu/paddress [127]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [127]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b13  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b14  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b15  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b16  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b17  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b18  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b19  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b2  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b20  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b21  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b22  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b23  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b24  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b25  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b26  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b27  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b28  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b29  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b3  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b30  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b31  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b32  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b33  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b34  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b35  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b36  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b37  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b38  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b39  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b4  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b40  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b41  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b42  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b43  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b44  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b45  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b46  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b47  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b48  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b49  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b5  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b50  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b51  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b52  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b53  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b54  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b55  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b56  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b57  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b58  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b59  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b6  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b60  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b61  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b62  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b63  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b64  (
    .clk(clk_pad),
    .d(\biu/paddress [64]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [64]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b65  (
    .clk(clk_pad),
    .d(\biu/paddress [65]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [65]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b66  (
    .clk(clk_pad),
    .d(\biu/paddress [66]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [66]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b67  (
    .clk(clk_pad),
    .d(\biu/paddress [67]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [67]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b68  (
    .clk(clk_pad),
    .d(\biu/paddress [68]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [68]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b69  (
    .clk(clk_pad),
    .d(\biu/paddress [69]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [69]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b7  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b70  (
    .clk(clk_pad),
    .d(\biu/paddress [70]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [70]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b71  (
    .clk(clk_pad),
    .d(\biu/paddress [71]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [71]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b72  (
    .clk(clk_pad),
    .d(\biu/paddress [72]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [72]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b73  (
    .clk(clk_pad),
    .d(\biu/paddress [73]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [73]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b74  (
    .clk(clk_pad),
    .d(\biu/paddress [74]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [74]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b75  (
    .clk(clk_pad),
    .d(\biu/paddress [75]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [75]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b76  (
    .clk(clk_pad),
    .d(\biu/paddress [76]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [76]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b77  (
    .clk(clk_pad),
    .d(\biu/paddress [77]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [77]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b78  (
    .clk(clk_pad),
    .d(\biu/paddress [78]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [78]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b79  (
    .clk(clk_pad),
    .d(\biu/paddress [79]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [79]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b8  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b80  (
    .clk(clk_pad),
    .d(\biu/paddress [80]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [80]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b81  (
    .clk(clk_pad),
    .d(\biu/paddress [81]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [81]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b82  (
    .clk(clk_pad),
    .d(\biu/paddress [82]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [82]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b83  (
    .clk(clk_pad),
    .d(\biu/paddress [83]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [83]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b84  (
    .clk(clk_pad),
    .d(\biu/paddress [84]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [84]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b85  (
    .clk(clk_pad),
    .d(\biu/paddress [85]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [85]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b86  (
    .clk(clk_pad),
    .d(\biu/paddress [86]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [86]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b87  (
    .clk(clk_pad),
    .d(\biu/paddress [87]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [87]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b88  (
    .clk(clk_pad),
    .d(\biu/paddress [88]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [88]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b89  (
    .clk(clk_pad),
    .d(\biu/paddress [89]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [89]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b9  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n166 [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b90  (
    .clk(clk_pad),
    .d(\biu/paddress [90]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [90]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b91  (
    .clk(clk_pad),
    .d(\biu/paddress [91]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [91]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b92  (
    .clk(clk_pad),
    .d(\biu/paddress [92]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [92]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b93  (
    .clk(clk_pad),
    .d(\biu/paddress [93]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [93]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b94  (
    .clk(clk_pad),
    .d(\biu/paddress [94]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [94]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b95  (
    .clk(clk_pad),
    .d(\biu/paddress [95]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [95]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b96  (
    .clk(clk_pad),
    .d(\biu/paddress [96]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [96]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b97  (
    .clk(clk_pad),
    .d(\biu/paddress [97]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [97]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b98  (
    .clk(clk_pad),
    .d(\biu/paddress [98]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [98]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b99  (
    .clk(clk_pad),
    .d(\biu/paddress [99]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [99]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b0  (
    .clk(clk_pad),
    .d(uncache_data[0]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b1  (
    .clk(clk_pad),
    .d(uncache_data[1]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b10  (
    .clk(clk_pad),
    .d(uncache_data[10]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b11  (
    .clk(clk_pad),
    .d(uncache_data[11]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b12  (
    .clk(clk_pad),
    .d(uncache_data[12]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b13  (
    .clk(clk_pad),
    .d(uncache_data[13]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b14  (
    .clk(clk_pad),
    .d(uncache_data[14]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b15  (
    .clk(clk_pad),
    .d(uncache_data[15]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b16  (
    .clk(clk_pad),
    .d(uncache_data[16]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b17  (
    .clk(clk_pad),
    .d(uncache_data[17]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b18  (
    .clk(clk_pad),
    .d(uncache_data[18]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b19  (
    .clk(clk_pad),
    .d(uncache_data[19]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b2  (
    .clk(clk_pad),
    .d(uncache_data[2]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b20  (
    .clk(clk_pad),
    .d(uncache_data[20]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b21  (
    .clk(clk_pad),
    .d(uncache_data[21]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b22  (
    .clk(clk_pad),
    .d(uncache_data[22]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b23  (
    .clk(clk_pad),
    .d(uncache_data[23]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b24  (
    .clk(clk_pad),
    .d(uncache_data[24]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b25  (
    .clk(clk_pad),
    .d(uncache_data[25]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b26  (
    .clk(clk_pad),
    .d(uncache_data[26]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b27  (
    .clk(clk_pad),
    .d(uncache_data[27]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b28  (
    .clk(clk_pad),
    .d(uncache_data[28]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b29  (
    .clk(clk_pad),
    .d(uncache_data[29]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b3  (
    .clk(clk_pad),
    .d(uncache_data[3]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b30  (
    .clk(clk_pad),
    .d(uncache_data[30]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b31  (
    .clk(clk_pad),
    .d(uncache_data[31]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b32  (
    .clk(clk_pad),
    .d(uncache_data[32]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b33  (
    .clk(clk_pad),
    .d(uncache_data[33]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b34  (
    .clk(clk_pad),
    .d(uncache_data[34]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b35  (
    .clk(clk_pad),
    .d(uncache_data[35]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b36  (
    .clk(clk_pad),
    .d(uncache_data[36]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b37  (
    .clk(clk_pad),
    .d(uncache_data[37]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b38  (
    .clk(clk_pad),
    .d(uncache_data[38]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b39  (
    .clk(clk_pad),
    .d(uncache_data[39]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b4  (
    .clk(clk_pad),
    .d(uncache_data[4]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b40  (
    .clk(clk_pad),
    .d(uncache_data[40]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b41  (
    .clk(clk_pad),
    .d(uncache_data[41]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b42  (
    .clk(clk_pad),
    .d(uncache_data[42]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b43  (
    .clk(clk_pad),
    .d(uncache_data[43]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b44  (
    .clk(clk_pad),
    .d(uncache_data[44]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b45  (
    .clk(clk_pad),
    .d(uncache_data[45]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b46  (
    .clk(clk_pad),
    .d(uncache_data[46]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b47  (
    .clk(clk_pad),
    .d(uncache_data[47]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b48  (
    .clk(clk_pad),
    .d(uncache_data[48]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b49  (
    .clk(clk_pad),
    .d(uncache_data[49]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b5  (
    .clk(clk_pad),
    .d(uncache_data[5]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b50  (
    .clk(clk_pad),
    .d(uncache_data[50]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b51  (
    .clk(clk_pad),
    .d(uncache_data[51]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b52  (
    .clk(clk_pad),
    .d(uncache_data[52]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b53  (
    .clk(clk_pad),
    .d(uncache_data[53]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b54  (
    .clk(clk_pad),
    .d(uncache_data[54]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b55  (
    .clk(clk_pad),
    .d(uncache_data[55]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b56  (
    .clk(clk_pad),
    .d(uncache_data[56]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b57  (
    .clk(clk_pad),
    .d(uncache_data[57]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b58  (
    .clk(clk_pad),
    .d(uncache_data[58]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b59  (
    .clk(clk_pad),
    .d(uncache_data[59]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b6  (
    .clk(clk_pad),
    .d(uncache_data[6]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b60  (
    .clk(clk_pad),
    .d(uncache_data[60]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b61  (
    .clk(clk_pad),
    .d(uncache_data[61]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b62  (
    .clk(clk_pad),
    .d(uncache_data[62]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b63  (
    .clk(clk_pad),
    .d(uncache_data[63]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b7  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n165 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b8  (
    .clk(clk_pad),
    .d(uncache_data[8]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b9  (
    .clk(clk_pad),
    .d(uncache_data[9]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg8_b0  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n132[0]_d ),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/statu [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg8_b1  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n131[1]_d ),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/statu [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg8_b2  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n132 [2]),
    .en(1'b1),
    .reset(~\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/statu [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg8_b3  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n132 [3]),
    .en(1'b1),
    .reset(~\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/statu [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg8_b4  (
    .clk(clk_pad),
    .d(\biu/cache_ctrl_logic/n127[4]_d ),
    .en(1'b1),
    .reset(~\biu/cache_ctrl_logic/mux44_b4_sel_is_2_o ),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/statu [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("DISABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u0  (
    .a(\cu_ru/tvec [4]),
    .b(\cu_ru/trap_cause [0]),
    .c(\cu_ru/add0_2/c0 ),
    .o({\cu_ru/add0_2/c1 ,\cu_ru/n43 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u1  (
    .a(\cu_ru/tvec [5]),
    .b(\cu_ru/trap_cause [1]),
    .c(\cu_ru/add0_2/c1 ),
    .o({\cu_ru/add0_2/c2 ,\cu_ru/n43 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u10  (
    .a(\cu_ru/tvec [14]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c10 ),
    .o({\cu_ru/add0_2/c11 ,\cu_ru/n43 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u11  (
    .a(\cu_ru/tvec [15]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c11 ),
    .o({\cu_ru/add0_2/c12 ,\cu_ru/n43 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u12  (
    .a(\cu_ru/tvec [16]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c12 ),
    .o({\cu_ru/add0_2/c13 ,\cu_ru/n43 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u13  (
    .a(\cu_ru/tvec [17]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c13 ),
    .o({\cu_ru/add0_2/c14 ,\cu_ru/n43 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u14  (
    .a(\cu_ru/tvec [18]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c14 ),
    .o({\cu_ru/add0_2/c15 ,\cu_ru/n43 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u15  (
    .a(\cu_ru/tvec [19]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c15 ),
    .o({\cu_ru/add0_2/c16 ,\cu_ru/n43 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u16  (
    .a(\cu_ru/tvec [20]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c16 ),
    .o({\cu_ru/add0_2/c17 ,\cu_ru/n43 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u17  (
    .a(\cu_ru/tvec [21]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c17 ),
    .o({\cu_ru/add0_2/c18 ,\cu_ru/n43 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u18  (
    .a(\cu_ru/tvec [22]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c18 ),
    .o({\cu_ru/add0_2/c19 ,\cu_ru/n43 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u19  (
    .a(\cu_ru/tvec [23]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c19 ),
    .o({\cu_ru/add0_2/c20 ,\cu_ru/n43 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u2  (
    .a(\cu_ru/tvec [6]),
    .b(\cu_ru/trap_cause [2]),
    .c(\cu_ru/add0_2/c2 ),
    .o({\cu_ru/add0_2/c3 ,\cu_ru/n43 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u20  (
    .a(\cu_ru/tvec [24]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c20 ),
    .o({\cu_ru/add0_2/c21 ,\cu_ru/n43 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u21  (
    .a(\cu_ru/tvec [25]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c21 ),
    .o({\cu_ru/add0_2/c22 ,\cu_ru/n43 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u22  (
    .a(\cu_ru/tvec [26]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c22 ),
    .o({\cu_ru/add0_2/c23 ,\cu_ru/n43 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u23  (
    .a(\cu_ru/tvec [27]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c23 ),
    .o({\cu_ru/add0_2/c24 ,\cu_ru/n43 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u24  (
    .a(\cu_ru/tvec [28]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c24 ),
    .o({\cu_ru/add0_2/c25 ,\cu_ru/n43 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u25  (
    .a(\cu_ru/tvec [29]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c25 ),
    .o({\cu_ru/add0_2/c26 ,\cu_ru/n43 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u26  (
    .a(\cu_ru/tvec [30]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c26 ),
    .o({\cu_ru/add0_2/c27 ,\cu_ru/n43 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u27  (
    .a(\cu_ru/tvec [31]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c27 ),
    .o({\cu_ru/add0_2/c28 ,\cu_ru/n43 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u28  (
    .a(\cu_ru/tvec [32]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c28 ),
    .o({\cu_ru/add0_2/c29 ,\cu_ru/n43 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u29  (
    .a(\cu_ru/tvec [33]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c29 ),
    .o({\cu_ru/add0_2/c30 ,\cu_ru/n43 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u3  (
    .a(\cu_ru/tvec [7]),
    .b(\cu_ru/trap_cause [3]),
    .c(\cu_ru/add0_2/c3 ),
    .o({\cu_ru/add0_2/c4 ,\cu_ru/n43 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u30  (
    .a(\cu_ru/tvec [34]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c30 ),
    .o({\cu_ru/add0_2/c31 ,\cu_ru/n43 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u31  (
    .a(\cu_ru/tvec [35]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c31 ),
    .o({\cu_ru/add0_2/c32 ,\cu_ru/n43 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u32  (
    .a(\cu_ru/tvec [36]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c32 ),
    .o({\cu_ru/add0_2/c33 ,\cu_ru/n43 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u33  (
    .a(\cu_ru/tvec [37]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c33 ),
    .o({\cu_ru/add0_2/c34 ,\cu_ru/n43 [33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u34  (
    .a(\cu_ru/tvec [38]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c34 ),
    .o({\cu_ru/add0_2/c35 ,\cu_ru/n43 [34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u35  (
    .a(\cu_ru/tvec [39]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c35 ),
    .o({\cu_ru/add0_2/c36 ,\cu_ru/n43 [35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u36  (
    .a(\cu_ru/tvec [40]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c36 ),
    .o({\cu_ru/add0_2/c37 ,\cu_ru/n43 [36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u37  (
    .a(\cu_ru/tvec [41]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c37 ),
    .o({\cu_ru/add0_2/c38 ,\cu_ru/n43 [37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u38  (
    .a(\cu_ru/tvec [42]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c38 ),
    .o({\cu_ru/add0_2/c39 ,\cu_ru/n43 [38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u39  (
    .a(\cu_ru/tvec [43]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c39 ),
    .o({\cu_ru/add0_2/c40 ,\cu_ru/n43 [39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u4  (
    .a(\cu_ru/tvec [8]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c4 ),
    .o({\cu_ru/add0_2/c5 ,\cu_ru/n43 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u40  (
    .a(\cu_ru/tvec [44]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c40 ),
    .o({\cu_ru/add0_2/c41 ,\cu_ru/n43 [40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u41  (
    .a(\cu_ru/tvec [45]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c41 ),
    .o({\cu_ru/add0_2/c42 ,\cu_ru/n43 [41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u42  (
    .a(\cu_ru/tvec [46]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c42 ),
    .o({\cu_ru/add0_2/c43 ,\cu_ru/n43 [42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u43  (
    .a(\cu_ru/tvec [47]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c43 ),
    .o({\cu_ru/add0_2/c44 ,\cu_ru/n43 [43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u44  (
    .a(\cu_ru/tvec [48]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c44 ),
    .o({\cu_ru/add0_2/c45 ,\cu_ru/n43 [44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u45  (
    .a(\cu_ru/tvec [49]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c45 ),
    .o({\cu_ru/add0_2/c46 ,\cu_ru/n43 [45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u46  (
    .a(\cu_ru/tvec [50]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c46 ),
    .o({\cu_ru/add0_2/c47 ,\cu_ru/n43 [46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u47  (
    .a(\cu_ru/tvec [51]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c47 ),
    .o({\cu_ru/add0_2/c48 ,\cu_ru/n43 [47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u48  (
    .a(\cu_ru/tvec [52]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c48 ),
    .o({\cu_ru/add0_2/c49 ,\cu_ru/n43 [48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u49  (
    .a(\cu_ru/tvec [53]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c49 ),
    .o({\cu_ru/add0_2/c50 ,\cu_ru/n43 [49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u5  (
    .a(\cu_ru/tvec [9]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c5 ),
    .o({\cu_ru/add0_2/c6 ,\cu_ru/n43 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u50  (
    .a(\cu_ru/tvec [54]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c50 ),
    .o({\cu_ru/add0_2/c51 ,\cu_ru/n43 [50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u51  (
    .a(\cu_ru/tvec [55]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c51 ),
    .o({\cu_ru/add0_2/c52 ,\cu_ru/n43 [51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u52  (
    .a(\cu_ru/tvec [56]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c52 ),
    .o({\cu_ru/add0_2/c53 ,\cu_ru/n43 [52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u53  (
    .a(\cu_ru/tvec [57]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c53 ),
    .o({\cu_ru/add0_2/c54 ,\cu_ru/n43 [53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u54  (
    .a(\cu_ru/tvec [58]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c54 ),
    .o({\cu_ru/add0_2/c55 ,\cu_ru/n43 [54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u55  (
    .a(\cu_ru/tvec [59]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c55 ),
    .o({\cu_ru/add0_2/c56 ,\cu_ru/n43 [55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u56  (
    .a(\cu_ru/tvec [60]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c56 ),
    .o({\cu_ru/add0_2/c57 ,\cu_ru/n43 [56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u57  (
    .a(\cu_ru/tvec [61]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c57 ),
    .o({\cu_ru/add0_2/c58 ,\cu_ru/n43 [57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u58  (
    .a(\cu_ru/tvec [62]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c58 ),
    .o({\cu_ru/add0_2/c59 ,\cu_ru/n43 [58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u59  (
    .a(\cu_ru/tvec [63]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c59 ),
    .o({\cu_ru/add0_2/c60 ,\cu_ru/n43 [59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u6  (
    .a(\cu_ru/tvec [10]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c6 ),
    .o({\cu_ru/add0_2/c7 ,\cu_ru/n43 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u7  (
    .a(\cu_ru/tvec [11]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c7 ),
    .o({\cu_ru/add0_2/c8 ,\cu_ru/n43 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u8  (
    .a(\cu_ru/tvec [12]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c8 ),
    .o({\cu_ru/add0_2/c9 ,\cu_ru/n43 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/u9  (
    .a(\cu_ru/tvec [13]),
    .b(1'b0),
    .c(\cu_ru/add0_2/c9 ),
    .o({\cu_ru/add0_2/c10 ,\cu_ru/n43 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \cu_ru/add0_2/ucin  (
    .a(1'b0),
    .o({\cu_ru/add0_2/c0 ,open_n6062}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/add0_2/ucout  (
    .c(\cu_ru/add0_2/c60 ),
    .o({open_n6065,\cu_ru/add0_2_co }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c0  (
    .di(data_rd[3:0]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_003 ,\cu_ru/al_ram_gpr_al_u0_do_i0_002 ,\cu_ru/al_ram_gpr_al_u0_do_i0_001 ,\cu_ru/al_ram_gpr_al_u0_do_i0_000 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c1  (
    .di(data_rd[7:4]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_007 ,\cu_ru/al_ram_gpr_al_u0_do_i0_006 ,\cu_ru/al_ram_gpr_al_u0_do_i0_005 ,\cu_ru/al_ram_gpr_al_u0_do_i0_004 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c10  (
    .di(data_rd[43:40]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_043 ,\cu_ru/al_ram_gpr_al_u0_do_i0_042 ,\cu_ru/al_ram_gpr_al_u0_do_i0_041 ,\cu_ru/al_ram_gpr_al_u0_do_i0_040 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c11  (
    .di(data_rd[47:44]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_047 ,\cu_ru/al_ram_gpr_al_u0_do_i0_046 ,\cu_ru/al_ram_gpr_al_u0_do_i0_045 ,\cu_ru/al_ram_gpr_al_u0_do_i0_044 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c12  (
    .di(data_rd[51:48]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_051 ,\cu_ru/al_ram_gpr_al_u0_do_i0_050 ,\cu_ru/al_ram_gpr_al_u0_do_i0_049 ,\cu_ru/al_ram_gpr_al_u0_do_i0_048 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c13  (
    .di(data_rd[55:52]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_055 ,\cu_ru/al_ram_gpr_al_u0_do_i0_054 ,\cu_ru/al_ram_gpr_al_u0_do_i0_053 ,\cu_ru/al_ram_gpr_al_u0_do_i0_052 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c14  (
    .di(data_rd[59:56]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_059 ,\cu_ru/al_ram_gpr_al_u0_do_i0_058 ,\cu_ru/al_ram_gpr_al_u0_do_i0_057 ,\cu_ru/al_ram_gpr_al_u0_do_i0_056 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c15  (
    .di(data_rd[63:60]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_063 ,\cu_ru/al_ram_gpr_al_u0_do_i0_062 ,\cu_ru/al_ram_gpr_al_u0_do_i0_061 ,\cu_ru/al_ram_gpr_al_u0_do_i0_060 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c2  (
    .di(data_rd[11:8]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_011 ,\cu_ru/al_ram_gpr_al_u0_do_i0_010 ,\cu_ru/al_ram_gpr_al_u0_do_i0_009 ,\cu_ru/al_ram_gpr_al_u0_do_i0_008 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c3  (
    .di(data_rd[15:12]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_015 ,\cu_ru/al_ram_gpr_al_u0_do_i0_014 ,\cu_ru/al_ram_gpr_al_u0_do_i0_013 ,\cu_ru/al_ram_gpr_al_u0_do_i0_012 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c4  (
    .di(data_rd[19:16]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_019 ,\cu_ru/al_ram_gpr_al_u0_do_i0_018 ,\cu_ru/al_ram_gpr_al_u0_do_i0_017 ,\cu_ru/al_ram_gpr_al_u0_do_i0_016 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c5  (
    .di(data_rd[23:20]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_023 ,\cu_ru/al_ram_gpr_al_u0_do_i0_022 ,\cu_ru/al_ram_gpr_al_u0_do_i0_021 ,\cu_ru/al_ram_gpr_al_u0_do_i0_020 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c6  (
    .di(data_rd[27:24]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_027 ,\cu_ru/al_ram_gpr_al_u0_do_i0_026 ,\cu_ru/al_ram_gpr_al_u0_do_i0_025 ,\cu_ru/al_ram_gpr_al_u0_do_i0_024 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c7  (
    .di(data_rd[31:28]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_031 ,\cu_ru/al_ram_gpr_al_u0_do_i0_030 ,\cu_ru/al_ram_gpr_al_u0_do_i0_029 ,\cu_ru/al_ram_gpr_al_u0_do_i0_028 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c8  (
    .di(data_rd[35:32]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_035 ,\cu_ru/al_ram_gpr_al_u0_do_i0_034 ,\cu_ru/al_ram_gpr_al_u0_do_i0_033 ,\cu_ru/al_ram_gpr_al_u0_do_i0_032 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r0_c9  (
    .di(data_rd[39:36]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i0_039 ,\cu_ru/al_ram_gpr_al_u0_do_i0_038 ,\cu_ru/al_ram_gpr_al_u0_do_i0_037 ,\cu_ru/al_ram_gpr_al_u0_do_i0_036 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c0  (
    .di(data_rd[3:0]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_003 ,\cu_ru/al_ram_gpr_al_u0_do_i1_002 ,\cu_ru/al_ram_gpr_al_u0_do_i1_001 ,\cu_ru/al_ram_gpr_al_u0_do_i1_000 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c1  (
    .di(data_rd[7:4]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_007 ,\cu_ru/al_ram_gpr_al_u0_do_i1_006 ,\cu_ru/al_ram_gpr_al_u0_do_i1_005 ,\cu_ru/al_ram_gpr_al_u0_do_i1_004 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c10  (
    .di(data_rd[43:40]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_043 ,\cu_ru/al_ram_gpr_al_u0_do_i1_042 ,\cu_ru/al_ram_gpr_al_u0_do_i1_041 ,\cu_ru/al_ram_gpr_al_u0_do_i1_040 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c11  (
    .di(data_rd[47:44]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_047 ,\cu_ru/al_ram_gpr_al_u0_do_i1_046 ,\cu_ru/al_ram_gpr_al_u0_do_i1_045 ,\cu_ru/al_ram_gpr_al_u0_do_i1_044 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c12  (
    .di(data_rd[51:48]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_051 ,\cu_ru/al_ram_gpr_al_u0_do_i1_050 ,\cu_ru/al_ram_gpr_al_u0_do_i1_049 ,\cu_ru/al_ram_gpr_al_u0_do_i1_048 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c13  (
    .di(data_rd[55:52]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_055 ,\cu_ru/al_ram_gpr_al_u0_do_i1_054 ,\cu_ru/al_ram_gpr_al_u0_do_i1_053 ,\cu_ru/al_ram_gpr_al_u0_do_i1_052 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c14  (
    .di(data_rd[59:56]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_059 ,\cu_ru/al_ram_gpr_al_u0_do_i1_058 ,\cu_ru/al_ram_gpr_al_u0_do_i1_057 ,\cu_ru/al_ram_gpr_al_u0_do_i1_056 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c15  (
    .di(data_rd[63:60]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_063 ,\cu_ru/al_ram_gpr_al_u0_do_i1_062 ,\cu_ru/al_ram_gpr_al_u0_do_i1_061 ,\cu_ru/al_ram_gpr_al_u0_do_i1_060 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c2  (
    .di(data_rd[11:8]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_011 ,\cu_ru/al_ram_gpr_al_u0_do_i1_010 ,\cu_ru/al_ram_gpr_al_u0_do_i1_009 ,\cu_ru/al_ram_gpr_al_u0_do_i1_008 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c3  (
    .di(data_rd[15:12]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_015 ,\cu_ru/al_ram_gpr_al_u0_do_i1_014 ,\cu_ru/al_ram_gpr_al_u0_do_i1_013 ,\cu_ru/al_ram_gpr_al_u0_do_i1_012 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c4  (
    .di(data_rd[19:16]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_019 ,\cu_ru/al_ram_gpr_al_u0_do_i1_018 ,\cu_ru/al_ram_gpr_al_u0_do_i1_017 ,\cu_ru/al_ram_gpr_al_u0_do_i1_016 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c5  (
    .di(data_rd[23:20]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_023 ,\cu_ru/al_ram_gpr_al_u0_do_i1_022 ,\cu_ru/al_ram_gpr_al_u0_do_i1_021 ,\cu_ru/al_ram_gpr_al_u0_do_i1_020 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c6  (
    .di(data_rd[27:24]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_027 ,\cu_ru/al_ram_gpr_al_u0_do_i1_026 ,\cu_ru/al_ram_gpr_al_u0_do_i1_025 ,\cu_ru/al_ram_gpr_al_u0_do_i1_024 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c7  (
    .di(data_rd[31:28]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_031 ,\cu_ru/al_ram_gpr_al_u0_do_i1_030 ,\cu_ru/al_ram_gpr_al_u0_do_i1_029 ,\cu_ru/al_ram_gpr_al_u0_do_i1_028 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c8  (
    .di(data_rd[35:32]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_035 ,\cu_ru/al_ram_gpr_al_u0_do_i1_034 ,\cu_ru/al_ram_gpr_al_u0_do_i1_033 ,\cu_ru/al_ram_gpr_al_u0_do_i1_032 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_al_u0_r1_c9  (
    .di(data_rd[39:36]),
    .raddr(\cu_ru/n49 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_al_u0_do_i1_039 ,\cu_ru/al_ram_gpr_al_u0_do_i1_038 ,\cu_ru/al_ram_gpr_al_u0_do_i1_037 ,\cu_ru/al_ram_gpr_al_u0_do_i1_036 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c0  (
    .di(data_rd[3:0]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_003 ,\cu_ru/al_ram_gpr_do_i0_002 ,\cu_ru/al_ram_gpr_do_i0_001 ,\cu_ru/al_ram_gpr_do_i0_000 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c1  (
    .di(data_rd[7:4]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_007 ,\cu_ru/al_ram_gpr_do_i0_006 ,\cu_ru/al_ram_gpr_do_i0_005 ,\cu_ru/al_ram_gpr_do_i0_004 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c10  (
    .di(data_rd[43:40]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_043 ,\cu_ru/al_ram_gpr_do_i0_042 ,\cu_ru/al_ram_gpr_do_i0_041 ,\cu_ru/al_ram_gpr_do_i0_040 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c11  (
    .di(data_rd[47:44]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_047 ,\cu_ru/al_ram_gpr_do_i0_046 ,\cu_ru/al_ram_gpr_do_i0_045 ,\cu_ru/al_ram_gpr_do_i0_044 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c12  (
    .di(data_rd[51:48]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_051 ,\cu_ru/al_ram_gpr_do_i0_050 ,\cu_ru/al_ram_gpr_do_i0_049 ,\cu_ru/al_ram_gpr_do_i0_048 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c13  (
    .di(data_rd[55:52]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_055 ,\cu_ru/al_ram_gpr_do_i0_054 ,\cu_ru/al_ram_gpr_do_i0_053 ,\cu_ru/al_ram_gpr_do_i0_052 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c14  (
    .di(data_rd[59:56]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_059 ,\cu_ru/al_ram_gpr_do_i0_058 ,\cu_ru/al_ram_gpr_do_i0_057 ,\cu_ru/al_ram_gpr_do_i0_056 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c15  (
    .di(data_rd[63:60]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_063 ,\cu_ru/al_ram_gpr_do_i0_062 ,\cu_ru/al_ram_gpr_do_i0_061 ,\cu_ru/al_ram_gpr_do_i0_060 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c2  (
    .di(data_rd[11:8]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_011 ,\cu_ru/al_ram_gpr_do_i0_010 ,\cu_ru/al_ram_gpr_do_i0_009 ,\cu_ru/al_ram_gpr_do_i0_008 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c3  (
    .di(data_rd[15:12]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_015 ,\cu_ru/al_ram_gpr_do_i0_014 ,\cu_ru/al_ram_gpr_do_i0_013 ,\cu_ru/al_ram_gpr_do_i0_012 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c4  (
    .di(data_rd[19:16]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_019 ,\cu_ru/al_ram_gpr_do_i0_018 ,\cu_ru/al_ram_gpr_do_i0_017 ,\cu_ru/al_ram_gpr_do_i0_016 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c5  (
    .di(data_rd[23:20]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_023 ,\cu_ru/al_ram_gpr_do_i0_022 ,\cu_ru/al_ram_gpr_do_i0_021 ,\cu_ru/al_ram_gpr_do_i0_020 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c6  (
    .di(data_rd[27:24]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_027 ,\cu_ru/al_ram_gpr_do_i0_026 ,\cu_ru/al_ram_gpr_do_i0_025 ,\cu_ru/al_ram_gpr_do_i0_024 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c7  (
    .di(data_rd[31:28]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_031 ,\cu_ru/al_ram_gpr_do_i0_030 ,\cu_ru/al_ram_gpr_do_i0_029 ,\cu_ru/al_ram_gpr_do_i0_028 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c8  (
    .di(data_rd[35:32]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_035 ,\cu_ru/al_ram_gpr_do_i0_034 ,\cu_ru/al_ram_gpr_do_i0_033 ,\cu_ru/al_ram_gpr_do_i0_032 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r0_c9  (
    .di(data_rd[39:36]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_0_al_n1985 ),
    .do({\cu_ru/al_ram_gpr_do_i0_039 ,\cu_ru/al_ram_gpr_do_i0_038 ,\cu_ru/al_ram_gpr_do_i0_037 ,\cu_ru/al_ram_gpr_do_i0_036 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c0  (
    .di(data_rd[3:0]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_003 ,\cu_ru/al_ram_gpr_do_i1_002 ,\cu_ru/al_ram_gpr_do_i1_001 ,\cu_ru/al_ram_gpr_do_i1_000 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c1  (
    .di(data_rd[7:4]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_007 ,\cu_ru/al_ram_gpr_do_i1_006 ,\cu_ru/al_ram_gpr_do_i1_005 ,\cu_ru/al_ram_gpr_do_i1_004 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c10  (
    .di(data_rd[43:40]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_043 ,\cu_ru/al_ram_gpr_do_i1_042 ,\cu_ru/al_ram_gpr_do_i1_041 ,\cu_ru/al_ram_gpr_do_i1_040 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c11  (
    .di(data_rd[47:44]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_047 ,\cu_ru/al_ram_gpr_do_i1_046 ,\cu_ru/al_ram_gpr_do_i1_045 ,\cu_ru/al_ram_gpr_do_i1_044 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c12  (
    .di(data_rd[51:48]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_051 ,\cu_ru/al_ram_gpr_do_i1_050 ,\cu_ru/al_ram_gpr_do_i1_049 ,\cu_ru/al_ram_gpr_do_i1_048 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c13  (
    .di(data_rd[55:52]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_055 ,\cu_ru/al_ram_gpr_do_i1_054 ,\cu_ru/al_ram_gpr_do_i1_053 ,\cu_ru/al_ram_gpr_do_i1_052 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c14  (
    .di(data_rd[59:56]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_059 ,\cu_ru/al_ram_gpr_do_i1_058 ,\cu_ru/al_ram_gpr_do_i1_057 ,\cu_ru/al_ram_gpr_do_i1_056 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c15  (
    .di(data_rd[63:60]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_063 ,\cu_ru/al_ram_gpr_do_i1_062 ,\cu_ru/al_ram_gpr_do_i1_061 ,\cu_ru/al_ram_gpr_do_i1_060 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c2  (
    .di(data_rd[11:8]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_011 ,\cu_ru/al_ram_gpr_do_i1_010 ,\cu_ru/al_ram_gpr_do_i1_009 ,\cu_ru/al_ram_gpr_do_i1_008 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c3  (
    .di(data_rd[15:12]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_015 ,\cu_ru/al_ram_gpr_do_i1_014 ,\cu_ru/al_ram_gpr_do_i1_013 ,\cu_ru/al_ram_gpr_do_i1_012 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c4  (
    .di(data_rd[19:16]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_019 ,\cu_ru/al_ram_gpr_do_i1_018 ,\cu_ru/al_ram_gpr_do_i1_017 ,\cu_ru/al_ram_gpr_do_i1_016 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c5  (
    .di(data_rd[23:20]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_023 ,\cu_ru/al_ram_gpr_do_i1_022 ,\cu_ru/al_ram_gpr_do_i1_021 ,\cu_ru/al_ram_gpr_do_i1_020 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c6  (
    .di(data_rd[27:24]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_027 ,\cu_ru/al_ram_gpr_do_i1_026 ,\cu_ru/al_ram_gpr_do_i1_025 ,\cu_ru/al_ram_gpr_do_i1_024 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c7  (
    .di(data_rd[31:28]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_031 ,\cu_ru/al_ram_gpr_do_i1_030 ,\cu_ru/al_ram_gpr_do_i1_029 ,\cu_ru/al_ram_gpr_do_i1_028 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c8  (
    .di(data_rd[35:32]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_035 ,\cu_ru/al_ram_gpr_do_i1_034 ,\cu_ru/al_ram_gpr_do_i1_033 ,\cu_ru/al_ram_gpr_do_i1_032 }));
  EG_LOGIC_DRAM16X4 \cu_ru/al_ram_gpr_r1_c9  (
    .di(data_rd[39:36]),
    .raddr(\cu_ru/n46 [3:0]),
    .waddr(\cu_ru/n52 [3:0]),
    .wclk(clk_pad),
    .we(\cu_ru/n53_1_al_n1986 ),
    .do({\cu_ru/al_ram_gpr_do_i1_039 ,\cu_ru/al_ram_gpr_do_i1_038 ,\cu_ru/al_ram_gpr_do_i1_037 ,\cu_ru/al_ram_gpr_do_i1_036 }));
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b0  (
    .clk(clk_pad),
    .d(data_csr[0]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[0]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b1  (
    .clk(clk_pad),
    .d(data_csr[1]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[1]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b10  (
    .clk(clk_pad),
    .d(data_csr[10]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[10]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b11  (
    .clk(clk_pad),
    .d(data_csr[11]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[11]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b12  (
    .clk(clk_pad),
    .d(data_csr[12]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[12]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b13  (
    .clk(clk_pad),
    .d(data_csr[13]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[13]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b14  (
    .clk(clk_pad),
    .d(data_csr[14]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[14]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b15  (
    .clk(clk_pad),
    .d(data_csr[15]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[15]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b16  (
    .clk(clk_pad),
    .d(data_csr[16]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[16]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b17  (
    .clk(clk_pad),
    .d(data_csr[17]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[17]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b18  (
    .clk(clk_pad),
    .d(data_csr[18]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[18]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b19  (
    .clk(clk_pad),
    .d(data_csr[19]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[19]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b2  (
    .clk(clk_pad),
    .d(data_csr[2]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[2]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b20  (
    .clk(clk_pad),
    .d(data_csr[20]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[20]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b21  (
    .clk(clk_pad),
    .d(data_csr[21]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[21]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b22  (
    .clk(clk_pad),
    .d(data_csr[22]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[22]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b23  (
    .clk(clk_pad),
    .d(data_csr[23]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[23]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b24  (
    .clk(clk_pad),
    .d(data_csr[24]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[24]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b25  (
    .clk(clk_pad),
    .d(data_csr[25]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[25]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b26  (
    .clk(clk_pad),
    .d(data_csr[26]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[26]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b27  (
    .clk(clk_pad),
    .d(data_csr[27]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[27]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b28  (
    .clk(clk_pad),
    .d(data_csr[28]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[28]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b29  (
    .clk(clk_pad),
    .d(data_csr[29]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[29]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b3  (
    .clk(clk_pad),
    .d(data_csr[3]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[3]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b30  (
    .clk(clk_pad),
    .d(data_csr[30]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[30]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b31  (
    .clk(clk_pad),
    .d(data_csr[31]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[31]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b32  (
    .clk(clk_pad),
    .d(data_csr[32]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[32]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b33  (
    .clk(clk_pad),
    .d(data_csr[33]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[33]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b34  (
    .clk(clk_pad),
    .d(data_csr[34]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[34]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b35  (
    .clk(clk_pad),
    .d(data_csr[35]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[35]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b36  (
    .clk(clk_pad),
    .d(data_csr[36]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[36]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b37  (
    .clk(clk_pad),
    .d(data_csr[37]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[37]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b38  (
    .clk(clk_pad),
    .d(data_csr[38]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[38]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b39  (
    .clk(clk_pad),
    .d(data_csr[39]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[39]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b4  (
    .clk(clk_pad),
    .d(data_csr[4]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[4]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b40  (
    .clk(clk_pad),
    .d(data_csr[40]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[40]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b41  (
    .clk(clk_pad),
    .d(data_csr[41]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[41]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b42  (
    .clk(clk_pad),
    .d(data_csr[42]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[42]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b43  (
    .clk(clk_pad),
    .d(data_csr[43]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[43]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b5  (
    .clk(clk_pad),
    .d(data_csr[5]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[5]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b6  (
    .clk(clk_pad),
    .d(data_csr[6]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[6]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b7  (
    .clk(clk_pad),
    .d(data_csr[7]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[7]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b8  (
    .clk(clk_pad),
    .d(data_csr[8]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[8]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b9  (
    .clk(clk_pad),
    .d(data_csr[9]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[9]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg1_b0  (
    .clk(clk_pad),
    .d(data_csr[60]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[60]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg1_b1  (
    .clk(clk_pad),
    .d(data_csr[61]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[61]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg1_b2  (
    .clk(clk_pad),
    .d(data_csr[62]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[62]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg1_b3  (
    .clk(clk_pad),
    .d(data_csr[63]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(satp[63]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u0  (
    .a(\cu_ru/mcycle [0]),
    .b(1'b1),
    .c(\cu_ru/m_cycle_event/add0/c0 ),
    .o({\cu_ru/m_cycle_event/add0/c1 ,\cu_ru/m_cycle_event/n2 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u1  (
    .a(\cu_ru/mcycle [1]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c1 ),
    .o({\cu_ru/m_cycle_event/add0/c2 ,\cu_ru/m_cycle_event/n2 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u10  (
    .a(\cu_ru/mcycle [10]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c10 ),
    .o({\cu_ru/m_cycle_event/add0/c11 ,\cu_ru/m_cycle_event/n2 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u11  (
    .a(\cu_ru/mcycle [11]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c11 ),
    .o({\cu_ru/m_cycle_event/add0/c12 ,\cu_ru/m_cycle_event/n2 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u12  (
    .a(\cu_ru/mcycle [12]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c12 ),
    .o({\cu_ru/m_cycle_event/add0/c13 ,\cu_ru/m_cycle_event/n2 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u13  (
    .a(\cu_ru/mcycle [13]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c13 ),
    .o({\cu_ru/m_cycle_event/add0/c14 ,\cu_ru/m_cycle_event/n2 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u14  (
    .a(\cu_ru/mcycle [14]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c14 ),
    .o({\cu_ru/m_cycle_event/add0/c15 ,\cu_ru/m_cycle_event/n2 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u15  (
    .a(\cu_ru/mcycle [15]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c15 ),
    .o({\cu_ru/m_cycle_event/add0/c16 ,\cu_ru/m_cycle_event/n2 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u16  (
    .a(\cu_ru/mcycle [16]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c16 ),
    .o({\cu_ru/m_cycle_event/add0/c17 ,\cu_ru/m_cycle_event/n2 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u17  (
    .a(\cu_ru/mcycle [17]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c17 ),
    .o({\cu_ru/m_cycle_event/add0/c18 ,\cu_ru/m_cycle_event/n2 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u18  (
    .a(\cu_ru/mcycle [18]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c18 ),
    .o({\cu_ru/m_cycle_event/add0/c19 ,\cu_ru/m_cycle_event/n2 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u19  (
    .a(\cu_ru/mcycle [19]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c19 ),
    .o({\cu_ru/m_cycle_event/add0/c20 ,\cu_ru/m_cycle_event/n2 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u2  (
    .a(\cu_ru/mcycle [2]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c2 ),
    .o({\cu_ru/m_cycle_event/add0/c3 ,\cu_ru/m_cycle_event/n2 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u20  (
    .a(\cu_ru/mcycle [20]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c20 ),
    .o({\cu_ru/m_cycle_event/add0/c21 ,\cu_ru/m_cycle_event/n2 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u21  (
    .a(\cu_ru/mcycle [21]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c21 ),
    .o({\cu_ru/m_cycle_event/add0/c22 ,\cu_ru/m_cycle_event/n2 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u22  (
    .a(\cu_ru/mcycle [22]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c22 ),
    .o({\cu_ru/m_cycle_event/add0/c23 ,\cu_ru/m_cycle_event/n2 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u23  (
    .a(\cu_ru/mcycle [23]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c23 ),
    .o({\cu_ru/m_cycle_event/add0/c24 ,\cu_ru/m_cycle_event/n2 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u24  (
    .a(\cu_ru/mcycle [24]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c24 ),
    .o({\cu_ru/m_cycle_event/add0/c25 ,\cu_ru/m_cycle_event/n2 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u25  (
    .a(\cu_ru/mcycle [25]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c25 ),
    .o({\cu_ru/m_cycle_event/add0/c26 ,\cu_ru/m_cycle_event/n2 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u26  (
    .a(\cu_ru/mcycle [26]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c26 ),
    .o({\cu_ru/m_cycle_event/add0/c27 ,\cu_ru/m_cycle_event/n2 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u27  (
    .a(\cu_ru/mcycle [27]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c27 ),
    .o({\cu_ru/m_cycle_event/add0/c28 ,\cu_ru/m_cycle_event/n2 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u28  (
    .a(\cu_ru/mcycle [28]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c28 ),
    .o({\cu_ru/m_cycle_event/add0/c29 ,\cu_ru/m_cycle_event/n2 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u29  (
    .a(\cu_ru/mcycle [29]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c29 ),
    .o({\cu_ru/m_cycle_event/add0/c30 ,\cu_ru/m_cycle_event/n2 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u3  (
    .a(\cu_ru/mcycle [3]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c3 ),
    .o({\cu_ru/m_cycle_event/add0/c4 ,\cu_ru/m_cycle_event/n2 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u30  (
    .a(\cu_ru/mcycle [30]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c30 ),
    .o({\cu_ru/m_cycle_event/add0/c31 ,\cu_ru/m_cycle_event/n2 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u31  (
    .a(\cu_ru/mcycle [31]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c31 ),
    .o({\cu_ru/m_cycle_event/add0/c32 ,\cu_ru/m_cycle_event/n2 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u32  (
    .a(\cu_ru/mcycle [32]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c32 ),
    .o({\cu_ru/m_cycle_event/add0/c33 ,\cu_ru/m_cycle_event/n2 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u33  (
    .a(\cu_ru/mcycle [33]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c33 ),
    .o({\cu_ru/m_cycle_event/add0/c34 ,\cu_ru/m_cycle_event/n2 [33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u34  (
    .a(\cu_ru/mcycle [34]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c34 ),
    .o({\cu_ru/m_cycle_event/add0/c35 ,\cu_ru/m_cycle_event/n2 [34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u35  (
    .a(\cu_ru/mcycle [35]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c35 ),
    .o({\cu_ru/m_cycle_event/add0/c36 ,\cu_ru/m_cycle_event/n2 [35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u36  (
    .a(\cu_ru/mcycle [36]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c36 ),
    .o({\cu_ru/m_cycle_event/add0/c37 ,\cu_ru/m_cycle_event/n2 [36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u37  (
    .a(\cu_ru/mcycle [37]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c37 ),
    .o({\cu_ru/m_cycle_event/add0/c38 ,\cu_ru/m_cycle_event/n2 [37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u38  (
    .a(\cu_ru/mcycle [38]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c38 ),
    .o({\cu_ru/m_cycle_event/add0/c39 ,\cu_ru/m_cycle_event/n2 [38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u39  (
    .a(\cu_ru/mcycle [39]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c39 ),
    .o({\cu_ru/m_cycle_event/add0/c40 ,\cu_ru/m_cycle_event/n2 [39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u4  (
    .a(\cu_ru/mcycle [4]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c4 ),
    .o({\cu_ru/m_cycle_event/add0/c5 ,\cu_ru/m_cycle_event/n2 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u40  (
    .a(\cu_ru/mcycle [40]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c40 ),
    .o({\cu_ru/m_cycle_event/add0/c41 ,\cu_ru/m_cycle_event/n2 [40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u41  (
    .a(\cu_ru/mcycle [41]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c41 ),
    .o({\cu_ru/m_cycle_event/add0/c42 ,\cu_ru/m_cycle_event/n2 [41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u42  (
    .a(\cu_ru/mcycle [42]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c42 ),
    .o({\cu_ru/m_cycle_event/add0/c43 ,\cu_ru/m_cycle_event/n2 [42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u43  (
    .a(\cu_ru/mcycle [43]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c43 ),
    .o({\cu_ru/m_cycle_event/add0/c44 ,\cu_ru/m_cycle_event/n2 [43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u44  (
    .a(\cu_ru/mcycle [44]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c44 ),
    .o({\cu_ru/m_cycle_event/add0/c45 ,\cu_ru/m_cycle_event/n2 [44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u45  (
    .a(\cu_ru/mcycle [45]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c45 ),
    .o({\cu_ru/m_cycle_event/add0/c46 ,\cu_ru/m_cycle_event/n2 [45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u46  (
    .a(\cu_ru/mcycle [46]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c46 ),
    .o({\cu_ru/m_cycle_event/add0/c47 ,\cu_ru/m_cycle_event/n2 [46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u47  (
    .a(\cu_ru/mcycle [47]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c47 ),
    .o({\cu_ru/m_cycle_event/add0/c48 ,\cu_ru/m_cycle_event/n2 [47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u48  (
    .a(\cu_ru/mcycle [48]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c48 ),
    .o({\cu_ru/m_cycle_event/add0/c49 ,\cu_ru/m_cycle_event/n2 [48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u49  (
    .a(\cu_ru/mcycle [49]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c49 ),
    .o({\cu_ru/m_cycle_event/add0/c50 ,\cu_ru/m_cycle_event/n2 [49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u5  (
    .a(\cu_ru/mcycle [5]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c5 ),
    .o({\cu_ru/m_cycle_event/add0/c6 ,\cu_ru/m_cycle_event/n2 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u50  (
    .a(\cu_ru/mcycle [50]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c50 ),
    .o({\cu_ru/m_cycle_event/add0/c51 ,\cu_ru/m_cycle_event/n2 [50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u51  (
    .a(\cu_ru/mcycle [51]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c51 ),
    .o({\cu_ru/m_cycle_event/add0/c52 ,\cu_ru/m_cycle_event/n2 [51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u52  (
    .a(\cu_ru/mcycle [52]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c52 ),
    .o({\cu_ru/m_cycle_event/add0/c53 ,\cu_ru/m_cycle_event/n2 [52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u53  (
    .a(\cu_ru/mcycle [53]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c53 ),
    .o({\cu_ru/m_cycle_event/add0/c54 ,\cu_ru/m_cycle_event/n2 [53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u54  (
    .a(\cu_ru/mcycle [54]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c54 ),
    .o({\cu_ru/m_cycle_event/add0/c55 ,\cu_ru/m_cycle_event/n2 [54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u55  (
    .a(\cu_ru/mcycle [55]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c55 ),
    .o({\cu_ru/m_cycle_event/add0/c56 ,\cu_ru/m_cycle_event/n2 [55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u56  (
    .a(\cu_ru/mcycle [56]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c56 ),
    .o({\cu_ru/m_cycle_event/add0/c57 ,\cu_ru/m_cycle_event/n2 [56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u57  (
    .a(\cu_ru/mcycle [57]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c57 ),
    .o({\cu_ru/m_cycle_event/add0/c58 ,\cu_ru/m_cycle_event/n2 [57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u58  (
    .a(\cu_ru/mcycle [58]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c58 ),
    .o({\cu_ru/m_cycle_event/add0/c59 ,\cu_ru/m_cycle_event/n2 [58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u59  (
    .a(\cu_ru/mcycle [59]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c59 ),
    .o({\cu_ru/m_cycle_event/add0/c60 ,\cu_ru/m_cycle_event/n2 [59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u6  (
    .a(\cu_ru/mcycle [6]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c6 ),
    .o({\cu_ru/m_cycle_event/add0/c7 ,\cu_ru/m_cycle_event/n2 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u60  (
    .a(\cu_ru/mcycle [60]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c60 ),
    .o({\cu_ru/m_cycle_event/add0/c61 ,\cu_ru/m_cycle_event/n2 [60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u61  (
    .a(\cu_ru/mcycle [61]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c61 ),
    .o({\cu_ru/m_cycle_event/add0/c62 ,\cu_ru/m_cycle_event/n2 [61]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u62  (
    .a(\cu_ru/mcycle [62]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c62 ),
    .o({\cu_ru/m_cycle_event/add0/c63 ,\cu_ru/m_cycle_event/n2 [62]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u63  (
    .a(\cu_ru/mcycle [63]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c63 ),
    .o({open_n6066,\cu_ru/m_cycle_event/n2 [63]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u7  (
    .a(\cu_ru/mcycle [7]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c7 ),
    .o({\cu_ru/m_cycle_event/add0/c8 ,\cu_ru/m_cycle_event/n2 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u8  (
    .a(\cu_ru/mcycle [8]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c8 ),
    .o({\cu_ru/m_cycle_event/add0/c9 ,\cu_ru/m_cycle_event/n2 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add0/u9  (
    .a(\cu_ru/mcycle [9]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add0/c9 ),
    .o({\cu_ru/m_cycle_event/add0/c10 ,\cu_ru/m_cycle_event/n2 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \cu_ru/m_cycle_event/add0/ucin  (
    .a(1'b0),
    .o({\cu_ru/m_cycle_event/add0/c0 ,open_n6069}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u0  (
    .a(\cu_ru/minstret [0]),
    .b(1'b1),
    .c(\cu_ru/m_cycle_event/add1/c0 ),
    .o({\cu_ru/m_cycle_event/add1/c1 ,\cu_ru/m_cycle_event/n4 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u1  (
    .a(\cu_ru/minstret [1]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c1 ),
    .o({\cu_ru/m_cycle_event/add1/c2 ,\cu_ru/m_cycle_event/n4 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u10  (
    .a(\cu_ru/minstret [10]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c10 ),
    .o({\cu_ru/m_cycle_event/add1/c11 ,\cu_ru/m_cycle_event/n4 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u11  (
    .a(\cu_ru/minstret [11]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c11 ),
    .o({\cu_ru/m_cycle_event/add1/c12 ,\cu_ru/m_cycle_event/n4 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u12  (
    .a(\cu_ru/minstret [12]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c12 ),
    .o({\cu_ru/m_cycle_event/add1/c13 ,\cu_ru/m_cycle_event/n4 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u13  (
    .a(\cu_ru/minstret [13]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c13 ),
    .o({\cu_ru/m_cycle_event/add1/c14 ,\cu_ru/m_cycle_event/n4 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u14  (
    .a(\cu_ru/minstret [14]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c14 ),
    .o({\cu_ru/m_cycle_event/add1/c15 ,\cu_ru/m_cycle_event/n4 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u15  (
    .a(\cu_ru/minstret [15]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c15 ),
    .o({\cu_ru/m_cycle_event/add1/c16 ,\cu_ru/m_cycle_event/n4 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u16  (
    .a(\cu_ru/minstret [16]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c16 ),
    .o({\cu_ru/m_cycle_event/add1/c17 ,\cu_ru/m_cycle_event/n4 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u17  (
    .a(\cu_ru/minstret [17]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c17 ),
    .o({\cu_ru/m_cycle_event/add1/c18 ,\cu_ru/m_cycle_event/n4 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u18  (
    .a(\cu_ru/minstret [18]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c18 ),
    .o({\cu_ru/m_cycle_event/add1/c19 ,\cu_ru/m_cycle_event/n4 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u19  (
    .a(\cu_ru/minstret [19]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c19 ),
    .o({\cu_ru/m_cycle_event/add1/c20 ,\cu_ru/m_cycle_event/n4 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u2  (
    .a(\cu_ru/minstret [2]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c2 ),
    .o({\cu_ru/m_cycle_event/add1/c3 ,\cu_ru/m_cycle_event/n4 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u20  (
    .a(\cu_ru/minstret [20]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c20 ),
    .o({\cu_ru/m_cycle_event/add1/c21 ,\cu_ru/m_cycle_event/n4 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u21  (
    .a(\cu_ru/minstret [21]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c21 ),
    .o({\cu_ru/m_cycle_event/add1/c22 ,\cu_ru/m_cycle_event/n4 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u22  (
    .a(\cu_ru/minstret [22]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c22 ),
    .o({\cu_ru/m_cycle_event/add1/c23 ,\cu_ru/m_cycle_event/n4 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u23  (
    .a(\cu_ru/minstret [23]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c23 ),
    .o({\cu_ru/m_cycle_event/add1/c24 ,\cu_ru/m_cycle_event/n4 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u24  (
    .a(\cu_ru/minstret [24]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c24 ),
    .o({\cu_ru/m_cycle_event/add1/c25 ,\cu_ru/m_cycle_event/n4 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u25  (
    .a(\cu_ru/minstret [25]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c25 ),
    .o({\cu_ru/m_cycle_event/add1/c26 ,\cu_ru/m_cycle_event/n4 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u26  (
    .a(\cu_ru/minstret [26]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c26 ),
    .o({\cu_ru/m_cycle_event/add1/c27 ,\cu_ru/m_cycle_event/n4 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u27  (
    .a(\cu_ru/minstret [27]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c27 ),
    .o({\cu_ru/m_cycle_event/add1/c28 ,\cu_ru/m_cycle_event/n4 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u28  (
    .a(\cu_ru/minstret [28]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c28 ),
    .o({\cu_ru/m_cycle_event/add1/c29 ,\cu_ru/m_cycle_event/n4 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u29  (
    .a(\cu_ru/minstret [29]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c29 ),
    .o({\cu_ru/m_cycle_event/add1/c30 ,\cu_ru/m_cycle_event/n4 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u3  (
    .a(\cu_ru/minstret [3]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c3 ),
    .o({\cu_ru/m_cycle_event/add1/c4 ,\cu_ru/m_cycle_event/n4 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u30  (
    .a(\cu_ru/minstret [30]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c30 ),
    .o({\cu_ru/m_cycle_event/add1/c31 ,\cu_ru/m_cycle_event/n4 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u31  (
    .a(\cu_ru/minstret [31]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c31 ),
    .o({\cu_ru/m_cycle_event/add1/c32 ,\cu_ru/m_cycle_event/n4 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u32  (
    .a(\cu_ru/minstret [32]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c32 ),
    .o({\cu_ru/m_cycle_event/add1/c33 ,\cu_ru/m_cycle_event/n4 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u33  (
    .a(\cu_ru/minstret [33]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c33 ),
    .o({\cu_ru/m_cycle_event/add1/c34 ,\cu_ru/m_cycle_event/n4 [33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u34  (
    .a(\cu_ru/minstret [34]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c34 ),
    .o({\cu_ru/m_cycle_event/add1/c35 ,\cu_ru/m_cycle_event/n4 [34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u35  (
    .a(\cu_ru/minstret [35]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c35 ),
    .o({\cu_ru/m_cycle_event/add1/c36 ,\cu_ru/m_cycle_event/n4 [35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u36  (
    .a(\cu_ru/minstret [36]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c36 ),
    .o({\cu_ru/m_cycle_event/add1/c37 ,\cu_ru/m_cycle_event/n4 [36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u37  (
    .a(\cu_ru/minstret [37]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c37 ),
    .o({\cu_ru/m_cycle_event/add1/c38 ,\cu_ru/m_cycle_event/n4 [37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u38  (
    .a(\cu_ru/minstret [38]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c38 ),
    .o({\cu_ru/m_cycle_event/add1/c39 ,\cu_ru/m_cycle_event/n4 [38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u39  (
    .a(\cu_ru/minstret [39]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c39 ),
    .o({\cu_ru/m_cycle_event/add1/c40 ,\cu_ru/m_cycle_event/n4 [39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u4  (
    .a(\cu_ru/minstret [4]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c4 ),
    .o({\cu_ru/m_cycle_event/add1/c5 ,\cu_ru/m_cycle_event/n4 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u40  (
    .a(\cu_ru/minstret [40]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c40 ),
    .o({\cu_ru/m_cycle_event/add1/c41 ,\cu_ru/m_cycle_event/n4 [40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u41  (
    .a(\cu_ru/minstret [41]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c41 ),
    .o({\cu_ru/m_cycle_event/add1/c42 ,\cu_ru/m_cycle_event/n4 [41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u42  (
    .a(\cu_ru/minstret [42]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c42 ),
    .o({\cu_ru/m_cycle_event/add1/c43 ,\cu_ru/m_cycle_event/n4 [42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u43  (
    .a(\cu_ru/minstret [43]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c43 ),
    .o({\cu_ru/m_cycle_event/add1/c44 ,\cu_ru/m_cycle_event/n4 [43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u44  (
    .a(\cu_ru/minstret [44]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c44 ),
    .o({\cu_ru/m_cycle_event/add1/c45 ,\cu_ru/m_cycle_event/n4 [44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u45  (
    .a(\cu_ru/minstret [45]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c45 ),
    .o({\cu_ru/m_cycle_event/add1/c46 ,\cu_ru/m_cycle_event/n4 [45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u46  (
    .a(\cu_ru/minstret [46]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c46 ),
    .o({\cu_ru/m_cycle_event/add1/c47 ,\cu_ru/m_cycle_event/n4 [46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u47  (
    .a(\cu_ru/minstret [47]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c47 ),
    .o({\cu_ru/m_cycle_event/add1/c48 ,\cu_ru/m_cycle_event/n4 [47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u48  (
    .a(\cu_ru/minstret [48]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c48 ),
    .o({\cu_ru/m_cycle_event/add1/c49 ,\cu_ru/m_cycle_event/n4 [48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u49  (
    .a(\cu_ru/minstret [49]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c49 ),
    .o({\cu_ru/m_cycle_event/add1/c50 ,\cu_ru/m_cycle_event/n4 [49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u5  (
    .a(\cu_ru/minstret [5]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c5 ),
    .o({\cu_ru/m_cycle_event/add1/c6 ,\cu_ru/m_cycle_event/n4 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u50  (
    .a(\cu_ru/minstret [50]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c50 ),
    .o({\cu_ru/m_cycle_event/add1/c51 ,\cu_ru/m_cycle_event/n4 [50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u51  (
    .a(\cu_ru/minstret [51]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c51 ),
    .o({\cu_ru/m_cycle_event/add1/c52 ,\cu_ru/m_cycle_event/n4 [51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u52  (
    .a(\cu_ru/minstret [52]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c52 ),
    .o({\cu_ru/m_cycle_event/add1/c53 ,\cu_ru/m_cycle_event/n4 [52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u53  (
    .a(\cu_ru/minstret [53]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c53 ),
    .o({\cu_ru/m_cycle_event/add1/c54 ,\cu_ru/m_cycle_event/n4 [53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u54  (
    .a(\cu_ru/minstret [54]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c54 ),
    .o({\cu_ru/m_cycle_event/add1/c55 ,\cu_ru/m_cycle_event/n4 [54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u55  (
    .a(\cu_ru/minstret [55]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c55 ),
    .o({\cu_ru/m_cycle_event/add1/c56 ,\cu_ru/m_cycle_event/n4 [55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u56  (
    .a(\cu_ru/minstret [56]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c56 ),
    .o({\cu_ru/m_cycle_event/add1/c57 ,\cu_ru/m_cycle_event/n4 [56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u57  (
    .a(\cu_ru/minstret [57]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c57 ),
    .o({\cu_ru/m_cycle_event/add1/c58 ,\cu_ru/m_cycle_event/n4 [57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u58  (
    .a(\cu_ru/minstret [58]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c58 ),
    .o({\cu_ru/m_cycle_event/add1/c59 ,\cu_ru/m_cycle_event/n4 [58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u59  (
    .a(\cu_ru/minstret [59]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c59 ),
    .o({\cu_ru/m_cycle_event/add1/c60 ,\cu_ru/m_cycle_event/n4 [59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u6  (
    .a(\cu_ru/minstret [6]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c6 ),
    .o({\cu_ru/m_cycle_event/add1/c7 ,\cu_ru/m_cycle_event/n4 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u60  (
    .a(\cu_ru/minstret [60]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c60 ),
    .o({\cu_ru/m_cycle_event/add1/c61 ,\cu_ru/m_cycle_event/n4 [60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u61  (
    .a(\cu_ru/minstret [61]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c61 ),
    .o({\cu_ru/m_cycle_event/add1/c62 ,\cu_ru/m_cycle_event/n4 [61]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u62  (
    .a(\cu_ru/minstret [62]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c62 ),
    .o({\cu_ru/m_cycle_event/add1/c63 ,\cu_ru/m_cycle_event/n4 [62]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u63  (
    .a(\cu_ru/minstret [63]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c63 ),
    .o({open_n6070,\cu_ru/m_cycle_event/n4 [63]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u7  (
    .a(\cu_ru/minstret [7]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c7 ),
    .o({\cu_ru/m_cycle_event/add1/c8 ,\cu_ru/m_cycle_event/n4 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u8  (
    .a(\cu_ru/minstret [8]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c8 ),
    .o({\cu_ru/m_cycle_event/add1/c9 ,\cu_ru/m_cycle_event/n4 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_cycle_event/add1/u9  (
    .a(\cu_ru/minstret [9]),
    .b(1'b0),
    .c(\cu_ru/m_cycle_event/add1/c9 ),
    .o({\cu_ru/m_cycle_event/add1/c10 ,\cu_ru/m_cycle_event/n4 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \cu_ru/m_cycle_event/add1/ucin  (
    .a(1'b0),
    .o({\cu_ru/m_cycle_event/add1/c0 ,open_n6073}));
  reg_sr_as_w1 \cu_ru/m_cycle_event/cy_reg  (
    .clk(clk_pad),
    .d(data_csr[0]),
    .en(\cu_ru/m_cycle_event/n13 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcountinhibit ));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(51)
  reg_sr_as_w1 \cu_ru/m_cycle_event/ir_reg  (
    .clk(clk_pad),
    .d(data_csr[2]),
    .en(\cu_ru/m_cycle_event/n13 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/m_cycle_event/mcountinhibit[2] ));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(51)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b0  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [0]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [0]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b1  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [1]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [1]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b10  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [10]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [10]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b11  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [11]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [11]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b12  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [12]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [12]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b13  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [13]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [13]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b14  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [14]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [14]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b15  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [15]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [15]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b16  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [16]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [16]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b17  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [17]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [17]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b18  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [18]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [18]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b19  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [19]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [19]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b2  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [2]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [2]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b20  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [20]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [20]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b21  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [21]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [21]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b22  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [22]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [22]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b23  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [23]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [23]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b24  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [24]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [24]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b25  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [25]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [25]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b26  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [26]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [26]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b27  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [27]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [27]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b28  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [28]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [28]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b29  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [29]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [29]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b3  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [3]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [3]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b30  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [30]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [30]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b31  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [31]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [31]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b32  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [32]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [32]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b33  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [33]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [33]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b34  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [34]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [34]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b35  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [35]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [35]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b36  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [36]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [36]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b37  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [37]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [37]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b38  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [38]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [38]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b39  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [39]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [39]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b4  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [4]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [4]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b40  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [40]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [40]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b41  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [41]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [41]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b42  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [42]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [42]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b43  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [43]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [43]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b44  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [44]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [44]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b45  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [45]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [45]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b46  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [46]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [46]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b47  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [47]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [47]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b48  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [48]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [48]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b49  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [49]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [49]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b5  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [5]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [5]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b50  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [50]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [50]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b51  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [51]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [51]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b52  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [52]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [52]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b53  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [53]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [53]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b54  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [54]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [54]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b55  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [55]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [55]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b56  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [56]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [56]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b57  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [57]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [57]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b58  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [58]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [58]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b59  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [59]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [59]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b6  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [6]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [6]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b60  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [60]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [60]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b61  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [61]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [61]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b62  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [62]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [62]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b63  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [63]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [63]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b7  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [7]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [7]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b8  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [8]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [8]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b9  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n4 [9]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/minstret [9]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b0  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [0]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b1  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [1]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b10  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [10]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b11  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [11]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b12  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [12]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b13  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [13]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b14  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [14]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b15  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [15]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b16  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [16]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b17  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [17]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b18  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [18]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b19  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [19]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b2  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [2]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b20  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [20]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b21  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [21]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b22  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [22]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b23  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [23]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b24  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [24]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b25  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [25]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b26  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [26]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b27  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [27]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b28  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [28]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b29  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [29]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b3  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [3]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b30  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [30]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b31  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [31]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b32  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [32]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b33  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [33]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b34  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [34]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b35  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [35]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b36  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [36]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b37  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [37]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b38  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [38]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b39  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [39]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b4  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [4]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b40  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [40]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b41  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [41]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b42  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [42]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b43  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [43]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b44  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [44]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b45  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [45]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b46  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [46]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b47  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [47]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b48  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [48]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b49  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [49]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b5  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [5]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b50  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [50]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b51  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [51]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b52  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [52]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b53  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [53]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b54  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [54]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b55  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [55]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b56  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [56]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b57  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [57]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b58  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [58]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b59  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [59]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b6  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [6]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b60  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [60]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b61  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [61]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b62  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [62]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b63  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [63]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b7  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [7]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b8  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [8]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b9  (
    .clk(clk_pad),
    .d(\cu_ru/m_cycle_event/n9 [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcycle [9]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b0  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [0]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b1  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [1]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b10  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [10]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b11  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [11]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b12  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [12]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b13  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [13]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b14  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [14]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b15  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [15]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b16  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [16]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b17  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [17]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b18  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [18]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b19  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [19]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b2  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [2]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b20  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [20]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b21  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [21]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b22  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [22]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b23  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [23]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b24  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [24]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b25  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [25]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b26  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [26]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b27  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [27]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b28  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [28]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b29  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [29]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b3  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [3]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b30  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [30]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b31  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [31]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b32  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [32]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b33  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [33]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b34  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [34]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b35  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [35]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b36  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [36]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b37  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [37]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b38  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [38]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b39  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [39]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b4  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [4]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b40  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [40]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b41  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [41]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b42  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [42]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b43  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [43]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b44  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [44]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b45  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [45]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b46  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [46]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b47  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [47]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b48  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [48]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b49  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [49]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b5  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [5]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b50  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [50]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b51  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [51]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b52  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [52]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b53  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [53]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b54  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [54]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b55  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [55]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b56  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [56]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b57  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [57]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b58  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [58]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b59  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [59]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b6  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [6]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b60  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [60]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b61  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [61]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b62  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [62]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b63  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [63]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b7  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [7]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b8  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [8]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b9  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n5 [9]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/scause [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b0  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n7 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcause [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b1  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n7 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcause [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b10  (
    .clk(clk_pad),
    .d(data_csr[10]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b11  (
    .clk(clk_pad),
    .d(data_csr[11]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b12  (
    .clk(clk_pad),
    .d(data_csr[12]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b13  (
    .clk(clk_pad),
    .d(data_csr[13]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b14  (
    .clk(clk_pad),
    .d(data_csr[14]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b15  (
    .clk(clk_pad),
    .d(data_csr[15]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b16  (
    .clk(clk_pad),
    .d(data_csr[16]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b17  (
    .clk(clk_pad),
    .d(data_csr[17]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b18  (
    .clk(clk_pad),
    .d(data_csr[18]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b19  (
    .clk(clk_pad),
    .d(data_csr[19]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b2  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n7 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcause [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b20  (
    .clk(clk_pad),
    .d(data_csr[20]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b21  (
    .clk(clk_pad),
    .d(data_csr[21]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b22  (
    .clk(clk_pad),
    .d(data_csr[22]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b23  (
    .clk(clk_pad),
    .d(data_csr[23]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b24  (
    .clk(clk_pad),
    .d(data_csr[24]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b25  (
    .clk(clk_pad),
    .d(data_csr[25]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b26  (
    .clk(clk_pad),
    .d(data_csr[26]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b27  (
    .clk(clk_pad),
    .d(data_csr[27]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b28  (
    .clk(clk_pad),
    .d(data_csr[28]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b29  (
    .clk(clk_pad),
    .d(data_csr[29]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b3  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n7 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcause [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b30  (
    .clk(clk_pad),
    .d(data_csr[30]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b31  (
    .clk(clk_pad),
    .d(data_csr[31]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b32  (
    .clk(clk_pad),
    .d(data_csr[32]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b33  (
    .clk(clk_pad),
    .d(data_csr[33]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b34  (
    .clk(clk_pad),
    .d(data_csr[34]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b35  (
    .clk(clk_pad),
    .d(data_csr[35]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b36  (
    .clk(clk_pad),
    .d(data_csr[36]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b37  (
    .clk(clk_pad),
    .d(data_csr[37]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b38  (
    .clk(clk_pad),
    .d(data_csr[38]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b39  (
    .clk(clk_pad),
    .d(data_csr[39]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b4  (
    .clk(clk_pad),
    .d(data_csr[4]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b40  (
    .clk(clk_pad),
    .d(data_csr[40]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b41  (
    .clk(clk_pad),
    .d(data_csr[41]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b42  (
    .clk(clk_pad),
    .d(data_csr[42]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b43  (
    .clk(clk_pad),
    .d(data_csr[43]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b44  (
    .clk(clk_pad),
    .d(data_csr[44]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b45  (
    .clk(clk_pad),
    .d(data_csr[45]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b46  (
    .clk(clk_pad),
    .d(data_csr[46]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b47  (
    .clk(clk_pad),
    .d(data_csr[47]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b48  (
    .clk(clk_pad),
    .d(data_csr[48]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b49  (
    .clk(clk_pad),
    .d(data_csr[49]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b5  (
    .clk(clk_pad),
    .d(data_csr[5]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b50  (
    .clk(clk_pad),
    .d(data_csr[50]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b51  (
    .clk(clk_pad),
    .d(data_csr[51]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b52  (
    .clk(clk_pad),
    .d(data_csr[52]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b53  (
    .clk(clk_pad),
    .d(data_csr[53]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b54  (
    .clk(clk_pad),
    .d(data_csr[54]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b55  (
    .clk(clk_pad),
    .d(data_csr[55]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b56  (
    .clk(clk_pad),
    .d(data_csr[56]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b57  (
    .clk(clk_pad),
    .d(data_csr[57]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b58  (
    .clk(clk_pad),
    .d(data_csr[58]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b59  (
    .clk(clk_pad),
    .d(data_csr[59]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b6  (
    .clk(clk_pad),
    .d(data_csr[6]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b60  (
    .clk(clk_pad),
    .d(data_csr[60]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b61  (
    .clk(clk_pad),
    .d(data_csr[61]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b62  (
    .clk(clk_pad),
    .d(data_csr[62]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b63  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_cause/n7 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mcause [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b7  (
    .clk(clk_pad),
    .d(data_csr[7]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b8  (
    .clk(clk_pad),
    .d(data_csr[8]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b9  (
    .clk(clk_pad),
    .d(data_csr[9]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u0  (
    .a(wb_ins_pc[2]),
    .b(1'b1),
    .c(\cu_ru/m_s_epc/add0/c0 ),
    .o({\cu_ru/m_s_epc/add0/c1 ,\cu_ru/m_s_epc/n0 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u1  (
    .a(wb_ins_pc[3]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c1 ),
    .o({\cu_ru/m_s_epc/add0/c2 ,\cu_ru/m_s_epc/n0 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u10  (
    .a(wb_ins_pc[12]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c10 ),
    .o({\cu_ru/m_s_epc/add0/c11 ,\cu_ru/m_s_epc/n0 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u11  (
    .a(wb_ins_pc[13]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c11 ),
    .o({\cu_ru/m_s_epc/add0/c12 ,\cu_ru/m_s_epc/n0 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u12  (
    .a(wb_ins_pc[14]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c12 ),
    .o({\cu_ru/m_s_epc/add0/c13 ,\cu_ru/m_s_epc/n0 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u13  (
    .a(wb_ins_pc[15]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c13 ),
    .o({\cu_ru/m_s_epc/add0/c14 ,\cu_ru/m_s_epc/n0 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u14  (
    .a(wb_ins_pc[16]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c14 ),
    .o({\cu_ru/m_s_epc/add0/c15 ,\cu_ru/m_s_epc/n0 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u15  (
    .a(wb_ins_pc[17]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c15 ),
    .o({\cu_ru/m_s_epc/add0/c16 ,\cu_ru/m_s_epc/n0 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u16  (
    .a(wb_ins_pc[18]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c16 ),
    .o({\cu_ru/m_s_epc/add0/c17 ,\cu_ru/m_s_epc/n0 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u17  (
    .a(wb_ins_pc[19]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c17 ),
    .o({\cu_ru/m_s_epc/add0/c18 ,\cu_ru/m_s_epc/n0 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u18  (
    .a(wb_ins_pc[20]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c18 ),
    .o({\cu_ru/m_s_epc/add0/c19 ,\cu_ru/m_s_epc/n0 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u19  (
    .a(wb_ins_pc[21]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c19 ),
    .o({\cu_ru/m_s_epc/add0/c20 ,\cu_ru/m_s_epc/n0 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u2  (
    .a(wb_ins_pc[4]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c2 ),
    .o({\cu_ru/m_s_epc/add0/c3 ,\cu_ru/m_s_epc/n0 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u20  (
    .a(wb_ins_pc[22]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c20 ),
    .o({\cu_ru/m_s_epc/add0/c21 ,\cu_ru/m_s_epc/n0 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u21  (
    .a(wb_ins_pc[23]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c21 ),
    .o({\cu_ru/m_s_epc/add0/c22 ,\cu_ru/m_s_epc/n0 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u22  (
    .a(wb_ins_pc[24]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c22 ),
    .o({\cu_ru/m_s_epc/add0/c23 ,\cu_ru/m_s_epc/n0 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u23  (
    .a(wb_ins_pc[25]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c23 ),
    .o({\cu_ru/m_s_epc/add0/c24 ,\cu_ru/m_s_epc/n0 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u24  (
    .a(wb_ins_pc[26]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c24 ),
    .o({\cu_ru/m_s_epc/add0/c25 ,\cu_ru/m_s_epc/n0 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u25  (
    .a(wb_ins_pc[27]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c25 ),
    .o({\cu_ru/m_s_epc/add0/c26 ,\cu_ru/m_s_epc/n0 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u26  (
    .a(wb_ins_pc[28]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c26 ),
    .o({\cu_ru/m_s_epc/add0/c27 ,\cu_ru/m_s_epc/n0 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u27  (
    .a(wb_ins_pc[29]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c27 ),
    .o({\cu_ru/m_s_epc/add0/c28 ,\cu_ru/m_s_epc/n0 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u28  (
    .a(wb_ins_pc[30]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c28 ),
    .o({\cu_ru/m_s_epc/add0/c29 ,\cu_ru/m_s_epc/n0 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u29  (
    .a(wb_ins_pc[31]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c29 ),
    .o({\cu_ru/m_s_epc/add0/c30 ,\cu_ru/m_s_epc/n0 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u3  (
    .a(wb_ins_pc[5]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c3 ),
    .o({\cu_ru/m_s_epc/add0/c4 ,\cu_ru/m_s_epc/n0 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u30  (
    .a(wb_ins_pc[32]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c30 ),
    .o({\cu_ru/m_s_epc/add0/c31 ,\cu_ru/m_s_epc/n0 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u31  (
    .a(wb_ins_pc[33]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c31 ),
    .o({\cu_ru/m_s_epc/add0/c32 ,\cu_ru/m_s_epc/n0 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u32  (
    .a(wb_ins_pc[34]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c32 ),
    .o({\cu_ru/m_s_epc/add0/c33 ,\cu_ru/m_s_epc/n0 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u33  (
    .a(wb_ins_pc[35]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c33 ),
    .o({\cu_ru/m_s_epc/add0/c34 ,\cu_ru/m_s_epc/n0 [33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u34  (
    .a(wb_ins_pc[36]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c34 ),
    .o({\cu_ru/m_s_epc/add0/c35 ,\cu_ru/m_s_epc/n0 [34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u35  (
    .a(wb_ins_pc[37]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c35 ),
    .o({\cu_ru/m_s_epc/add0/c36 ,\cu_ru/m_s_epc/n0 [35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u36  (
    .a(wb_ins_pc[38]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c36 ),
    .o({\cu_ru/m_s_epc/add0/c37 ,\cu_ru/m_s_epc/n0 [36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u37  (
    .a(wb_ins_pc[39]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c37 ),
    .o({\cu_ru/m_s_epc/add0/c38 ,\cu_ru/m_s_epc/n0 [37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u38  (
    .a(wb_ins_pc[40]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c38 ),
    .o({\cu_ru/m_s_epc/add0/c39 ,\cu_ru/m_s_epc/n0 [38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u39  (
    .a(wb_ins_pc[41]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c39 ),
    .o({\cu_ru/m_s_epc/add0/c40 ,\cu_ru/m_s_epc/n0 [39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u4  (
    .a(wb_ins_pc[6]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c4 ),
    .o({\cu_ru/m_s_epc/add0/c5 ,\cu_ru/m_s_epc/n0 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u40  (
    .a(wb_ins_pc[42]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c40 ),
    .o({\cu_ru/m_s_epc/add0/c41 ,\cu_ru/m_s_epc/n0 [40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u41  (
    .a(wb_ins_pc[43]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c41 ),
    .o({\cu_ru/m_s_epc/add0/c42 ,\cu_ru/m_s_epc/n0 [41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u42  (
    .a(wb_ins_pc[44]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c42 ),
    .o({\cu_ru/m_s_epc/add0/c43 ,\cu_ru/m_s_epc/n0 [42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u43  (
    .a(wb_ins_pc[45]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c43 ),
    .o({\cu_ru/m_s_epc/add0/c44 ,\cu_ru/m_s_epc/n0 [43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u44  (
    .a(wb_ins_pc[46]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c44 ),
    .o({\cu_ru/m_s_epc/add0/c45 ,\cu_ru/m_s_epc/n0 [44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u45  (
    .a(wb_ins_pc[47]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c45 ),
    .o({\cu_ru/m_s_epc/add0/c46 ,\cu_ru/m_s_epc/n0 [45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u46  (
    .a(wb_ins_pc[48]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c46 ),
    .o({\cu_ru/m_s_epc/add0/c47 ,\cu_ru/m_s_epc/n0 [46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u47  (
    .a(wb_ins_pc[49]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c47 ),
    .o({\cu_ru/m_s_epc/add0/c48 ,\cu_ru/m_s_epc/n0 [47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u48  (
    .a(wb_ins_pc[50]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c48 ),
    .o({\cu_ru/m_s_epc/add0/c49 ,\cu_ru/m_s_epc/n0 [48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u49  (
    .a(wb_ins_pc[51]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c49 ),
    .o({\cu_ru/m_s_epc/add0/c50 ,\cu_ru/m_s_epc/n0 [49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u5  (
    .a(wb_ins_pc[7]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c5 ),
    .o({\cu_ru/m_s_epc/add0/c6 ,\cu_ru/m_s_epc/n0 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u50  (
    .a(wb_ins_pc[52]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c50 ),
    .o({\cu_ru/m_s_epc/add0/c51 ,\cu_ru/m_s_epc/n0 [50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u51  (
    .a(wb_ins_pc[53]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c51 ),
    .o({\cu_ru/m_s_epc/add0/c52 ,\cu_ru/m_s_epc/n0 [51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u52  (
    .a(wb_ins_pc[54]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c52 ),
    .o({\cu_ru/m_s_epc/add0/c53 ,\cu_ru/m_s_epc/n0 [52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u53  (
    .a(wb_ins_pc[55]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c53 ),
    .o({\cu_ru/m_s_epc/add0/c54 ,\cu_ru/m_s_epc/n0 [53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u54  (
    .a(wb_ins_pc[56]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c54 ),
    .o({\cu_ru/m_s_epc/add0/c55 ,\cu_ru/m_s_epc/n0 [54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u55  (
    .a(wb_ins_pc[57]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c55 ),
    .o({\cu_ru/m_s_epc/add0/c56 ,\cu_ru/m_s_epc/n0 [55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u56  (
    .a(wb_ins_pc[58]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c56 ),
    .o({\cu_ru/m_s_epc/add0/c57 ,\cu_ru/m_s_epc/n0 [56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u57  (
    .a(wb_ins_pc[59]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c57 ),
    .o({\cu_ru/m_s_epc/add0/c58 ,\cu_ru/m_s_epc/n0 [57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u58  (
    .a(wb_ins_pc[60]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c58 ),
    .o({\cu_ru/m_s_epc/add0/c59 ,\cu_ru/m_s_epc/n0 [58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u59  (
    .a(wb_ins_pc[61]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c59 ),
    .o({\cu_ru/m_s_epc/add0/c60 ,\cu_ru/m_s_epc/n0 [59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u6  (
    .a(wb_ins_pc[8]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c6 ),
    .o({\cu_ru/m_s_epc/add0/c7 ,\cu_ru/m_s_epc/n0 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u60  (
    .a(wb_ins_pc[62]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c60 ),
    .o({\cu_ru/m_s_epc/add0/c61 ,\cu_ru/m_s_epc/n0 [60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u61  (
    .a(wb_ins_pc[63]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c61 ),
    .o({open_n6074,\cu_ru/m_s_epc/n0 [61]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u7  (
    .a(wb_ins_pc[9]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c7 ),
    .o({\cu_ru/m_s_epc/add0/c8 ,\cu_ru/m_s_epc/n0 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u8  (
    .a(wb_ins_pc[10]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c8 ),
    .o({\cu_ru/m_s_epc/add0/c9 ,\cu_ru/m_s_epc/n0 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \cu_ru/m_s_epc/add0/u9  (
    .a(wb_ins_pc[11]),
    .b(1'b0),
    .c(\cu_ru/m_s_epc/add0/c9 ),
    .o({\cu_ru/m_s_epc/add0/c10 ,\cu_ru/m_s_epc/n0 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \cu_ru/m_s_epc/add0/ucin  (
    .a(1'b0),
    .o({\cu_ru/m_s_epc/add0/c0 ,open_n6077}));
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b0  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [0]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b1  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [1]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b10  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [10]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b11  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [11]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b12  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [12]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b13  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [13]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b14  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [14]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b15  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [15]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b16  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [16]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b17  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [17]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b18  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [18]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b19  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [19]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b2  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [2]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b20  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [20]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b21  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [21]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b22  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [22]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b23  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [23]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b24  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [24]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b25  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [25]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b26  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [26]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b27  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [27]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b28  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [28]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b29  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [29]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b3  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [3]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b30  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [30]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b31  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [31]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b32  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [32]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b33  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [33]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b34  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [34]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b35  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [35]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b36  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [36]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b37  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [37]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b38  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [38]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b39  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [39]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b4  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [4]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b40  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [40]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b41  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [41]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b42  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [42]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b43  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [43]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b44  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [44]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b45  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [45]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b46  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [46]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b47  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [47]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b48  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [48]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b49  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [49]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b5  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [5]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b50  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [50]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b51  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [51]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b52  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [52]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b53  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [53]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b54  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [54]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b55  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [55]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b56  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [56]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b57  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [57]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b58  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [58]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b59  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [59]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b6  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [6]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b60  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [60]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b61  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [61]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b62  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [62]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b63  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [63]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b7  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [7]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b8  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [8]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b9  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n8 [9]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sepc [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b0  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b1  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b10  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b11  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b12  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b13  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b14  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b15  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b16  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b17  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b18  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b19  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b2  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b20  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b21  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b22  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b23  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b24  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b25  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b26  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b27  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b28  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b29  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b3  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b30  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b31  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b32  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b33  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b34  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b35  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b36  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b37  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b38  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b39  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b4  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b40  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b41  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b42  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b43  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b44  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b45  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b46  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b47  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b48  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b49  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b5  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b50  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b51  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b52  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b53  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b54  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b55  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b56  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b57  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b58  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b59  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b6  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b60  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b61  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b62  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b63  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b7  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b8  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b9  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_epc/n10 [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mepc [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_ie/meie_reg  (
    .clk(clk_pad),
    .d(data_csr[11]),
    .en(\cu_ru/m_s_ie/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/m_sie [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  reg_sr_as_w1 \cu_ru/m_s_ie/msie_reg  (
    .clk(clk_pad),
    .d(data_csr[3]),
    .en(\cu_ru/m_s_ie/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/m_sie [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  reg_sr_as_w1 \cu_ru/m_s_ie/mtie_reg  (
    .clk(clk_pad),
    .d(data_csr[7]),
    .en(\cu_ru/m_s_ie/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/m_sie [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  reg_sr_as_w1 \cu_ru/m_s_ie/seie_reg  (
    .clk(clk_pad),
    .d(data_csr[9]),
    .en(~\cu_ru/m_s_ie/u11_sel_is_0_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/m_sie [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  reg_sr_as_w1 \cu_ru/m_s_ie/ssie_reg  (
    .clk(clk_pad),
    .d(data_csr[1]),
    .en(~\cu_ru/m_s_ie/u11_sel_is_0_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/m_sie [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  reg_sr_as_w1 \cu_ru/m_s_ie/stie_reg  (
    .clk(clk_pad),
    .d(data_csr[5]),
    .en(~\cu_ru/m_s_ie/u11_sel_is_0_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/m_sie [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IDDRPIPEMODE("NONE"),
    .INCEMUX("INV"),
    .INPCLKMUX("CLK"),
    .INRSTMUX("RST"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("RESET"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .SRMODE("SYNC"),
    .TSMUX("1"))
    \cu_ru/m_s_ip/meip_reg_IN  (
    .ce(\cu_ru/m_s_ip/u12_sel_is_2_o ),
    .ipad(m_ext_int),
    .ipclk(clk_pad),
    .rst(rst_pad),
    .diq({open_n6087,open_n6088,open_n6089,\cu_ru/m_sip [11]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IDDRPIPEMODE("NONE"),
    .INCEMUX("INV"),
    .INPCLKMUX("CLK"),
    .INRSTMUX("RST"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("RESET"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .SRMODE("SYNC"),
    .TSMUX("1"))
    \cu_ru/m_s_ip/msip_reg_IN  (
    .ce(\cu_ru/m_s_ip/u12_sel_is_2_o ),
    .ipad(m_soft_int),
    .ipclk(clk_pad),
    .rst(rst_pad),
    .diq({open_n6101,open_n6102,open_n6103,\cu_ru/m_sip [3]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IDDRPIPEMODE("NONE"),
    .INCEMUX("INV"),
    .INPCLKMUX("CLK"),
    .INRSTMUX("RST"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("RESET"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .SRMODE("SYNC"),
    .TSMUX("1"))
    \cu_ru/m_s_ip/mtip_reg_IN  (
    .ce(\cu_ru/m_s_ip/u12_sel_is_2_o ),
    .ipad(m_time_int),
    .ipclk(clk_pad),
    .rst(rst_pad),
    .diq({open_n6115,open_n6116,open_n6117,\cu_ru/m_sip [7]}));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  reg_sr_as_w1 \cu_ru/m_s_ip/seip_reg  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_ip/n1 ),
    .en(\cu_ru/m_s_ip/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/m_s_ip/seip ));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  reg_sr_as_w1 \cu_ru/m_s_ip/ssip_reg  (
    .clk(clk_pad),
    .d(data_csr[1]),
    .en(~\cu_ru/m_s_ip/u11_sel_is_0_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/m_sip [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  reg_sr_as_w1 \cu_ru/m_s_ip/stip_reg  (
    .clk(clk_pad),
    .d(data_csr[5]),
    .en(\cu_ru/m_s_ip/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/m_sip [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b0  (
    .clk(clk_pad),
    .d(data_csr[0]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b1  (
    .clk(clk_pad),
    .d(data_csr[1]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b10  (
    .clk(clk_pad),
    .d(data_csr[10]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b11  (
    .clk(clk_pad),
    .d(data_csr[11]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b12  (
    .clk(clk_pad),
    .d(data_csr[12]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b13  (
    .clk(clk_pad),
    .d(data_csr[13]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b14  (
    .clk(clk_pad),
    .d(data_csr[14]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b15  (
    .clk(clk_pad),
    .d(data_csr[15]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b16  (
    .clk(clk_pad),
    .d(data_csr[16]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b17  (
    .clk(clk_pad),
    .d(data_csr[17]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b18  (
    .clk(clk_pad),
    .d(data_csr[18]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b19  (
    .clk(clk_pad),
    .d(data_csr[19]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b2  (
    .clk(clk_pad),
    .d(data_csr[2]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b20  (
    .clk(clk_pad),
    .d(data_csr[20]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b21  (
    .clk(clk_pad),
    .d(data_csr[21]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b22  (
    .clk(clk_pad),
    .d(data_csr[22]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b23  (
    .clk(clk_pad),
    .d(data_csr[23]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b24  (
    .clk(clk_pad),
    .d(data_csr[24]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b25  (
    .clk(clk_pad),
    .d(data_csr[25]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b26  (
    .clk(clk_pad),
    .d(data_csr[26]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b27  (
    .clk(clk_pad),
    .d(data_csr[27]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b28  (
    .clk(clk_pad),
    .d(data_csr[28]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b29  (
    .clk(clk_pad),
    .d(data_csr[29]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b3  (
    .clk(clk_pad),
    .d(data_csr[3]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b30  (
    .clk(clk_pad),
    .d(data_csr[30]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b31  (
    .clk(clk_pad),
    .d(data_csr[31]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b32  (
    .clk(clk_pad),
    .d(data_csr[32]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b33  (
    .clk(clk_pad),
    .d(data_csr[33]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b34  (
    .clk(clk_pad),
    .d(data_csr[34]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b35  (
    .clk(clk_pad),
    .d(data_csr[35]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b36  (
    .clk(clk_pad),
    .d(data_csr[36]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b37  (
    .clk(clk_pad),
    .d(data_csr[37]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b38  (
    .clk(clk_pad),
    .d(data_csr[38]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b39  (
    .clk(clk_pad),
    .d(data_csr[39]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b4  (
    .clk(clk_pad),
    .d(data_csr[4]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b40  (
    .clk(clk_pad),
    .d(data_csr[40]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b41  (
    .clk(clk_pad),
    .d(data_csr[41]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b42  (
    .clk(clk_pad),
    .d(data_csr[42]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b43  (
    .clk(clk_pad),
    .d(data_csr[43]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b44  (
    .clk(clk_pad),
    .d(data_csr[44]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b45  (
    .clk(clk_pad),
    .d(data_csr[45]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b46  (
    .clk(clk_pad),
    .d(data_csr[46]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b47  (
    .clk(clk_pad),
    .d(data_csr[47]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b48  (
    .clk(clk_pad),
    .d(data_csr[48]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b49  (
    .clk(clk_pad),
    .d(data_csr[49]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b5  (
    .clk(clk_pad),
    .d(data_csr[5]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b50  (
    .clk(clk_pad),
    .d(data_csr[50]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b51  (
    .clk(clk_pad),
    .d(data_csr[51]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b52  (
    .clk(clk_pad),
    .d(data_csr[52]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b53  (
    .clk(clk_pad),
    .d(data_csr[53]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b54  (
    .clk(clk_pad),
    .d(data_csr[54]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b55  (
    .clk(clk_pad),
    .d(data_csr[55]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b56  (
    .clk(clk_pad),
    .d(data_csr[56]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b57  (
    .clk(clk_pad),
    .d(data_csr[57]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b58  (
    .clk(clk_pad),
    .d(data_csr[58]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b59  (
    .clk(clk_pad),
    .d(data_csr[59]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b6  (
    .clk(clk_pad),
    .d(data_csr[6]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b60  (
    .clk(clk_pad),
    .d(data_csr[60]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b61  (
    .clk(clk_pad),
    .d(data_csr[61]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b62  (
    .clk(clk_pad),
    .d(data_csr[62]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b63  (
    .clk(clk_pad),
    .d(data_csr[63]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b7  (
    .clk(clk_pad),
    .d(data_csr[7]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b8  (
    .clk(clk_pad),
    .d(data_csr[8]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b9  (
    .clk(clk_pad),
    .d(data_csr[9]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mscratch [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b0  (
    .clk(clk_pad),
    .d(data_csr[0]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b1  (
    .clk(clk_pad),
    .d(data_csr[1]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b10  (
    .clk(clk_pad),
    .d(data_csr[10]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b11  (
    .clk(clk_pad),
    .d(data_csr[11]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b12  (
    .clk(clk_pad),
    .d(data_csr[12]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b13  (
    .clk(clk_pad),
    .d(data_csr[13]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b14  (
    .clk(clk_pad),
    .d(data_csr[14]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b15  (
    .clk(clk_pad),
    .d(data_csr[15]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b16  (
    .clk(clk_pad),
    .d(data_csr[16]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b17  (
    .clk(clk_pad),
    .d(data_csr[17]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b18  (
    .clk(clk_pad),
    .d(data_csr[18]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b19  (
    .clk(clk_pad),
    .d(data_csr[19]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b2  (
    .clk(clk_pad),
    .d(data_csr[2]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b20  (
    .clk(clk_pad),
    .d(data_csr[20]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b21  (
    .clk(clk_pad),
    .d(data_csr[21]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b22  (
    .clk(clk_pad),
    .d(data_csr[22]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b23  (
    .clk(clk_pad),
    .d(data_csr[23]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b24  (
    .clk(clk_pad),
    .d(data_csr[24]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b25  (
    .clk(clk_pad),
    .d(data_csr[25]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b26  (
    .clk(clk_pad),
    .d(data_csr[26]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b27  (
    .clk(clk_pad),
    .d(data_csr[27]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b28  (
    .clk(clk_pad),
    .d(data_csr[28]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b29  (
    .clk(clk_pad),
    .d(data_csr[29]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b3  (
    .clk(clk_pad),
    .d(data_csr[3]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b30  (
    .clk(clk_pad),
    .d(data_csr[30]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b31  (
    .clk(clk_pad),
    .d(data_csr[31]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b32  (
    .clk(clk_pad),
    .d(data_csr[32]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b33  (
    .clk(clk_pad),
    .d(data_csr[33]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b34  (
    .clk(clk_pad),
    .d(data_csr[34]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b35  (
    .clk(clk_pad),
    .d(data_csr[35]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b36  (
    .clk(clk_pad),
    .d(data_csr[36]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b37  (
    .clk(clk_pad),
    .d(data_csr[37]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b38  (
    .clk(clk_pad),
    .d(data_csr[38]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b39  (
    .clk(clk_pad),
    .d(data_csr[39]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b4  (
    .clk(clk_pad),
    .d(data_csr[4]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b40  (
    .clk(clk_pad),
    .d(data_csr[40]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b41  (
    .clk(clk_pad),
    .d(data_csr[41]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b42  (
    .clk(clk_pad),
    .d(data_csr[42]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b43  (
    .clk(clk_pad),
    .d(data_csr[43]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b44  (
    .clk(clk_pad),
    .d(data_csr[44]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b45  (
    .clk(clk_pad),
    .d(data_csr[45]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b46  (
    .clk(clk_pad),
    .d(data_csr[46]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b47  (
    .clk(clk_pad),
    .d(data_csr[47]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b48  (
    .clk(clk_pad),
    .d(data_csr[48]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b49  (
    .clk(clk_pad),
    .d(data_csr[49]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b5  (
    .clk(clk_pad),
    .d(data_csr[5]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b50  (
    .clk(clk_pad),
    .d(data_csr[50]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b51  (
    .clk(clk_pad),
    .d(data_csr[51]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b52  (
    .clk(clk_pad),
    .d(data_csr[52]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b53  (
    .clk(clk_pad),
    .d(data_csr[53]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b54  (
    .clk(clk_pad),
    .d(data_csr[54]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b55  (
    .clk(clk_pad),
    .d(data_csr[55]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b56  (
    .clk(clk_pad),
    .d(data_csr[56]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b57  (
    .clk(clk_pad),
    .d(data_csr[57]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b58  (
    .clk(clk_pad),
    .d(data_csr[58]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b59  (
    .clk(clk_pad),
    .d(data_csr[59]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b6  (
    .clk(clk_pad),
    .d(data_csr[6]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b60  (
    .clk(clk_pad),
    .d(data_csr[60]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b61  (
    .clk(clk_pad),
    .d(data_csr[61]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b62  (
    .clk(clk_pad),
    .d(data_csr[62]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b63  (
    .clk(clk_pad),
    .d(data_csr[63]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b7  (
    .clk(clk_pad),
    .d(data_csr[7]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b8  (
    .clk(clk_pad),
    .d(data_csr[8]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b9  (
    .clk(clk_pad),
    .d(data_csr[9]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/sscratch [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_status/mie_reg  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_status/n37 ),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mie ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/mpie_reg  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_status/n45 ),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mstatus [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/mprv_reg  (
    .clk(clk_pad),
    .d(data_csr[17]),
    .en(\cu_ru/m_s_status/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(mprv));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/mxr_reg  (
    .clk(clk_pad),
    .d(data_csr[19]),
    .en(~\cu_ru/m_s_status/u34_sel_is_0_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(mxr));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/reg0_b0  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_status/n47 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mstatus [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/reg0_b1  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_status/n47 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mstatus [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/reg1_b0  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_status/n64 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(priv[0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  reg_sr_as_w1 \cu_ru/m_s_status/reg1_b1  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_status/n64 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(priv[1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  reg_ar_ss_w1 \cu_ru/m_s_status/reg1_b3  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_status/n64 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(rst_pad),
    .q(priv[3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  reg_sr_as_w1 \cu_ru/m_s_status/sie_reg  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_status/n36 ),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mstatus [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/spie_reg  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_status/n44 ),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mstatus [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/spp_reg  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_status/n46 ),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mstatus [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/sum_reg  (
    .clk(clk_pad),
    .d(data_csr[18]),
    .en(~\cu_ru/m_s_status/u34_sel_is_0_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(sum));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/tsr_reg  (
    .clk(clk_pad),
    .d(data_csr[22]),
    .en(\cu_ru/m_s_status/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(tsr));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/tvm_reg  (
    .clk(clk_pad),
    .d(data_csr[20]),
    .en(\cu_ru/m_s_status/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(tvm));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/tw_reg  (
    .clk(clk_pad),
    .d(data_csr[21]),
    .en(\cu_ru/m_s_status/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(tw));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b0  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [0]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b1  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [1]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b10  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [10]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b11  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [11]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b12  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [12]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b13  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [13]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b14  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [14]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b15  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [15]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b16  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [16]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b17  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [17]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b18  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [18]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b19  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [19]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b2  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [2]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b20  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [20]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b21  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [21]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b22  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [22]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b23  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [23]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b24  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [24]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b25  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [25]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b26  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [26]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b27  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [27]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b28  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [28]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b29  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [29]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b3  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [3]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b30  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [30]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b31  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [31]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b32  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [32]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b33  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [33]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b34  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [34]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b35  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [35]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b36  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [36]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b37  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [37]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b38  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [38]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b39  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [39]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b4  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [4]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b40  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [40]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b41  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [41]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b42  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [42]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b43  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [43]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b44  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [44]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b45  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [45]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b46  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [46]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b47  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [47]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b48  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [48]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b49  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [49]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b5  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [5]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b50  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [50]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b51  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [51]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b52  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [52]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b53  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [53]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b54  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [54]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b55  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [55]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b56  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [56]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b57  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [57]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b58  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [58]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b59  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [59]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b6  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [6]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b60  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [60]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b61  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [61]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b62  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [62]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b63  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [63]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b7  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [7]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b8  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [8]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b9  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n9 [9]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stval [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b0  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b1  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b10  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b11  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b12  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b13  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b14  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b15  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b16  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b17  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b18  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b19  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b2  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b20  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b21  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b22  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b23  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b24  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b25  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b26  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b27  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b28  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b29  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b3  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b30  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b31  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b32  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b33  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b34  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b35  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b36  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b37  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b38  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b39  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b4  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b40  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b41  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b42  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b43  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b44  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b45  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b46  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b47  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b48  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b49  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b5  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b50  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b51  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b52  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b53  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b54  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b55  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b56  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b57  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b58  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b59  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b6  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b60  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b61  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b62  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b63  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b7  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b8  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b9  (
    .clk(clk_pad),
    .d(\cu_ru/m_s_tval/n11 [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtval [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b0  (
    .clk(clk_pad),
    .d(csr_data[0]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b1  (
    .clk(clk_pad),
    .d(csr_data[1]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b10  (
    .clk(clk_pad),
    .d(csr_data[10]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b11  (
    .clk(clk_pad),
    .d(csr_data[11]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b12  (
    .clk(clk_pad),
    .d(csr_data[12]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b13  (
    .clk(clk_pad),
    .d(csr_data[13]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b14  (
    .clk(clk_pad),
    .d(csr_data[14]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b15  (
    .clk(clk_pad),
    .d(csr_data[15]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b16  (
    .clk(clk_pad),
    .d(csr_data[16]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b17  (
    .clk(clk_pad),
    .d(csr_data[17]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b18  (
    .clk(clk_pad),
    .d(csr_data[18]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b19  (
    .clk(clk_pad),
    .d(csr_data[19]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b2  (
    .clk(clk_pad),
    .d(csr_data[2]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b20  (
    .clk(clk_pad),
    .d(csr_data[20]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b21  (
    .clk(clk_pad),
    .d(csr_data[21]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b22  (
    .clk(clk_pad),
    .d(csr_data[22]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b23  (
    .clk(clk_pad),
    .d(csr_data[23]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b24  (
    .clk(clk_pad),
    .d(csr_data[24]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b25  (
    .clk(clk_pad),
    .d(csr_data[25]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b26  (
    .clk(clk_pad),
    .d(csr_data[26]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b27  (
    .clk(clk_pad),
    .d(csr_data[27]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b28  (
    .clk(clk_pad),
    .d(csr_data[28]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b29  (
    .clk(clk_pad),
    .d(csr_data[29]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b3  (
    .clk(clk_pad),
    .d(csr_data[3]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b30  (
    .clk(clk_pad),
    .d(csr_data[30]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b31  (
    .clk(clk_pad),
    .d(csr_data[31]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b32  (
    .clk(clk_pad),
    .d(csr_data[32]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b33  (
    .clk(clk_pad),
    .d(csr_data[33]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b34  (
    .clk(clk_pad),
    .d(csr_data[34]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b35  (
    .clk(clk_pad),
    .d(csr_data[35]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b36  (
    .clk(clk_pad),
    .d(csr_data[36]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b37  (
    .clk(clk_pad),
    .d(csr_data[37]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b38  (
    .clk(clk_pad),
    .d(csr_data[38]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b39  (
    .clk(clk_pad),
    .d(csr_data[39]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b4  (
    .clk(clk_pad),
    .d(csr_data[4]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b40  (
    .clk(clk_pad),
    .d(csr_data[40]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b41  (
    .clk(clk_pad),
    .d(csr_data[41]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b42  (
    .clk(clk_pad),
    .d(csr_data[42]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b43  (
    .clk(clk_pad),
    .d(csr_data[43]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b44  (
    .clk(clk_pad),
    .d(csr_data[44]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b45  (
    .clk(clk_pad),
    .d(csr_data[45]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b46  (
    .clk(clk_pad),
    .d(csr_data[46]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b47  (
    .clk(clk_pad),
    .d(csr_data[47]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b48  (
    .clk(clk_pad),
    .d(csr_data[48]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b49  (
    .clk(clk_pad),
    .d(csr_data[49]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b5  (
    .clk(clk_pad),
    .d(csr_data[5]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b50  (
    .clk(clk_pad),
    .d(csr_data[50]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b51  (
    .clk(clk_pad),
    .d(csr_data[51]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b52  (
    .clk(clk_pad),
    .d(csr_data[52]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b53  (
    .clk(clk_pad),
    .d(csr_data[53]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b54  (
    .clk(clk_pad),
    .d(csr_data[54]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b55  (
    .clk(clk_pad),
    .d(csr_data[55]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b56  (
    .clk(clk_pad),
    .d(csr_data[56]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b57  (
    .clk(clk_pad),
    .d(csr_data[57]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b58  (
    .clk(clk_pad),
    .d(csr_data[58]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b59  (
    .clk(clk_pad),
    .d(csr_data[59]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b6  (
    .clk(clk_pad),
    .d(csr_data[6]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b60  (
    .clk(clk_pad),
    .d(csr_data[60]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b61  (
    .clk(clk_pad),
    .d(csr_data[61]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b62  (
    .clk(clk_pad),
    .d(csr_data[62]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b63  (
    .clk(clk_pad),
    .d(csr_data[63]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b7  (
    .clk(clk_pad),
    .d(csr_data[7]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b8  (
    .clk(clk_pad),
    .d(csr_data[8]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b9  (
    .clk(clk_pad),
    .d(csr_data[9]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/stvec [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b0  (
    .clk(clk_pad),
    .d(csr_data[0]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b1  (
    .clk(clk_pad),
    .d(csr_data[1]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b10  (
    .clk(clk_pad),
    .d(csr_data[10]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b11  (
    .clk(clk_pad),
    .d(csr_data[11]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b12  (
    .clk(clk_pad),
    .d(csr_data[12]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b13  (
    .clk(clk_pad),
    .d(csr_data[13]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b14  (
    .clk(clk_pad),
    .d(csr_data[14]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b15  (
    .clk(clk_pad),
    .d(csr_data[15]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b16  (
    .clk(clk_pad),
    .d(csr_data[16]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b17  (
    .clk(clk_pad),
    .d(csr_data[17]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b18  (
    .clk(clk_pad),
    .d(csr_data[18]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b19  (
    .clk(clk_pad),
    .d(csr_data[19]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b2  (
    .clk(clk_pad),
    .d(csr_data[2]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b20  (
    .clk(clk_pad),
    .d(csr_data[20]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b21  (
    .clk(clk_pad),
    .d(csr_data[21]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b22  (
    .clk(clk_pad),
    .d(csr_data[22]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b23  (
    .clk(clk_pad),
    .d(csr_data[23]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b24  (
    .clk(clk_pad),
    .d(csr_data[24]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b25  (
    .clk(clk_pad),
    .d(csr_data[25]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b26  (
    .clk(clk_pad),
    .d(csr_data[26]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b27  (
    .clk(clk_pad),
    .d(csr_data[27]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b28  (
    .clk(clk_pad),
    .d(csr_data[28]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b29  (
    .clk(clk_pad),
    .d(csr_data[29]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b3  (
    .clk(clk_pad),
    .d(csr_data[3]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b30  (
    .clk(clk_pad),
    .d(csr_data[30]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b31  (
    .clk(clk_pad),
    .d(csr_data[31]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b32  (
    .clk(clk_pad),
    .d(csr_data[32]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b33  (
    .clk(clk_pad),
    .d(csr_data[33]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b34  (
    .clk(clk_pad),
    .d(csr_data[34]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b35  (
    .clk(clk_pad),
    .d(csr_data[35]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b36  (
    .clk(clk_pad),
    .d(csr_data[36]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b37  (
    .clk(clk_pad),
    .d(csr_data[37]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b38  (
    .clk(clk_pad),
    .d(csr_data[38]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b39  (
    .clk(clk_pad),
    .d(csr_data[39]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b4  (
    .clk(clk_pad),
    .d(csr_data[4]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b40  (
    .clk(clk_pad),
    .d(csr_data[40]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b41  (
    .clk(clk_pad),
    .d(csr_data[41]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b42  (
    .clk(clk_pad),
    .d(csr_data[42]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b43  (
    .clk(clk_pad),
    .d(csr_data[43]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b44  (
    .clk(clk_pad),
    .d(csr_data[44]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b45  (
    .clk(clk_pad),
    .d(csr_data[45]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b46  (
    .clk(clk_pad),
    .d(csr_data[46]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b47  (
    .clk(clk_pad),
    .d(csr_data[47]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b48  (
    .clk(clk_pad),
    .d(csr_data[48]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b49  (
    .clk(clk_pad),
    .d(csr_data[49]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b5  (
    .clk(clk_pad),
    .d(csr_data[5]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b50  (
    .clk(clk_pad),
    .d(csr_data[50]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b51  (
    .clk(clk_pad),
    .d(csr_data[51]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b52  (
    .clk(clk_pad),
    .d(csr_data[52]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b53  (
    .clk(clk_pad),
    .d(csr_data[53]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b54  (
    .clk(clk_pad),
    .d(csr_data[54]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b55  (
    .clk(clk_pad),
    .d(csr_data[55]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b56  (
    .clk(clk_pad),
    .d(csr_data[56]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b57  (
    .clk(clk_pad),
    .d(csr_data[57]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b58  (
    .clk(clk_pad),
    .d(csr_data[58]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b59  (
    .clk(clk_pad),
    .d(csr_data[59]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b6  (
    .clk(clk_pad),
    .d(csr_data[6]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b60  (
    .clk(clk_pad),
    .d(csr_data[60]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b61  (
    .clk(clk_pad),
    .d(csr_data[61]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b62  (
    .clk(clk_pad),
    .d(csr_data[62]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b63  (
    .clk(clk_pad),
    .d(csr_data[63]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b7  (
    .clk(clk_pad),
    .d(csr_data[7]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b8  (
    .clk(clk_pad),
    .d(csr_data[8]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b9  (
    .clk(clk_pad),
    .d(csr_data[9]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mtvec [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dbk_reg  (
    .clk(clk_pad),
    .d(data_csr[3]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [3]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/decs_reg  (
    .clk(clk_pad),
    .d(data_csr[9]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [9]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/decu_reg  (
    .clk(clk_pad),
    .d(data_csr[8]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [8]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/diaf_reg  (
    .clk(clk_pad),
    .d(data_csr[1]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [1]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/diam_reg  (
    .clk(clk_pad),
    .d(data_csr[0]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [0]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dii_reg  (
    .clk(clk_pad),
    .d(data_csr[2]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [2]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dipf_reg  (
    .clk(clk_pad),
    .d(data_csr[12]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [12]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dlaf_reg  (
    .clk(clk_pad),
    .d(data_csr[5]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [5]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dlam_reg  (
    .clk(clk_pad),
    .d(data_csr[4]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [4]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dlpf_reg  (
    .clk(clk_pad),
    .d(data_csr[13]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [13]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dsaf_reg  (
    .clk(clk_pad),
    .d(data_csr[7]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [7]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dsam_reg  (
    .clk(clk_pad),
    .d(data_csr[6]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [6]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dspf_reg  (
    .clk(clk_pad),
    .d(data_csr[15]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/medeleg [15]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/mideleg_int_ctrl/dsei_reg  (
    .clk(clk_pad),
    .d(data_csr[9]),
    .en(\cu_ru/mideleg_int_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mideleg [9]));  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  reg_sr_as_w1 \cu_ru/mideleg_int_ctrl/dssi_reg  (
    .clk(clk_pad),
    .d(data_csr[1]),
    .en(\cu_ru/mideleg_int_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mideleg [1]));  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  reg_sr_as_w1 \cu_ru/mideleg_int_ctrl/dsti_reg  (
    .clk(clk_pad),
    .d(data_csr[5]),
    .en(\cu_ru/mideleg_int_ctrl/n0 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\cu_ru/mideleg [5]));  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub0/u0  (
    .a(id_rs1_index[0]),
    .b(1'b1),
    .c(\cu_ru/sub0/c0 ),
    .o({\cu_ru/sub0/c1 ,\cu_ru/n46 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub0/u1  (
    .a(id_rs1_index[1]),
    .b(1'b0),
    .c(\cu_ru/sub0/c1 ),
    .o({\cu_ru/sub0/c2 ,\cu_ru/n46 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub0/u2  (
    .a(id_rs1_index[2]),
    .b(1'b0),
    .c(\cu_ru/sub0/c2 ),
    .o({\cu_ru/sub0/c3 ,\cu_ru/n46 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub0/u3  (
    .a(id_rs1_index[3]),
    .b(1'b0),
    .c(\cu_ru/sub0/c3 ),
    .o({\cu_ru/sub0/c4 ,\cu_ru/n46 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub0/u4  (
    .a(id_rs1_index[4]),
    .b(1'b0),
    .c(\cu_ru/sub0/c4 ),
    .o({open_n6120,\cu_ru/n46 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \cu_ru/sub0/ucin  (
    .a(1'b0),
    .o({\cu_ru/sub0/c0 ,open_n6123}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub1/u0  (
    .a(id_rs2_index[0]),
    .b(1'b1),
    .c(\cu_ru/sub1/c0 ),
    .o({\cu_ru/sub1/c1 ,\cu_ru/n49 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub1/u1  (
    .a(id_rs2_index[1]),
    .b(1'b0),
    .c(\cu_ru/sub1/c1 ),
    .o({\cu_ru/sub1/c2 ,\cu_ru/n49 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub1/u2  (
    .a(id_rs2_index[2]),
    .b(1'b0),
    .c(\cu_ru/sub1/c2 ),
    .o({\cu_ru/sub1/c3 ,\cu_ru/n49 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub1/u3  (
    .a(id_rs2_index[3]),
    .b(1'b0),
    .c(\cu_ru/sub1/c3 ),
    .o({\cu_ru/sub1/c4 ,\cu_ru/n49 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub1/u4  (
    .a(id_rs2_index[4]),
    .b(1'b0),
    .c(\cu_ru/sub1/c4 ),
    .o({open_n6124,\cu_ru/n49 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \cu_ru/sub1/ucin  (
    .a(1'b0),
    .o({\cu_ru/sub1/c0 ,open_n6127}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub2/u0  (
    .a(wb_rd_index[0]),
    .b(1'b1),
    .c(\cu_ru/sub2/c0 ),
    .o({\cu_ru/sub2/c1 ,\cu_ru/n52 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub2/u1  (
    .a(wb_rd_index[1]),
    .b(1'b0),
    .c(\cu_ru/sub2/c1 ),
    .o({\cu_ru/sub2/c2 ,\cu_ru/n52 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub2/u2  (
    .a(wb_rd_index[2]),
    .b(1'b0),
    .c(\cu_ru/sub2/c2 ),
    .o({\cu_ru/sub2/c3 ,\cu_ru/n52 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub2/u3  (
    .a(wb_rd_index[3]),
    .b(1'b0),
    .c(\cu_ru/sub2/c3 ),
    .o({\cu_ru/sub2/c4 ,\cu_ru/n52 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \cu_ru/sub2/u4  (
    .a(wb_rd_index[4]),
    .b(1'b0),
    .c(\cu_ru/sub2/c4 ),
    .o({open_n6128,\cu_ru/n52 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \cu_ru/sub2/ucin  (
    .a(1'b0),
    .o({\cu_ru/sub2/c0 ,open_n6131}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u0  (
    .a(ds1[0]),
    .b(\exu/alu_au/n17 [0]),
    .c(\exu/alu_au/add0/c0 ),
    .o({\exu/alu_au/add0/c1 ,\exu/alu_au/add_64 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u1  (
    .a(ds1[1]),
    .b(\exu/alu_au/n17 [1]),
    .c(\exu/alu_au/add0/c1 ),
    .o({\exu/alu_au/add0/c2 ,\exu/alu_au/add_64 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u10  (
    .a(ds1[10]),
    .b(\exu/alu_au/n17 [10]),
    .c(\exu/alu_au/add0/c10 ),
    .o({\exu/alu_au/add0/c11 ,\exu/alu_au/add_64 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u11  (
    .a(ds1[11]),
    .b(\exu/alu_au/n17 [11]),
    .c(\exu/alu_au/add0/c11 ),
    .o({\exu/alu_au/add0/c12 ,\exu/alu_au/add_64 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u12  (
    .a(ds1[12]),
    .b(\exu/alu_au/n17 [12]),
    .c(\exu/alu_au/add0/c12 ),
    .o({\exu/alu_au/add0/c13 ,\exu/alu_au/add_64 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u13  (
    .a(ds1[13]),
    .b(\exu/alu_au/n17 [13]),
    .c(\exu/alu_au/add0/c13 ),
    .o({\exu/alu_au/add0/c14 ,\exu/alu_au/add_64 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u14  (
    .a(ds1[14]),
    .b(\exu/alu_au/n17 [14]),
    .c(\exu/alu_au/add0/c14 ),
    .o({\exu/alu_au/add0/c15 ,\exu/alu_au/add_64 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u15  (
    .a(ds1[15]),
    .b(\exu/alu_au/n17 [15]),
    .c(\exu/alu_au/add0/c15 ),
    .o({\exu/alu_au/add0/c16 ,\exu/alu_au/add_64 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u16  (
    .a(ds1[16]),
    .b(\exu/alu_au/n17 [16]),
    .c(\exu/alu_au/add0/c16 ),
    .o({\exu/alu_au/add0/c17 ,\exu/alu_au/add_64 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u17  (
    .a(ds1[17]),
    .b(\exu/alu_au/n17 [17]),
    .c(\exu/alu_au/add0/c17 ),
    .o({\exu/alu_au/add0/c18 ,\exu/alu_au/add_64 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u18  (
    .a(ds1[18]),
    .b(\exu/alu_au/n17 [18]),
    .c(\exu/alu_au/add0/c18 ),
    .o({\exu/alu_au/add0/c19 ,\exu/alu_au/add_64 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u19  (
    .a(ds1[19]),
    .b(\exu/alu_au/n17 [19]),
    .c(\exu/alu_au/add0/c19 ),
    .o({\exu/alu_au/add0/c20 ,\exu/alu_au/add_64 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u2  (
    .a(ds1[2]),
    .b(\exu/alu_au/n17 [2]),
    .c(\exu/alu_au/add0/c2 ),
    .o({\exu/alu_au/add0/c3 ,\exu/alu_au/add_64 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u20  (
    .a(ds1[20]),
    .b(\exu/alu_au/n17 [20]),
    .c(\exu/alu_au/add0/c20 ),
    .o({\exu/alu_au/add0/c21 ,\exu/alu_au/add_64 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u21  (
    .a(ds1[21]),
    .b(\exu/alu_au/n17 [21]),
    .c(\exu/alu_au/add0/c21 ),
    .o({\exu/alu_au/add0/c22 ,\exu/alu_au/add_64 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u22  (
    .a(ds1[22]),
    .b(\exu/alu_au/n17 [22]),
    .c(\exu/alu_au/add0/c22 ),
    .o({\exu/alu_au/add0/c23 ,\exu/alu_au/add_64 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u23  (
    .a(ds1[23]),
    .b(\exu/alu_au/n17 [23]),
    .c(\exu/alu_au/add0/c23 ),
    .o({\exu/alu_au/add0/c24 ,\exu/alu_au/add_64 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u24  (
    .a(ds1[24]),
    .b(\exu/alu_au/n17 [24]),
    .c(\exu/alu_au/add0/c24 ),
    .o({\exu/alu_au/add0/c25 ,\exu/alu_au/add_64 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u25  (
    .a(ds1[25]),
    .b(\exu/alu_au/n17 [25]),
    .c(\exu/alu_au/add0/c25 ),
    .o({\exu/alu_au/add0/c26 ,\exu/alu_au/add_64 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u26  (
    .a(ds1[26]),
    .b(\exu/alu_au/n17 [26]),
    .c(\exu/alu_au/add0/c26 ),
    .o({\exu/alu_au/add0/c27 ,\exu/alu_au/add_64 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u27  (
    .a(ds1[27]),
    .b(\exu/alu_au/n17 [27]),
    .c(\exu/alu_au/add0/c27 ),
    .o({\exu/alu_au/add0/c28 ,\exu/alu_au/add_64 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u28  (
    .a(ds1[28]),
    .b(\exu/alu_au/n17 [28]),
    .c(\exu/alu_au/add0/c28 ),
    .o({\exu/alu_au/add0/c29 ,\exu/alu_au/add_64 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u29  (
    .a(ds1[29]),
    .b(\exu/alu_au/n17 [29]),
    .c(\exu/alu_au/add0/c29 ),
    .o({\exu/alu_au/add0/c30 ,\exu/alu_au/add_64 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u3  (
    .a(ds1[3]),
    .b(\exu/alu_au/n17 [3]),
    .c(\exu/alu_au/add0/c3 ),
    .o({\exu/alu_au/add0/c4 ,\exu/alu_au/add_64 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u30  (
    .a(ds1[30]),
    .b(\exu/alu_au/n17 [30]),
    .c(\exu/alu_au/add0/c30 ),
    .o({\exu/alu_au/add0/c31 ,\exu/alu_au/add_64 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u31  (
    .a(ds1[31]),
    .b(\exu/alu_au/n17 [31]),
    .c(\exu/alu_au/add0/c31 ),
    .o({\exu/alu_au/add0/c32 ,\exu/alu_au/add_64 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u32  (
    .a(ds1[32]),
    .b(\exu/alu_au/n17 [32]),
    .c(\exu/alu_au/add0/c32 ),
    .o({\exu/alu_au/add0/c33 ,\exu/alu_au/add_64 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u33  (
    .a(ds1[33]),
    .b(\exu/alu_au/n17 [33]),
    .c(\exu/alu_au/add0/c33 ),
    .o({\exu/alu_au/add0/c34 ,\exu/alu_au/add_64 [33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u34  (
    .a(ds1[34]),
    .b(\exu/alu_au/n17 [34]),
    .c(\exu/alu_au/add0/c34 ),
    .o({\exu/alu_au/add0/c35 ,\exu/alu_au/add_64 [34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u35  (
    .a(ds1[35]),
    .b(\exu/alu_au/n17 [35]),
    .c(\exu/alu_au/add0/c35 ),
    .o({\exu/alu_au/add0/c36 ,\exu/alu_au/add_64 [35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u36  (
    .a(ds1[36]),
    .b(\exu/alu_au/n17 [36]),
    .c(\exu/alu_au/add0/c36 ),
    .o({\exu/alu_au/add0/c37 ,\exu/alu_au/add_64 [36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u37  (
    .a(ds1[37]),
    .b(\exu/alu_au/n17 [37]),
    .c(\exu/alu_au/add0/c37 ),
    .o({\exu/alu_au/add0/c38 ,\exu/alu_au/add_64 [37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u38  (
    .a(ds1[38]),
    .b(\exu/alu_au/n17 [38]),
    .c(\exu/alu_au/add0/c38 ),
    .o({\exu/alu_au/add0/c39 ,\exu/alu_au/add_64 [38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u39  (
    .a(ds1[39]),
    .b(\exu/alu_au/n17 [39]),
    .c(\exu/alu_au/add0/c39 ),
    .o({\exu/alu_au/add0/c40 ,\exu/alu_au/add_64 [39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u4  (
    .a(ds1[4]),
    .b(\exu/alu_au/n17 [4]),
    .c(\exu/alu_au/add0/c4 ),
    .o({\exu/alu_au/add0/c5 ,\exu/alu_au/add_64 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u40  (
    .a(ds1[40]),
    .b(\exu/alu_au/n17 [40]),
    .c(\exu/alu_au/add0/c40 ),
    .o({\exu/alu_au/add0/c41 ,\exu/alu_au/add_64 [40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u41  (
    .a(ds1[41]),
    .b(\exu/alu_au/n17 [41]),
    .c(\exu/alu_au/add0/c41 ),
    .o({\exu/alu_au/add0/c42 ,\exu/alu_au/add_64 [41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u42  (
    .a(ds1[42]),
    .b(\exu/alu_au/n17 [42]),
    .c(\exu/alu_au/add0/c42 ),
    .o({\exu/alu_au/add0/c43 ,\exu/alu_au/add_64 [42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u43  (
    .a(ds1[43]),
    .b(\exu/alu_au/n17 [43]),
    .c(\exu/alu_au/add0/c43 ),
    .o({\exu/alu_au/add0/c44 ,\exu/alu_au/add_64 [43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u44  (
    .a(ds1[44]),
    .b(\exu/alu_au/n17 [44]),
    .c(\exu/alu_au/add0/c44 ),
    .o({\exu/alu_au/add0/c45 ,\exu/alu_au/add_64 [44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u45  (
    .a(ds1[45]),
    .b(\exu/alu_au/n17 [45]),
    .c(\exu/alu_au/add0/c45 ),
    .o({\exu/alu_au/add0/c46 ,\exu/alu_au/add_64 [45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u46  (
    .a(ds1[46]),
    .b(\exu/alu_au/n17 [46]),
    .c(\exu/alu_au/add0/c46 ),
    .o({\exu/alu_au/add0/c47 ,\exu/alu_au/add_64 [46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u47  (
    .a(ds1[47]),
    .b(\exu/alu_au/n17 [47]),
    .c(\exu/alu_au/add0/c47 ),
    .o({\exu/alu_au/add0/c48 ,\exu/alu_au/add_64 [47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u48  (
    .a(ds1[48]),
    .b(\exu/alu_au/n17 [48]),
    .c(\exu/alu_au/add0/c48 ),
    .o({\exu/alu_au/add0/c49 ,\exu/alu_au/add_64 [48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u49  (
    .a(ds1[49]),
    .b(\exu/alu_au/n17 [49]),
    .c(\exu/alu_au/add0/c49 ),
    .o({\exu/alu_au/add0/c50 ,\exu/alu_au/add_64 [49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u5  (
    .a(ds1[5]),
    .b(\exu/alu_au/n17 [5]),
    .c(\exu/alu_au/add0/c5 ),
    .o({\exu/alu_au/add0/c6 ,\exu/alu_au/add_64 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u50  (
    .a(ds1[50]),
    .b(\exu/alu_au/n17 [50]),
    .c(\exu/alu_au/add0/c50 ),
    .o({\exu/alu_au/add0/c51 ,\exu/alu_au/add_64 [50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u51  (
    .a(ds1[51]),
    .b(\exu/alu_au/n17 [51]),
    .c(\exu/alu_au/add0/c51 ),
    .o({\exu/alu_au/add0/c52 ,\exu/alu_au/add_64 [51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u52  (
    .a(ds1[52]),
    .b(\exu/alu_au/n17 [52]),
    .c(\exu/alu_au/add0/c52 ),
    .o({\exu/alu_au/add0/c53 ,\exu/alu_au/add_64 [52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u53  (
    .a(ds1[53]),
    .b(\exu/alu_au/n17 [53]),
    .c(\exu/alu_au/add0/c53 ),
    .o({\exu/alu_au/add0/c54 ,\exu/alu_au/add_64 [53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u54  (
    .a(ds1[54]),
    .b(\exu/alu_au/n17 [54]),
    .c(\exu/alu_au/add0/c54 ),
    .o({\exu/alu_au/add0/c55 ,\exu/alu_au/add_64 [54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u55  (
    .a(ds1[55]),
    .b(\exu/alu_au/n17 [55]),
    .c(\exu/alu_au/add0/c55 ),
    .o({\exu/alu_au/add0/c56 ,\exu/alu_au/add_64 [55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u56  (
    .a(ds1[56]),
    .b(\exu/alu_au/n17 [56]),
    .c(\exu/alu_au/add0/c56 ),
    .o({\exu/alu_au/add0/c57 ,\exu/alu_au/add_64 [56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u57  (
    .a(ds1[57]),
    .b(\exu/alu_au/n17 [57]),
    .c(\exu/alu_au/add0/c57 ),
    .o({\exu/alu_au/add0/c58 ,\exu/alu_au/add_64 [57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u58  (
    .a(ds1[58]),
    .b(\exu/alu_au/n17 [58]),
    .c(\exu/alu_au/add0/c58 ),
    .o({\exu/alu_au/add0/c59 ,\exu/alu_au/add_64 [58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u59  (
    .a(ds1[59]),
    .b(\exu/alu_au/n17 [59]),
    .c(\exu/alu_au/add0/c59 ),
    .o({\exu/alu_au/add0/c60 ,\exu/alu_au/add_64 [59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u6  (
    .a(ds1[6]),
    .b(\exu/alu_au/n17 [6]),
    .c(\exu/alu_au/add0/c6 ),
    .o({\exu/alu_au/add0/c7 ,\exu/alu_au/add_64 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u60  (
    .a(ds1[60]),
    .b(\exu/alu_au/n17 [60]),
    .c(\exu/alu_au/add0/c60 ),
    .o({\exu/alu_au/add0/c61 ,\exu/alu_au/add_64 [60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u61  (
    .a(ds1[61]),
    .b(\exu/alu_au/n17 [61]),
    .c(\exu/alu_au/add0/c61 ),
    .o({\exu/alu_au/add0/c62 ,\exu/alu_au/add_64 [61]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u62  (
    .a(ds1[62]),
    .b(\exu/alu_au/n17 [62]),
    .c(\exu/alu_au/add0/c62 ),
    .o({\exu/alu_au/add0/c63 ,\exu/alu_au/add_64 [62]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u63  (
    .a(ds1[63]),
    .b(\exu/alu_au/n17 [63]),
    .c(\exu/alu_au/add0/c63 ),
    .o({open_n6132,\exu/alu_au/add_64 [63]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u7  (
    .a(ds1[7]),
    .b(\exu/alu_au/n17 [7]),
    .c(\exu/alu_au/add0/c7 ),
    .o({\exu/alu_au/add0/c8 ,\exu/alu_au/add_64 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u8  (
    .a(ds1[8]),
    .b(\exu/alu_au/n17 [8]),
    .c(\exu/alu_au/add0/c8 ),
    .o({\exu/alu_au/add0/c9 ,\exu/alu_au/add_64 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add0/u9  (
    .a(ds1[9]),
    .b(\exu/alu_au/n17 [9]),
    .c(\exu/alu_au/add0/c9 ),
    .o({\exu/alu_au/add0/c10 ,\exu/alu_au/add_64 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \exu/alu_au/add0/ucin  (
    .a(1'b0),
    .o({\exu/alu_au/add0/c0 ,open_n6135}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u0  (
    .a(\exu/alu_au/add_64 [0]),
    .b(1'b1),
    .c(\exu/alu_au/add1/c0 ),
    .o({\exu/alu_au/add1/c1 ,\exu/alu_au/sub_64 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u1  (
    .a(\exu/alu_au/add_64 [1]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c1 ),
    .o({\exu/alu_au/add1/c2 ,\exu/alu_au/sub_64 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u10  (
    .a(\exu/alu_au/add_64 [10]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c10 ),
    .o({\exu/alu_au/add1/c11 ,\exu/alu_au/sub_64 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u11  (
    .a(\exu/alu_au/add_64 [11]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c11 ),
    .o({\exu/alu_au/add1/c12 ,\exu/alu_au/sub_64 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u12  (
    .a(\exu/alu_au/add_64 [12]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c12 ),
    .o({\exu/alu_au/add1/c13 ,\exu/alu_au/sub_64 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u13  (
    .a(\exu/alu_au/add_64 [13]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c13 ),
    .o({\exu/alu_au/add1/c14 ,\exu/alu_au/sub_64 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u14  (
    .a(\exu/alu_au/add_64 [14]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c14 ),
    .o({\exu/alu_au/add1/c15 ,\exu/alu_au/sub_64 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u15  (
    .a(\exu/alu_au/add_64 [15]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c15 ),
    .o({\exu/alu_au/add1/c16 ,\exu/alu_au/sub_64 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u16  (
    .a(\exu/alu_au/add_64 [16]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c16 ),
    .o({\exu/alu_au/add1/c17 ,\exu/alu_au/sub_64 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u17  (
    .a(\exu/alu_au/add_64 [17]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c17 ),
    .o({\exu/alu_au/add1/c18 ,\exu/alu_au/sub_64 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u18  (
    .a(\exu/alu_au/add_64 [18]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c18 ),
    .o({\exu/alu_au/add1/c19 ,\exu/alu_au/sub_64 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u19  (
    .a(\exu/alu_au/add_64 [19]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c19 ),
    .o({\exu/alu_au/add1/c20 ,\exu/alu_au/sub_64 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u2  (
    .a(\exu/alu_au/add_64 [2]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c2 ),
    .o({\exu/alu_au/add1/c3 ,\exu/alu_au/sub_64 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u20  (
    .a(\exu/alu_au/add_64 [20]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c20 ),
    .o({\exu/alu_au/add1/c21 ,\exu/alu_au/sub_64 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u21  (
    .a(\exu/alu_au/add_64 [21]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c21 ),
    .o({\exu/alu_au/add1/c22 ,\exu/alu_au/sub_64 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u22  (
    .a(\exu/alu_au/add_64 [22]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c22 ),
    .o({\exu/alu_au/add1/c23 ,\exu/alu_au/sub_64 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u23  (
    .a(\exu/alu_au/add_64 [23]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c23 ),
    .o({\exu/alu_au/add1/c24 ,\exu/alu_au/sub_64 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u24  (
    .a(\exu/alu_au/add_64 [24]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c24 ),
    .o({\exu/alu_au/add1/c25 ,\exu/alu_au/sub_64 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u25  (
    .a(\exu/alu_au/add_64 [25]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c25 ),
    .o({\exu/alu_au/add1/c26 ,\exu/alu_au/sub_64 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u26  (
    .a(\exu/alu_au/add_64 [26]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c26 ),
    .o({\exu/alu_au/add1/c27 ,\exu/alu_au/sub_64 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u27  (
    .a(\exu/alu_au/add_64 [27]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c27 ),
    .o({\exu/alu_au/add1/c28 ,\exu/alu_au/sub_64 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u28  (
    .a(\exu/alu_au/add_64 [28]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c28 ),
    .o({\exu/alu_au/add1/c29 ,\exu/alu_au/sub_64 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u29  (
    .a(\exu/alu_au/add_64 [29]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c29 ),
    .o({\exu/alu_au/add1/c30 ,\exu/alu_au/sub_64 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u3  (
    .a(\exu/alu_au/add_64 [3]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c3 ),
    .o({\exu/alu_au/add1/c4 ,\exu/alu_au/sub_64 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u30  (
    .a(\exu/alu_au/add_64 [30]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c30 ),
    .o({\exu/alu_au/add1/c31 ,\exu/alu_au/sub_64 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u31  (
    .a(\exu/alu_au/add_64 [31]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c31 ),
    .o({open_n6136,\exu/alu_au/sub_64 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u4  (
    .a(\exu/alu_au/add_64 [4]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c4 ),
    .o({\exu/alu_au/add1/c5 ,\exu/alu_au/sub_64 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u5  (
    .a(\exu/alu_au/add_64 [5]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c5 ),
    .o({\exu/alu_au/add1/c6 ,\exu/alu_au/sub_64 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u6  (
    .a(\exu/alu_au/add_64 [6]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c6 ),
    .o({\exu/alu_au/add1/c7 ,\exu/alu_au/sub_64 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u7  (
    .a(\exu/alu_au/add_64 [7]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c7 ),
    .o({\exu/alu_au/add1/c8 ,\exu/alu_au/sub_64 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u8  (
    .a(\exu/alu_au/add_64 [8]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c8 ),
    .o({\exu/alu_au/add1/c9 ,\exu/alu_au/sub_64 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add1/u9  (
    .a(\exu/alu_au/add_64 [9]),
    .b(1'b0),
    .c(\exu/alu_au/add1/c9 ),
    .o({\exu/alu_au/add1/c10 ,\exu/alu_au/sub_64 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \exu/alu_au/add1/ucin  (
    .a(1'b0),
    .o({\exu/alu_au/add1/c0 ,open_n6139}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u0  (
    .a(as1[0]),
    .b(as2[0]),
    .c(\exu/alu_au/add2/c0 ),
    .o({\exu/alu_au/add2/c1 ,addr_ex[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u1  (
    .a(as1[1]),
    .b(as2[1]),
    .c(\exu/alu_au/add2/c1 ),
    .o({\exu/alu_au/add2/c2 ,addr_ex[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u10  (
    .a(as1[10]),
    .b(as2[10]),
    .c(\exu/alu_au/add2/c10 ),
    .o({\exu/alu_au/add2/c11 ,addr_ex[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u11  (
    .a(as1[11]),
    .b(as2[11]),
    .c(\exu/alu_au/add2/c11 ),
    .o({\exu/alu_au/add2/c12 ,addr_ex[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u12  (
    .a(as1[12]),
    .b(as2[12]),
    .c(\exu/alu_au/add2/c12 ),
    .o({\exu/alu_au/add2/c13 ,addr_ex[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u13  (
    .a(as1[13]),
    .b(as2[13]),
    .c(\exu/alu_au/add2/c13 ),
    .o({\exu/alu_au/add2/c14 ,addr_ex[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u14  (
    .a(as1[14]),
    .b(as2[14]),
    .c(\exu/alu_au/add2/c14 ),
    .o({\exu/alu_au/add2/c15 ,addr_ex[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u15  (
    .a(as1[15]),
    .b(as2[15]),
    .c(\exu/alu_au/add2/c15 ),
    .o({\exu/alu_au/add2/c16 ,addr_ex[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u16  (
    .a(as1[16]),
    .b(as2[16]),
    .c(\exu/alu_au/add2/c16 ),
    .o({\exu/alu_au/add2/c17 ,addr_ex[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u17  (
    .a(as1[17]),
    .b(as2[17]),
    .c(\exu/alu_au/add2/c17 ),
    .o({\exu/alu_au/add2/c18 ,addr_ex[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u18  (
    .a(as1[18]),
    .b(as2[18]),
    .c(\exu/alu_au/add2/c18 ),
    .o({\exu/alu_au/add2/c19 ,addr_ex[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u19  (
    .a(as1[19]),
    .b(as2[19]),
    .c(\exu/alu_au/add2/c19 ),
    .o({\exu/alu_au/add2/c20 ,addr_ex[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u2  (
    .a(as1[2]),
    .b(as2[2]),
    .c(\exu/alu_au/add2/c2 ),
    .o({\exu/alu_au/add2/c3 ,addr_ex[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u20  (
    .a(as1[20]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c20 ),
    .o({\exu/alu_au/add2/c21 ,addr_ex[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u21  (
    .a(as1[21]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c21 ),
    .o({\exu/alu_au/add2/c22 ,addr_ex[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u22  (
    .a(as1[22]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c22 ),
    .o({\exu/alu_au/add2/c23 ,addr_ex[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u23  (
    .a(as1[23]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c23 ),
    .o({\exu/alu_au/add2/c24 ,addr_ex[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u24  (
    .a(as1[24]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c24 ),
    .o({\exu/alu_au/add2/c25 ,addr_ex[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u25  (
    .a(as1[25]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c25 ),
    .o({\exu/alu_au/add2/c26 ,addr_ex[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u26  (
    .a(as1[26]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c26 ),
    .o({\exu/alu_au/add2/c27 ,addr_ex[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u27  (
    .a(as1[27]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c27 ),
    .o({\exu/alu_au/add2/c28 ,addr_ex[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u28  (
    .a(as1[28]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c28 ),
    .o({\exu/alu_au/add2/c29 ,addr_ex[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u29  (
    .a(as1[29]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c29 ),
    .o({\exu/alu_au/add2/c30 ,addr_ex[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u3  (
    .a(as1[3]),
    .b(as2[3]),
    .c(\exu/alu_au/add2/c3 ),
    .o({\exu/alu_au/add2/c4 ,addr_ex[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u30  (
    .a(as1[30]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c30 ),
    .o({\exu/alu_au/add2/c31 ,addr_ex[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u31  (
    .a(as1[31]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c31 ),
    .o({\exu/alu_au/add2/c32 ,addr_ex[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u32  (
    .a(as1[32]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c32 ),
    .o({\exu/alu_au/add2/c33 ,addr_ex[32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u33  (
    .a(as1[33]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c33 ),
    .o({\exu/alu_au/add2/c34 ,addr_ex[33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u34  (
    .a(as1[34]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c34 ),
    .o({\exu/alu_au/add2/c35 ,addr_ex[34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u35  (
    .a(as1[35]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c35 ),
    .o({\exu/alu_au/add2/c36 ,addr_ex[35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u36  (
    .a(as1[36]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c36 ),
    .o({\exu/alu_au/add2/c37 ,addr_ex[36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u37  (
    .a(as1[37]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c37 ),
    .o({\exu/alu_au/add2/c38 ,addr_ex[37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u38  (
    .a(as1[38]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c38 ),
    .o({\exu/alu_au/add2/c39 ,addr_ex[38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u39  (
    .a(as1[39]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c39 ),
    .o({\exu/alu_au/add2/c40 ,addr_ex[39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u4  (
    .a(as1[4]),
    .b(as2[4]),
    .c(\exu/alu_au/add2/c4 ),
    .o({\exu/alu_au/add2/c5 ,addr_ex[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u40  (
    .a(as1[40]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c40 ),
    .o({\exu/alu_au/add2/c41 ,addr_ex[40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u41  (
    .a(as1[41]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c41 ),
    .o({\exu/alu_au/add2/c42 ,addr_ex[41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u42  (
    .a(as1[42]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c42 ),
    .o({\exu/alu_au/add2/c43 ,addr_ex[42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u43  (
    .a(as1[43]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c43 ),
    .o({\exu/alu_au/add2/c44 ,addr_ex[43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u44  (
    .a(as1[44]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c44 ),
    .o({\exu/alu_au/add2/c45 ,addr_ex[44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u45  (
    .a(as1[45]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c45 ),
    .o({\exu/alu_au/add2/c46 ,addr_ex[45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u46  (
    .a(as1[46]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c46 ),
    .o({\exu/alu_au/add2/c47 ,addr_ex[46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u47  (
    .a(as1[47]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c47 ),
    .o({\exu/alu_au/add2/c48 ,addr_ex[47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u48  (
    .a(as1[48]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c48 ),
    .o({\exu/alu_au/add2/c49 ,addr_ex[48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u49  (
    .a(as1[49]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c49 ),
    .o({\exu/alu_au/add2/c50 ,addr_ex[49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u5  (
    .a(as1[5]),
    .b(as2[5]),
    .c(\exu/alu_au/add2/c5 ),
    .o({\exu/alu_au/add2/c6 ,addr_ex[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u50  (
    .a(as1[50]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c50 ),
    .o({\exu/alu_au/add2/c51 ,addr_ex[50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u51  (
    .a(as1[51]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c51 ),
    .o({\exu/alu_au/add2/c52 ,addr_ex[51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u52  (
    .a(as1[52]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c52 ),
    .o({\exu/alu_au/add2/c53 ,addr_ex[52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u53  (
    .a(as1[53]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c53 ),
    .o({\exu/alu_au/add2/c54 ,addr_ex[53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u54  (
    .a(as1[54]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c54 ),
    .o({\exu/alu_au/add2/c55 ,addr_ex[54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u55  (
    .a(as1[55]),
    .b(as2[20]),
    .c(\exu/alu_au/add2/c55 ),
    .o({\exu/alu_au/add2/c56 ,addr_ex[55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u56  (
    .a(as1[56]),
    .b(as2[56]),
    .c(\exu/alu_au/add2/c56 ),
    .o({\exu/alu_au/add2/c57 ,addr_ex[56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u57  (
    .a(as1[57]),
    .b(as2[56]),
    .c(\exu/alu_au/add2/c57 ),
    .o({\exu/alu_au/add2/c58 ,addr_ex[57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u58  (
    .a(as1[58]),
    .b(as2[56]),
    .c(\exu/alu_au/add2/c58 ),
    .o({\exu/alu_au/add2/c59 ,addr_ex[58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u59  (
    .a(as1[59]),
    .b(as2[56]),
    .c(\exu/alu_au/add2/c59 ),
    .o({\exu/alu_au/add2/c60 ,addr_ex[59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u6  (
    .a(as1[6]),
    .b(as2[6]),
    .c(\exu/alu_au/add2/c6 ),
    .o({\exu/alu_au/add2/c7 ,addr_ex[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u60  (
    .a(as1[60]),
    .b(as2[56]),
    .c(\exu/alu_au/add2/c60 ),
    .o({\exu/alu_au/add2/c61 ,addr_ex[60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u61  (
    .a(as1[61]),
    .b(as2[56]),
    .c(\exu/alu_au/add2/c61 ),
    .o({\exu/alu_au/add2/c62 ,addr_ex[61]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u62  (
    .a(as1[62]),
    .b(as2[56]),
    .c(\exu/alu_au/add2/c62 ),
    .o({\exu/alu_au/add2/c63 ,addr_ex[62]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u63  (
    .a(as1[63]),
    .b(as2[56]),
    .c(\exu/alu_au/add2/c63 ),
    .o({open_n6140,addr_ex[63]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u7  (
    .a(as1[7]),
    .b(as2[7]),
    .c(\exu/alu_au/add2/c7 ),
    .o({\exu/alu_au/add2/c8 ,addr_ex[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u8  (
    .a(as1[8]),
    .b(as2[8]),
    .c(\exu/alu_au/add2/c8 ),
    .o({\exu/alu_au/add2/c9 ,addr_ex[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \exu/alu_au/add2/u9  (
    .a(as1[9]),
    .b(as2[9]),
    .c(\exu/alu_au/add2/c9 ),
    .o({\exu/alu_au/add2/c10 ,addr_ex[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \exu/alu_au/add2/ucin  (
    .a(1'b0),
    .o({\exu/alu_au/add2/c0 ,open_n6143}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_0  (
    .a(ds1[0]),
    .b(ds2[0]),
    .c(\exu/alu_au/lt0_c0 ),
    .o({\exu/alu_au/lt0_c1 ,open_n6144}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_1  (
    .a(ds1[1]),
    .b(ds2[1]),
    .c(\exu/alu_au/lt0_c1 ),
    .o({\exu/alu_au/lt0_c2 ,open_n6145}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_10  (
    .a(ds1[10]),
    .b(ds2[10]),
    .c(\exu/alu_au/lt0_c10 ),
    .o({\exu/alu_au/lt0_c11 ,open_n6146}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_11  (
    .a(ds1[11]),
    .b(ds2[11]),
    .c(\exu/alu_au/lt0_c11 ),
    .o({\exu/alu_au/lt0_c12 ,open_n6147}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_12  (
    .a(ds1[12]),
    .b(ds2[12]),
    .c(\exu/alu_au/lt0_c12 ),
    .o({\exu/alu_au/lt0_c13 ,open_n6148}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_13  (
    .a(ds1[13]),
    .b(ds2[13]),
    .c(\exu/alu_au/lt0_c13 ),
    .o({\exu/alu_au/lt0_c14 ,open_n6149}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_14  (
    .a(ds1[14]),
    .b(ds2[14]),
    .c(\exu/alu_au/lt0_c14 ),
    .o({\exu/alu_au/lt0_c15 ,open_n6150}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_15  (
    .a(ds1[15]),
    .b(ds2[15]),
    .c(\exu/alu_au/lt0_c15 ),
    .o({\exu/alu_au/lt0_c16 ,open_n6151}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_16  (
    .a(ds1[16]),
    .b(ds2[16]),
    .c(\exu/alu_au/lt0_c16 ),
    .o({\exu/alu_au/lt0_c17 ,open_n6152}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_17  (
    .a(ds1[17]),
    .b(ds2[17]),
    .c(\exu/alu_au/lt0_c17 ),
    .o({\exu/alu_au/lt0_c18 ,open_n6153}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_18  (
    .a(ds1[18]),
    .b(ds2[18]),
    .c(\exu/alu_au/lt0_c18 ),
    .o({\exu/alu_au/lt0_c19 ,open_n6154}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_19  (
    .a(ds1[19]),
    .b(ds2[19]),
    .c(\exu/alu_au/lt0_c19 ),
    .o({\exu/alu_au/lt0_c20 ,open_n6155}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_2  (
    .a(ds1[2]),
    .b(ds2[2]),
    .c(\exu/alu_au/lt0_c2 ),
    .o({\exu/alu_au/lt0_c3 ,open_n6156}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_20  (
    .a(ds1[20]),
    .b(ds2[20]),
    .c(\exu/alu_au/lt0_c20 ),
    .o({\exu/alu_au/lt0_c21 ,open_n6157}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_21  (
    .a(ds1[21]),
    .b(ds2[21]),
    .c(\exu/alu_au/lt0_c21 ),
    .o({\exu/alu_au/lt0_c22 ,open_n6158}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_22  (
    .a(ds1[22]),
    .b(ds2[22]),
    .c(\exu/alu_au/lt0_c22 ),
    .o({\exu/alu_au/lt0_c23 ,open_n6159}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_23  (
    .a(ds1[23]),
    .b(ds2[23]),
    .c(\exu/alu_au/lt0_c23 ),
    .o({\exu/alu_au/lt0_c24 ,open_n6160}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_24  (
    .a(ds1[24]),
    .b(ds2[24]),
    .c(\exu/alu_au/lt0_c24 ),
    .o({\exu/alu_au/lt0_c25 ,open_n6161}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_25  (
    .a(ds1[25]),
    .b(ds2[25]),
    .c(\exu/alu_au/lt0_c25 ),
    .o({\exu/alu_au/lt0_c26 ,open_n6162}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_26  (
    .a(ds1[26]),
    .b(ds2[26]),
    .c(\exu/alu_au/lt0_c26 ),
    .o({\exu/alu_au/lt0_c27 ,open_n6163}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_27  (
    .a(ds1[27]),
    .b(ds2[27]),
    .c(\exu/alu_au/lt0_c27 ),
    .o({\exu/alu_au/lt0_c28 ,open_n6164}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_28  (
    .a(ds1[28]),
    .b(ds2[28]),
    .c(\exu/alu_au/lt0_c28 ),
    .o({\exu/alu_au/lt0_c29 ,open_n6165}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_29  (
    .a(ds1[29]),
    .b(ds2[29]),
    .c(\exu/alu_au/lt0_c29 ),
    .o({\exu/alu_au/lt0_c30 ,open_n6166}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_3  (
    .a(ds1[3]),
    .b(ds2[3]),
    .c(\exu/alu_au/lt0_c3 ),
    .o({\exu/alu_au/lt0_c4 ,open_n6167}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_30  (
    .a(ds1[30]),
    .b(ds2[30]),
    .c(\exu/alu_au/lt0_c30 ),
    .o({\exu/alu_au/lt0_c31 ,open_n6168}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_31  (
    .a(ds1[31]),
    .b(ds2[31]),
    .c(\exu/alu_au/lt0_c31 ),
    .o({\exu/alu_au/lt0_c32 ,open_n6169}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_32  (
    .a(ds1[32]),
    .b(ds2[32]),
    .c(\exu/alu_au/lt0_c32 ),
    .o({\exu/alu_au/lt0_c33 ,open_n6170}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_33  (
    .a(ds1[33]),
    .b(ds2[33]),
    .c(\exu/alu_au/lt0_c33 ),
    .o({\exu/alu_au/lt0_c34 ,open_n6171}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_34  (
    .a(ds1[34]),
    .b(ds2[34]),
    .c(\exu/alu_au/lt0_c34 ),
    .o({\exu/alu_au/lt0_c35 ,open_n6172}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_35  (
    .a(ds1[35]),
    .b(ds2[35]),
    .c(\exu/alu_au/lt0_c35 ),
    .o({\exu/alu_au/lt0_c36 ,open_n6173}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_36  (
    .a(ds1[36]),
    .b(ds2[36]),
    .c(\exu/alu_au/lt0_c36 ),
    .o({\exu/alu_au/lt0_c37 ,open_n6174}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_37  (
    .a(ds1[37]),
    .b(ds2[37]),
    .c(\exu/alu_au/lt0_c37 ),
    .o({\exu/alu_au/lt0_c38 ,open_n6175}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_38  (
    .a(ds1[38]),
    .b(ds2[38]),
    .c(\exu/alu_au/lt0_c38 ),
    .o({\exu/alu_au/lt0_c39 ,open_n6176}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_39  (
    .a(ds1[39]),
    .b(ds2[39]),
    .c(\exu/alu_au/lt0_c39 ),
    .o({\exu/alu_au/lt0_c40 ,open_n6177}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_4  (
    .a(ds1[4]),
    .b(ds2[4]),
    .c(\exu/alu_au/lt0_c4 ),
    .o({\exu/alu_au/lt0_c5 ,open_n6178}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_40  (
    .a(ds1[40]),
    .b(ds2[40]),
    .c(\exu/alu_au/lt0_c40 ),
    .o({\exu/alu_au/lt0_c41 ,open_n6179}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_41  (
    .a(ds1[41]),
    .b(ds2[41]),
    .c(\exu/alu_au/lt0_c41 ),
    .o({\exu/alu_au/lt0_c42 ,open_n6180}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_42  (
    .a(ds1[42]),
    .b(ds2[42]),
    .c(\exu/alu_au/lt0_c42 ),
    .o({\exu/alu_au/lt0_c43 ,open_n6181}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_43  (
    .a(ds1[43]),
    .b(ds2[43]),
    .c(\exu/alu_au/lt0_c43 ),
    .o({\exu/alu_au/lt0_c44 ,open_n6182}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_44  (
    .a(ds1[44]),
    .b(ds2[44]),
    .c(\exu/alu_au/lt0_c44 ),
    .o({\exu/alu_au/lt0_c45 ,open_n6183}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_45  (
    .a(ds1[45]),
    .b(ds2[45]),
    .c(\exu/alu_au/lt0_c45 ),
    .o({\exu/alu_au/lt0_c46 ,open_n6184}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_46  (
    .a(ds1[46]),
    .b(ds2[46]),
    .c(\exu/alu_au/lt0_c46 ),
    .o({\exu/alu_au/lt0_c47 ,open_n6185}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_47  (
    .a(ds1[47]),
    .b(ds2[47]),
    .c(\exu/alu_au/lt0_c47 ),
    .o({\exu/alu_au/lt0_c48 ,open_n6186}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_48  (
    .a(ds1[48]),
    .b(ds2[48]),
    .c(\exu/alu_au/lt0_c48 ),
    .o({\exu/alu_au/lt0_c49 ,open_n6187}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_49  (
    .a(ds1[49]),
    .b(ds2[49]),
    .c(\exu/alu_au/lt0_c49 ),
    .o({\exu/alu_au/lt0_c50 ,open_n6188}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_5  (
    .a(ds1[5]),
    .b(ds2[5]),
    .c(\exu/alu_au/lt0_c5 ),
    .o({\exu/alu_au/lt0_c6 ,open_n6189}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_50  (
    .a(ds1[50]),
    .b(ds2[50]),
    .c(\exu/alu_au/lt0_c50 ),
    .o({\exu/alu_au/lt0_c51 ,open_n6190}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_51  (
    .a(ds1[51]),
    .b(ds2[51]),
    .c(\exu/alu_au/lt0_c51 ),
    .o({\exu/alu_au/lt0_c52 ,open_n6191}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_52  (
    .a(ds1[52]),
    .b(ds2[52]),
    .c(\exu/alu_au/lt0_c52 ),
    .o({\exu/alu_au/lt0_c53 ,open_n6192}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_53  (
    .a(ds1[53]),
    .b(ds2[53]),
    .c(\exu/alu_au/lt0_c53 ),
    .o({\exu/alu_au/lt0_c54 ,open_n6193}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_54  (
    .a(ds1[54]),
    .b(ds2[54]),
    .c(\exu/alu_au/lt0_c54 ),
    .o({\exu/alu_au/lt0_c55 ,open_n6194}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_55  (
    .a(ds1[55]),
    .b(ds2[55]),
    .c(\exu/alu_au/lt0_c55 ),
    .o({\exu/alu_au/lt0_c56 ,open_n6195}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_56  (
    .a(ds1[56]),
    .b(ds2[56]),
    .c(\exu/alu_au/lt0_c56 ),
    .o({\exu/alu_au/lt0_c57 ,open_n6196}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_57  (
    .a(ds1[57]),
    .b(ds2[57]),
    .c(\exu/alu_au/lt0_c57 ),
    .o({\exu/alu_au/lt0_c58 ,open_n6197}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_58  (
    .a(ds1[58]),
    .b(ds2[58]),
    .c(\exu/alu_au/lt0_c58 ),
    .o({\exu/alu_au/lt0_c59 ,open_n6198}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_59  (
    .a(ds1[59]),
    .b(ds2[59]),
    .c(\exu/alu_au/lt0_c59 ),
    .o({\exu/alu_au/lt0_c60 ,open_n6199}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_6  (
    .a(ds1[6]),
    .b(ds2[6]),
    .c(\exu/alu_au/lt0_c6 ),
    .o({\exu/alu_au/lt0_c7 ,open_n6200}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_60  (
    .a(ds1[60]),
    .b(ds2[60]),
    .c(\exu/alu_au/lt0_c60 ),
    .o({\exu/alu_au/lt0_c61 ,open_n6201}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_61  (
    .a(ds1[61]),
    .b(ds2[61]),
    .c(\exu/alu_au/lt0_c61 ),
    .o({\exu/alu_au/lt0_c62 ,open_n6202}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_62  (
    .a(ds1[62]),
    .b(ds2[62]),
    .c(\exu/alu_au/lt0_c62 ),
    .o({\exu/alu_au/lt0_c63 ,open_n6203}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_63  (
    .a(ds1[63]),
    .b(ds2[63]),
    .c(\exu/alu_au/lt0_c63 ),
    .o({\exu/alu_au/lt0_c64 ,open_n6204}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_7  (
    .a(ds1[7]),
    .b(ds2[7]),
    .c(\exu/alu_au/lt0_c7 ),
    .o({\exu/alu_au/lt0_c8 ,open_n6205}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_8  (
    .a(ds1[8]),
    .b(ds2[8]),
    .c(\exu/alu_au/lt0_c8 ),
    .o({\exu/alu_au/lt0_c9 ,open_n6206}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_9  (
    .a(ds1[9]),
    .b(ds2[9]),
    .c(\exu/alu_au/lt0_c9 ),
    .o({\exu/alu_au/lt0_c10 ,open_n6207}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \exu/alu_au/lt0_cin  (
    .a(1'b0),
    .o({\exu/alu_au/lt0_c0 ,open_n6210}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt0_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\exu/alu_au/lt0_c64 ),
    .o({open_n6211,\exu/alu_au/n5 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_0  (
    .a(ds2[0]),
    .b(ds1[0]),
    .c(\exu/alu_au/lt1_c0 ),
    .o({\exu/alu_au/lt1_c1 ,open_n6212}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_1  (
    .a(ds2[1]),
    .b(ds1[1]),
    .c(\exu/alu_au/lt1_c1 ),
    .o({\exu/alu_au/lt1_c2 ,open_n6213}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_10  (
    .a(ds2[10]),
    .b(ds1[10]),
    .c(\exu/alu_au/lt1_c10 ),
    .o({\exu/alu_au/lt1_c11 ,open_n6214}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_11  (
    .a(ds2[11]),
    .b(ds1[11]),
    .c(\exu/alu_au/lt1_c11 ),
    .o({\exu/alu_au/lt1_c12 ,open_n6215}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_12  (
    .a(ds2[12]),
    .b(ds1[12]),
    .c(\exu/alu_au/lt1_c12 ),
    .o({\exu/alu_au/lt1_c13 ,open_n6216}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_13  (
    .a(ds2[13]),
    .b(ds1[13]),
    .c(\exu/alu_au/lt1_c13 ),
    .o({\exu/alu_au/lt1_c14 ,open_n6217}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_14  (
    .a(ds2[14]),
    .b(ds1[14]),
    .c(\exu/alu_au/lt1_c14 ),
    .o({\exu/alu_au/lt1_c15 ,open_n6218}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_15  (
    .a(ds2[15]),
    .b(ds1[15]),
    .c(\exu/alu_au/lt1_c15 ),
    .o({\exu/alu_au/lt1_c16 ,open_n6219}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_16  (
    .a(ds2[16]),
    .b(ds1[16]),
    .c(\exu/alu_au/lt1_c16 ),
    .o({\exu/alu_au/lt1_c17 ,open_n6220}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_17  (
    .a(ds2[17]),
    .b(ds1[17]),
    .c(\exu/alu_au/lt1_c17 ),
    .o({\exu/alu_au/lt1_c18 ,open_n6221}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_18  (
    .a(ds2[18]),
    .b(ds1[18]),
    .c(\exu/alu_au/lt1_c18 ),
    .o({\exu/alu_au/lt1_c19 ,open_n6222}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_19  (
    .a(ds2[19]),
    .b(ds1[19]),
    .c(\exu/alu_au/lt1_c19 ),
    .o({\exu/alu_au/lt1_c20 ,open_n6223}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_2  (
    .a(ds2[2]),
    .b(ds1[2]),
    .c(\exu/alu_au/lt1_c2 ),
    .o({\exu/alu_au/lt1_c3 ,open_n6224}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_20  (
    .a(ds2[20]),
    .b(ds1[20]),
    .c(\exu/alu_au/lt1_c20 ),
    .o({\exu/alu_au/lt1_c21 ,open_n6225}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_21  (
    .a(ds2[21]),
    .b(ds1[21]),
    .c(\exu/alu_au/lt1_c21 ),
    .o({\exu/alu_au/lt1_c22 ,open_n6226}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_22  (
    .a(ds2[22]),
    .b(ds1[22]),
    .c(\exu/alu_au/lt1_c22 ),
    .o({\exu/alu_au/lt1_c23 ,open_n6227}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_23  (
    .a(ds2[23]),
    .b(ds1[23]),
    .c(\exu/alu_au/lt1_c23 ),
    .o({\exu/alu_au/lt1_c24 ,open_n6228}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_24  (
    .a(ds2[24]),
    .b(ds1[24]),
    .c(\exu/alu_au/lt1_c24 ),
    .o({\exu/alu_au/lt1_c25 ,open_n6229}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_25  (
    .a(ds2[25]),
    .b(ds1[25]),
    .c(\exu/alu_au/lt1_c25 ),
    .o({\exu/alu_au/lt1_c26 ,open_n6230}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_26  (
    .a(ds2[26]),
    .b(ds1[26]),
    .c(\exu/alu_au/lt1_c26 ),
    .o({\exu/alu_au/lt1_c27 ,open_n6231}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_27  (
    .a(ds2[27]),
    .b(ds1[27]),
    .c(\exu/alu_au/lt1_c27 ),
    .o({\exu/alu_au/lt1_c28 ,open_n6232}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_28  (
    .a(ds2[28]),
    .b(ds1[28]),
    .c(\exu/alu_au/lt1_c28 ),
    .o({\exu/alu_au/lt1_c29 ,open_n6233}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_29  (
    .a(ds2[29]),
    .b(ds1[29]),
    .c(\exu/alu_au/lt1_c29 ),
    .o({\exu/alu_au/lt1_c30 ,open_n6234}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_3  (
    .a(ds2[3]),
    .b(ds1[3]),
    .c(\exu/alu_au/lt1_c3 ),
    .o({\exu/alu_au/lt1_c4 ,open_n6235}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_30  (
    .a(ds2[30]),
    .b(ds1[30]),
    .c(\exu/alu_au/lt1_c30 ),
    .o({\exu/alu_au/lt1_c31 ,open_n6236}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_31  (
    .a(ds2[31]),
    .b(ds1[31]),
    .c(\exu/alu_au/lt1_c31 ),
    .o({\exu/alu_au/lt1_c32 ,open_n6237}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_32  (
    .a(ds2[32]),
    .b(ds1[32]),
    .c(\exu/alu_au/lt1_c32 ),
    .o({\exu/alu_au/lt1_c33 ,open_n6238}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_33  (
    .a(ds2[33]),
    .b(ds1[33]),
    .c(\exu/alu_au/lt1_c33 ),
    .o({\exu/alu_au/lt1_c34 ,open_n6239}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_34  (
    .a(ds2[34]),
    .b(ds1[34]),
    .c(\exu/alu_au/lt1_c34 ),
    .o({\exu/alu_au/lt1_c35 ,open_n6240}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_35  (
    .a(ds2[35]),
    .b(ds1[35]),
    .c(\exu/alu_au/lt1_c35 ),
    .o({\exu/alu_au/lt1_c36 ,open_n6241}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_36  (
    .a(ds2[36]),
    .b(ds1[36]),
    .c(\exu/alu_au/lt1_c36 ),
    .o({\exu/alu_au/lt1_c37 ,open_n6242}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_37  (
    .a(ds2[37]),
    .b(ds1[37]),
    .c(\exu/alu_au/lt1_c37 ),
    .o({\exu/alu_au/lt1_c38 ,open_n6243}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_38  (
    .a(ds2[38]),
    .b(ds1[38]),
    .c(\exu/alu_au/lt1_c38 ),
    .o({\exu/alu_au/lt1_c39 ,open_n6244}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_39  (
    .a(ds2[39]),
    .b(ds1[39]),
    .c(\exu/alu_au/lt1_c39 ),
    .o({\exu/alu_au/lt1_c40 ,open_n6245}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_4  (
    .a(ds2[4]),
    .b(ds1[4]),
    .c(\exu/alu_au/lt1_c4 ),
    .o({\exu/alu_au/lt1_c5 ,open_n6246}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_40  (
    .a(ds2[40]),
    .b(ds1[40]),
    .c(\exu/alu_au/lt1_c40 ),
    .o({\exu/alu_au/lt1_c41 ,open_n6247}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_41  (
    .a(ds2[41]),
    .b(ds1[41]),
    .c(\exu/alu_au/lt1_c41 ),
    .o({\exu/alu_au/lt1_c42 ,open_n6248}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_42  (
    .a(ds2[42]),
    .b(ds1[42]),
    .c(\exu/alu_au/lt1_c42 ),
    .o({\exu/alu_au/lt1_c43 ,open_n6249}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_43  (
    .a(ds2[43]),
    .b(ds1[43]),
    .c(\exu/alu_au/lt1_c43 ),
    .o({\exu/alu_au/lt1_c44 ,open_n6250}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_44  (
    .a(ds2[44]),
    .b(ds1[44]),
    .c(\exu/alu_au/lt1_c44 ),
    .o({\exu/alu_au/lt1_c45 ,open_n6251}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_45  (
    .a(ds2[45]),
    .b(ds1[45]),
    .c(\exu/alu_au/lt1_c45 ),
    .o({\exu/alu_au/lt1_c46 ,open_n6252}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_46  (
    .a(ds2[46]),
    .b(ds1[46]),
    .c(\exu/alu_au/lt1_c46 ),
    .o({\exu/alu_au/lt1_c47 ,open_n6253}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_47  (
    .a(ds2[47]),
    .b(ds1[47]),
    .c(\exu/alu_au/lt1_c47 ),
    .o({\exu/alu_au/lt1_c48 ,open_n6254}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_48  (
    .a(ds2[48]),
    .b(ds1[48]),
    .c(\exu/alu_au/lt1_c48 ),
    .o({\exu/alu_au/lt1_c49 ,open_n6255}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_49  (
    .a(ds2[49]),
    .b(ds1[49]),
    .c(\exu/alu_au/lt1_c49 ),
    .o({\exu/alu_au/lt1_c50 ,open_n6256}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_5  (
    .a(ds2[5]),
    .b(ds1[5]),
    .c(\exu/alu_au/lt1_c5 ),
    .o({\exu/alu_au/lt1_c6 ,open_n6257}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_50  (
    .a(ds2[50]),
    .b(ds1[50]),
    .c(\exu/alu_au/lt1_c50 ),
    .o({\exu/alu_au/lt1_c51 ,open_n6258}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_51  (
    .a(ds2[51]),
    .b(ds1[51]),
    .c(\exu/alu_au/lt1_c51 ),
    .o({\exu/alu_au/lt1_c52 ,open_n6259}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_52  (
    .a(ds2[52]),
    .b(ds1[52]),
    .c(\exu/alu_au/lt1_c52 ),
    .o({\exu/alu_au/lt1_c53 ,open_n6260}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_53  (
    .a(ds2[53]),
    .b(ds1[53]),
    .c(\exu/alu_au/lt1_c53 ),
    .o({\exu/alu_au/lt1_c54 ,open_n6261}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_54  (
    .a(ds2[54]),
    .b(ds1[54]),
    .c(\exu/alu_au/lt1_c54 ),
    .o({\exu/alu_au/lt1_c55 ,open_n6262}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_55  (
    .a(ds2[55]),
    .b(ds1[55]),
    .c(\exu/alu_au/lt1_c55 ),
    .o({\exu/alu_au/lt1_c56 ,open_n6263}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_56  (
    .a(ds2[56]),
    .b(ds1[56]),
    .c(\exu/alu_au/lt1_c56 ),
    .o({\exu/alu_au/lt1_c57 ,open_n6264}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_57  (
    .a(ds2[57]),
    .b(ds1[57]),
    .c(\exu/alu_au/lt1_c57 ),
    .o({\exu/alu_au/lt1_c58 ,open_n6265}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_58  (
    .a(ds2[58]),
    .b(ds1[58]),
    .c(\exu/alu_au/lt1_c58 ),
    .o({\exu/alu_au/lt1_c59 ,open_n6266}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_59  (
    .a(ds2[59]),
    .b(ds1[59]),
    .c(\exu/alu_au/lt1_c59 ),
    .o({\exu/alu_au/lt1_c60 ,open_n6267}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_6  (
    .a(ds2[6]),
    .b(ds1[6]),
    .c(\exu/alu_au/lt1_c6 ),
    .o({\exu/alu_au/lt1_c7 ,open_n6268}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_60  (
    .a(ds2[60]),
    .b(ds1[60]),
    .c(\exu/alu_au/lt1_c60 ),
    .o({\exu/alu_au/lt1_c61 ,open_n6269}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_61  (
    .a(ds2[61]),
    .b(ds1[61]),
    .c(\exu/alu_au/lt1_c61 ),
    .o({\exu/alu_au/lt1_c62 ,open_n6270}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_62  (
    .a(ds2[62]),
    .b(ds1[62]),
    .c(\exu/alu_au/lt1_c62 ),
    .o({\exu/alu_au/lt1_c63 ,open_n6271}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_63  (
    .a(ds2[63]),
    .b(ds1[63]),
    .c(\exu/alu_au/lt1_c63 ),
    .o({\exu/alu_au/lt1_c64 ,open_n6272}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_7  (
    .a(ds2[7]),
    .b(ds1[7]),
    .c(\exu/alu_au/lt1_c7 ),
    .o({\exu/alu_au/lt1_c8 ,open_n6273}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_8  (
    .a(ds2[8]),
    .b(ds1[8]),
    .c(\exu/alu_au/lt1_c8 ),
    .o({\exu/alu_au/lt1_c9 ,open_n6274}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_9  (
    .a(ds2[9]),
    .b(ds1[9]),
    .c(\exu/alu_au/lt1_c9 ),
    .o({\exu/alu_au/lt1_c10 ,open_n6275}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \exu/alu_au/lt1_cin  (
    .a(1'b0),
    .o({\exu/alu_au/lt1_c0 ,open_n6278}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \exu/alu_au/lt1_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\exu/alu_au/lt1_c64 ),
    .o({open_n6279,\exu/alu_au/n12 }));
  reg_sr_as_w1 \exu/csr_write_reg  (
    .clk(clk_pad),
    .d(ex_csr_write),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_csr_write));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/ebreak_reg  (
    .clk(clk_pad),
    .d(ex_ebreak),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ebreak));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ecall_reg  (
    .clk(clk_pad),
    .d(ex_ecall),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ecall));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/gpr_write_reg  (
    .clk(clk_pad),
    .d(ex_gpr_write),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_gpr_write));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/id_jmp_reg  (
    .clk(clk_pad),
    .d(ex_jmp),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_jmp));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/id_system_reg  (
    .clk(clk_pad),
    .d(ex_system),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_system));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ill_ins_reg  (
    .clk(clk_pad),
    .d(ex_ill_ins),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ill_ins));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ins_acc_fault_reg  (
    .clk(clk_pad),
    .d(ex_ins_acc_fault),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ins_acc_fault));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ins_addr_mis_reg  (
    .clk(clk_pad),
    .d(ex_ins_addr_mis),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ins_addr_mis));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ins_page_fault_reg  (
    .clk(clk_pad),
    .d(ex_ins_page_fault),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ins_page_fault));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/int_acc_reg  (
    .clk(clk_pad),
    .d(ex_int_acc),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_int_acc));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ld_acc_fault_reg  (
    .clk(clk_pad),
    .d(load_acc_fault),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ld_acc_fault));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ld_addr_mis_reg  (
    .clk(clk_pad),
    .d(\exu/load_addr_mis ),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ld_addr_mis));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ld_page_fault_reg  (
    .clk(clk_pad),
    .d(load_page_fault),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ld_page_fault));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/m_ret_reg  (
    .clk(clk_pad),
    .d(ex_m_ret),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_m_ret));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/pc_jmp_reg  (
    .clk(clk_pad),
    .d(jmp),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(pc_jmp));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg0_b0  (
    .clk(clk_pad),
    .d(\exu/n52 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/shift_count [0]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b1  (
    .clk(clk_pad),
    .d(\exu/n52 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/shift_count [1]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b2  (
    .clk(clk_pad),
    .d(\exu/n52 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/shift_count [2]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b3  (
    .clk(clk_pad),
    .d(\exu/n52 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/shift_count [3]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b4  (
    .clk(clk_pad),
    .d(\exu/n52 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/shift_count [4]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b5  (
    .clk(clk_pad),
    .d(\exu/n52 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/shift_count [5]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b6  (
    .clk(clk_pad),
    .d(\exu/n52 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/shift_count [6]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b7  (
    .clk(clk_pad),
    .d(\exu/n52 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/shift_count [7]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg1_b0  (
    .clk(clk_pad),
    .d(\exu/n64 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[0]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b1  (
    .clk(clk_pad),
    .d(\exu/n64 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[1]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b10  (
    .clk(clk_pad),
    .d(\exu/n64 [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[10]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b11  (
    .clk(clk_pad),
    .d(\exu/n64 [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[11]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b12  (
    .clk(clk_pad),
    .d(\exu/n64 [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[12]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b13  (
    .clk(clk_pad),
    .d(\exu/n64 [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[13]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b14  (
    .clk(clk_pad),
    .d(\exu/n64 [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[14]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b15  (
    .clk(clk_pad),
    .d(\exu/n64 [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[15]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b16  (
    .clk(clk_pad),
    .d(\exu/n64 [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[16]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b17  (
    .clk(clk_pad),
    .d(\exu/n64 [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[17]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b18  (
    .clk(clk_pad),
    .d(\exu/n64 [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[18]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b19  (
    .clk(clk_pad),
    .d(\exu/n64 [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[19]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b2  (
    .clk(clk_pad),
    .d(\exu/n64 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[2]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b20  (
    .clk(clk_pad),
    .d(\exu/n64 [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[20]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b21  (
    .clk(clk_pad),
    .d(\exu/n64 [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[21]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b22  (
    .clk(clk_pad),
    .d(\exu/n64 [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[22]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b23  (
    .clk(clk_pad),
    .d(\exu/n64 [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[23]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b24  (
    .clk(clk_pad),
    .d(\exu/n64 [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[24]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b25  (
    .clk(clk_pad),
    .d(\exu/n64 [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[25]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b26  (
    .clk(clk_pad),
    .d(\exu/n64 [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[26]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b27  (
    .clk(clk_pad),
    .d(\exu/n64 [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[27]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b28  (
    .clk(clk_pad),
    .d(\exu/n64 [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[28]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b29  (
    .clk(clk_pad),
    .d(\exu/n64 [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[29]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b3  (
    .clk(clk_pad),
    .d(\exu/n64 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[3]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b30  (
    .clk(clk_pad),
    .d(\exu/n64 [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[30]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b31  (
    .clk(clk_pad),
    .d(\exu/n64 [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[31]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b32  (
    .clk(clk_pad),
    .d(\exu/n64 [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[32]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b33  (
    .clk(clk_pad),
    .d(\exu/n64 [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[33]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b34  (
    .clk(clk_pad),
    .d(\exu/n64 [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[34]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b35  (
    .clk(clk_pad),
    .d(\exu/n64 [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[35]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b36  (
    .clk(clk_pad),
    .d(\exu/n64 [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[36]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b37  (
    .clk(clk_pad),
    .d(\exu/n64 [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[37]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b38  (
    .clk(clk_pad),
    .d(\exu/n64 [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[38]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b39  (
    .clk(clk_pad),
    .d(\exu/n64 [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[39]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b4  (
    .clk(clk_pad),
    .d(\exu/n64 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[4]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b40  (
    .clk(clk_pad),
    .d(\exu/n64 [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[40]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b41  (
    .clk(clk_pad),
    .d(\exu/n64 [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[41]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b42  (
    .clk(clk_pad),
    .d(\exu/n64 [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[42]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b43  (
    .clk(clk_pad),
    .d(\exu/n64 [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[43]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b44  (
    .clk(clk_pad),
    .d(\exu/n64 [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[44]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b45  (
    .clk(clk_pad),
    .d(\exu/n64 [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[45]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b46  (
    .clk(clk_pad),
    .d(\exu/n64 [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[46]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b47  (
    .clk(clk_pad),
    .d(\exu/n64 [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[47]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b48  (
    .clk(clk_pad),
    .d(\exu/n64 [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[48]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b49  (
    .clk(clk_pad),
    .d(\exu/n64 [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[49]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b5  (
    .clk(clk_pad),
    .d(\exu/n64 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[5]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b50  (
    .clk(clk_pad),
    .d(\exu/n64 [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[50]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b51  (
    .clk(clk_pad),
    .d(\exu/n64 [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[51]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b52  (
    .clk(clk_pad),
    .d(\exu/n64 [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[52]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b53  (
    .clk(clk_pad),
    .d(\exu/n64 [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[53]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b54  (
    .clk(clk_pad),
    .d(\exu/n64 [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[54]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b55  (
    .clk(clk_pad),
    .d(\exu/n64 [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[55]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b56  (
    .clk(clk_pad),
    .d(\exu/n64 [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[56]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b57  (
    .clk(clk_pad),
    .d(\exu/n64 [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[57]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b58  (
    .clk(clk_pad),
    .d(\exu/n64 [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[58]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b59  (
    .clk(clk_pad),
    .d(\exu/n64 [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[59]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b6  (
    .clk(clk_pad),
    .d(\exu/n64 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[6]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b60  (
    .clk(clk_pad),
    .d(\exu/n64 [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[60]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b61  (
    .clk(clk_pad),
    .d(\exu/n64 [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[61]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b62  (
    .clk(clk_pad),
    .d(\exu/n64 [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[62]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b63  (
    .clk(clk_pad),
    .d(\exu/n64 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[63]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b7  (
    .clk(clk_pad),
    .d(\exu/n64 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[7]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b8  (
    .clk(clk_pad),
    .d(\exu/n64 [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[8]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b9  (
    .clk(clk_pad),
    .d(\exu/n64 [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_rd[9]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg2_b0  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[0]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b1  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[1]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b10  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[10]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b11  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[11]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b12  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[12]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b13  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[13]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b14  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[14]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b15  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[15]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b16  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[16]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b17  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[17]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b18  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[18]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b19  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[19]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b2  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[2]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b20  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[20]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b21  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[21]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b22  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[22]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b23  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[23]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b24  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[24]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b25  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[25]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b26  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[26]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b27  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[27]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b28  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[28]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b29  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[29]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b3  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[3]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b30  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[30]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b31  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[31]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b32  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[32]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b33  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[33]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b34  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[34]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b35  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[35]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b36  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[36]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b37  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[37]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b38  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[38]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b39  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[39]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b4  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[4]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b40  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[40]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b41  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[41]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b42  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[42]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b43  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[43]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b44  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[44]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b45  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[45]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b46  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[46]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b47  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[47]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b48  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[48]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b49  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[49]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b5  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[5]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b50  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[50]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b51  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[51]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b52  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[52]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b53  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[53]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b54  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[54]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b55  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[55]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b56  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[56]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b57  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[57]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b58  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[58]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b59  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[59]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b6  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[6]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b60  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[60]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b61  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[61]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b62  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[62]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b63  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[63]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b7  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[7]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b8  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[8]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b9  (
    .clk(clk_pad),
    .d(\exu/alu_data_mem_csr [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(data_csr[9]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b0  (
    .clk(clk_pad),
    .d(addr_ex[0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[0]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b1  (
    .clk(clk_pad),
    .d(addr_ex[1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[1]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b10  (
    .clk(clk_pad),
    .d(addr_ex[10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[10]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b11  (
    .clk(clk_pad),
    .d(addr_ex[11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[11]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b12  (
    .clk(clk_pad),
    .d(addr_ex[12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[12]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b13  (
    .clk(clk_pad),
    .d(addr_ex[13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[13]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b14  (
    .clk(clk_pad),
    .d(addr_ex[14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[14]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b15  (
    .clk(clk_pad),
    .d(addr_ex[15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[15]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b16  (
    .clk(clk_pad),
    .d(addr_ex[16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[16]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b17  (
    .clk(clk_pad),
    .d(addr_ex[17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[17]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b18  (
    .clk(clk_pad),
    .d(addr_ex[18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[18]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b19  (
    .clk(clk_pad),
    .d(addr_ex[19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[19]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b2  (
    .clk(clk_pad),
    .d(addr_ex[2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[2]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b20  (
    .clk(clk_pad),
    .d(addr_ex[20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[20]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b21  (
    .clk(clk_pad),
    .d(addr_ex[21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[21]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b22  (
    .clk(clk_pad),
    .d(addr_ex[22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[22]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b23  (
    .clk(clk_pad),
    .d(addr_ex[23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[23]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b24  (
    .clk(clk_pad),
    .d(addr_ex[24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[24]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b25  (
    .clk(clk_pad),
    .d(addr_ex[25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[25]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b26  (
    .clk(clk_pad),
    .d(addr_ex[26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[26]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b27  (
    .clk(clk_pad),
    .d(addr_ex[27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[27]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b28  (
    .clk(clk_pad),
    .d(addr_ex[28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[28]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b29  (
    .clk(clk_pad),
    .d(addr_ex[29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[29]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b3  (
    .clk(clk_pad),
    .d(addr_ex[3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[3]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b30  (
    .clk(clk_pad),
    .d(addr_ex[30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[30]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b31  (
    .clk(clk_pad),
    .d(addr_ex[31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[31]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b32  (
    .clk(clk_pad),
    .d(addr_ex[32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[32]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b33  (
    .clk(clk_pad),
    .d(addr_ex[33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[33]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b34  (
    .clk(clk_pad),
    .d(addr_ex[34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[34]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b35  (
    .clk(clk_pad),
    .d(addr_ex[35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[35]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b36  (
    .clk(clk_pad),
    .d(addr_ex[36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[36]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b37  (
    .clk(clk_pad),
    .d(addr_ex[37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[37]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b38  (
    .clk(clk_pad),
    .d(addr_ex[38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[38]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b39  (
    .clk(clk_pad),
    .d(addr_ex[39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[39]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b4  (
    .clk(clk_pad),
    .d(addr_ex[4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[4]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b40  (
    .clk(clk_pad),
    .d(addr_ex[40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[40]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b41  (
    .clk(clk_pad),
    .d(addr_ex[41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[41]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b42  (
    .clk(clk_pad),
    .d(addr_ex[42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[42]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b43  (
    .clk(clk_pad),
    .d(addr_ex[43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[43]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b44  (
    .clk(clk_pad),
    .d(addr_ex[44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[44]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b45  (
    .clk(clk_pad),
    .d(addr_ex[45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[45]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b46  (
    .clk(clk_pad),
    .d(addr_ex[46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[46]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b47  (
    .clk(clk_pad),
    .d(addr_ex[47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[47]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b48  (
    .clk(clk_pad),
    .d(addr_ex[48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[48]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b49  (
    .clk(clk_pad),
    .d(addr_ex[49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[49]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b5  (
    .clk(clk_pad),
    .d(addr_ex[5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[5]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b50  (
    .clk(clk_pad),
    .d(addr_ex[50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[50]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b51  (
    .clk(clk_pad),
    .d(addr_ex[51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[51]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b52  (
    .clk(clk_pad),
    .d(addr_ex[52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[52]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b53  (
    .clk(clk_pad),
    .d(addr_ex[53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[53]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b54  (
    .clk(clk_pad),
    .d(addr_ex[54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[54]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b55  (
    .clk(clk_pad),
    .d(addr_ex[55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[55]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b56  (
    .clk(clk_pad),
    .d(addr_ex[56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[56]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b57  (
    .clk(clk_pad),
    .d(addr_ex[57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[57]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b58  (
    .clk(clk_pad),
    .d(addr_ex[58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[58]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b59  (
    .clk(clk_pad),
    .d(addr_ex[59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[59]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b6  (
    .clk(clk_pad),
    .d(addr_ex[6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[6]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b60  (
    .clk(clk_pad),
    .d(addr_ex[60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[60]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b61  (
    .clk(clk_pad),
    .d(addr_ex[61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[61]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b62  (
    .clk(clk_pad),
    .d(addr_ex[62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[62]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b63  (
    .clk(clk_pad),
    .d(addr_ex[63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[63]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b7  (
    .clk(clk_pad),
    .d(addr_ex[7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[7]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b8  (
    .clk(clk_pad),
    .d(addr_ex[8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[8]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b9  (
    .clk(clk_pad),
    .d(addr_ex[9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(new_pc[9]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg4_b0  (
    .clk(clk_pad),
    .d(ex_ins_pc[0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[0]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b1  (
    .clk(clk_pad),
    .d(ex_ins_pc[1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[1]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b10  (
    .clk(clk_pad),
    .d(ex_ins_pc[10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[10]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b11  (
    .clk(clk_pad),
    .d(ex_ins_pc[11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[11]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b12  (
    .clk(clk_pad),
    .d(ex_ins_pc[12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[12]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b13  (
    .clk(clk_pad),
    .d(ex_ins_pc[13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[13]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b14  (
    .clk(clk_pad),
    .d(ex_ins_pc[14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[14]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b15  (
    .clk(clk_pad),
    .d(ex_ins_pc[15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[15]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b16  (
    .clk(clk_pad),
    .d(ex_ins_pc[16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[16]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b17  (
    .clk(clk_pad),
    .d(ex_ins_pc[17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[17]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b18  (
    .clk(clk_pad),
    .d(ex_ins_pc[18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[18]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b19  (
    .clk(clk_pad),
    .d(ex_ins_pc[19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[19]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b2  (
    .clk(clk_pad),
    .d(ex_ins_pc[2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[2]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b20  (
    .clk(clk_pad),
    .d(ex_ins_pc[20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[20]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b21  (
    .clk(clk_pad),
    .d(ex_ins_pc[21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[21]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b22  (
    .clk(clk_pad),
    .d(ex_ins_pc[22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[22]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b23  (
    .clk(clk_pad),
    .d(ex_ins_pc[23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[23]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b24  (
    .clk(clk_pad),
    .d(ex_ins_pc[24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[24]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b25  (
    .clk(clk_pad),
    .d(ex_ins_pc[25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[25]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b26  (
    .clk(clk_pad),
    .d(ex_ins_pc[26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[26]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b27  (
    .clk(clk_pad),
    .d(ex_ins_pc[27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[27]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b28  (
    .clk(clk_pad),
    .d(ex_ins_pc[28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[28]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b29  (
    .clk(clk_pad),
    .d(ex_ins_pc[29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[29]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b3  (
    .clk(clk_pad),
    .d(ex_ins_pc[3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[3]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b30  (
    .clk(clk_pad),
    .d(ex_ins_pc[30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[30]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b31  (
    .clk(clk_pad),
    .d(ex_ins_pc[31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[31]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b32  (
    .clk(clk_pad),
    .d(ex_ins_pc[32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[32]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b33  (
    .clk(clk_pad),
    .d(ex_ins_pc[33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[33]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b34  (
    .clk(clk_pad),
    .d(ex_ins_pc[34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[34]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b35  (
    .clk(clk_pad),
    .d(ex_ins_pc[35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[35]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b36  (
    .clk(clk_pad),
    .d(ex_ins_pc[36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[36]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b37  (
    .clk(clk_pad),
    .d(ex_ins_pc[37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[37]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b38  (
    .clk(clk_pad),
    .d(ex_ins_pc[38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[38]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b39  (
    .clk(clk_pad),
    .d(ex_ins_pc[39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[39]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b4  (
    .clk(clk_pad),
    .d(ex_ins_pc[4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[4]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b40  (
    .clk(clk_pad),
    .d(ex_ins_pc[40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[40]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b41  (
    .clk(clk_pad),
    .d(ex_ins_pc[41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[41]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b42  (
    .clk(clk_pad),
    .d(ex_ins_pc[42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[42]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b43  (
    .clk(clk_pad),
    .d(ex_ins_pc[43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[43]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b44  (
    .clk(clk_pad),
    .d(ex_ins_pc[44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[44]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b45  (
    .clk(clk_pad),
    .d(ex_ins_pc[45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[45]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b46  (
    .clk(clk_pad),
    .d(ex_ins_pc[46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[46]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b47  (
    .clk(clk_pad),
    .d(ex_ins_pc[47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[47]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b48  (
    .clk(clk_pad),
    .d(ex_ins_pc[48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[48]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b49  (
    .clk(clk_pad),
    .d(ex_ins_pc[49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[49]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b5  (
    .clk(clk_pad),
    .d(ex_ins_pc[5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[5]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b50  (
    .clk(clk_pad),
    .d(ex_ins_pc[50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[50]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b51  (
    .clk(clk_pad),
    .d(ex_ins_pc[51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[51]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b52  (
    .clk(clk_pad),
    .d(ex_ins_pc[52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[52]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b53  (
    .clk(clk_pad),
    .d(ex_ins_pc[53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[53]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b54  (
    .clk(clk_pad),
    .d(ex_ins_pc[54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[54]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b55  (
    .clk(clk_pad),
    .d(ex_ins_pc[55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[55]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b56  (
    .clk(clk_pad),
    .d(ex_ins_pc[56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[56]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b57  (
    .clk(clk_pad),
    .d(ex_ins_pc[57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[57]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b58  (
    .clk(clk_pad),
    .d(ex_ins_pc[58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[58]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b59  (
    .clk(clk_pad),
    .d(ex_ins_pc[59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[59]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b6  (
    .clk(clk_pad),
    .d(ex_ins_pc[6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[6]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b60  (
    .clk(clk_pad),
    .d(ex_ins_pc[60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[60]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b61  (
    .clk(clk_pad),
    .d(ex_ins_pc[61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[61]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b62  (
    .clk(clk_pad),
    .d(ex_ins_pc[62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[62]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b63  (
    .clk(clk_pad),
    .d(ex_ins_pc[63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[63]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b7  (
    .clk(clk_pad),
    .d(ex_ins_pc[7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[7]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b8  (
    .clk(clk_pad),
    .d(ex_ins_pc[8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[8]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b9  (
    .clk(clk_pad),
    .d(ex_ins_pc[9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_ins_pc[9]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b0  (
    .clk(clk_pad),
    .d(\exu/n71 [0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[0]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b1  (
    .clk(clk_pad),
    .d(\exu/n71 [1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[1]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b10  (
    .clk(clk_pad),
    .d(\exu/n71 [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[10]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b11  (
    .clk(clk_pad),
    .d(\exu/n71 [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[11]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b12  (
    .clk(clk_pad),
    .d(\exu/n71 [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[12]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b13  (
    .clk(clk_pad),
    .d(\exu/n71 [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[13]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b14  (
    .clk(clk_pad),
    .d(\exu/n71 [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[14]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b15  (
    .clk(clk_pad),
    .d(\exu/n71 [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[15]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b16  (
    .clk(clk_pad),
    .d(\exu/n71 [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[16]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b17  (
    .clk(clk_pad),
    .d(\exu/n71 [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[17]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b18  (
    .clk(clk_pad),
    .d(\exu/n71 [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[18]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b19  (
    .clk(clk_pad),
    .d(\exu/n71 [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[19]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b2  (
    .clk(clk_pad),
    .d(\exu/n71 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[2]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b20  (
    .clk(clk_pad),
    .d(\exu/n71 [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[20]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b21  (
    .clk(clk_pad),
    .d(\exu/n71 [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[21]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b22  (
    .clk(clk_pad),
    .d(\exu/n71 [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[22]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b23  (
    .clk(clk_pad),
    .d(\exu/n71 [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[23]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b24  (
    .clk(clk_pad),
    .d(\exu/n71 [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[24]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b25  (
    .clk(clk_pad),
    .d(\exu/n71 [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[25]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b26  (
    .clk(clk_pad),
    .d(\exu/n71 [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[26]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b27  (
    .clk(clk_pad),
    .d(\exu/n71 [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[27]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b28  (
    .clk(clk_pad),
    .d(\exu/n71 [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[28]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b29  (
    .clk(clk_pad),
    .d(\exu/n71 [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[29]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b3  (
    .clk(clk_pad),
    .d(\exu/n71 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[3]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b30  (
    .clk(clk_pad),
    .d(\exu/n71 [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[30]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b31  (
    .clk(clk_pad),
    .d(\exu/n71 [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[31]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b32  (
    .clk(clk_pad),
    .d(\exu/n71 [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[32]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b33  (
    .clk(clk_pad),
    .d(\exu/n71 [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[33]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b34  (
    .clk(clk_pad),
    .d(\exu/n71 [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[34]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b35  (
    .clk(clk_pad),
    .d(\exu/n71 [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[35]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b36  (
    .clk(clk_pad),
    .d(\exu/n71 [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[36]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b37  (
    .clk(clk_pad),
    .d(\exu/n71 [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[37]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b38  (
    .clk(clk_pad),
    .d(\exu/n71 [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[38]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b39  (
    .clk(clk_pad),
    .d(\exu/n71 [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[39]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b4  (
    .clk(clk_pad),
    .d(\exu/n71 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[4]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b40  (
    .clk(clk_pad),
    .d(\exu/n71 [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[40]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b41  (
    .clk(clk_pad),
    .d(\exu/n71 [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[41]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b42  (
    .clk(clk_pad),
    .d(\exu/n71 [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[42]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b43  (
    .clk(clk_pad),
    .d(\exu/n71 [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[43]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b44  (
    .clk(clk_pad),
    .d(\exu/n71 [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[44]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b45  (
    .clk(clk_pad),
    .d(\exu/n71 [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[45]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b46  (
    .clk(clk_pad),
    .d(\exu/n71 [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[46]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b47  (
    .clk(clk_pad),
    .d(\exu/n71 [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[47]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b48  (
    .clk(clk_pad),
    .d(\exu/n71 [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[48]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b49  (
    .clk(clk_pad),
    .d(\exu/n71 [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[49]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b5  (
    .clk(clk_pad),
    .d(\exu/n71 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[5]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b50  (
    .clk(clk_pad),
    .d(\exu/n71 [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[50]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b51  (
    .clk(clk_pad),
    .d(\exu/n71 [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[51]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b52  (
    .clk(clk_pad),
    .d(\exu/n71 [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[52]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b53  (
    .clk(clk_pad),
    .d(\exu/n71 [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[53]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b54  (
    .clk(clk_pad),
    .d(\exu/n71 [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[54]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b55  (
    .clk(clk_pad),
    .d(\exu/n71 [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[55]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b56  (
    .clk(clk_pad),
    .d(\exu/n71 [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[56]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b57  (
    .clk(clk_pad),
    .d(\exu/n71 [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[57]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b58  (
    .clk(clk_pad),
    .d(\exu/n71 [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[58]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b59  (
    .clk(clk_pad),
    .d(\exu/n71 [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[59]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b6  (
    .clk(clk_pad),
    .d(\exu/n71 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[6]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b60  (
    .clk(clk_pad),
    .d(\exu/n71 [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[60]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b61  (
    .clk(clk_pad),
    .d(\exu/n71 [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[61]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b62  (
    .clk(clk_pad),
    .d(\exu/n71 [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[62]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b63  (
    .clk(clk_pad),
    .d(\exu/n71 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[63]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b7  (
    .clk(clk_pad),
    .d(\exu/n71 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[7]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b8  (
    .clk(clk_pad),
    .d(\exu/n71 [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[8]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b9  (
    .clk(clk_pad),
    .d(\exu/n71 [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_exc_code[9]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg6_b0  (
    .clk(clk_pad),
    .d(ex_csr_index[0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[0]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b1  (
    .clk(clk_pad),
    .d(ex_csr_index[1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[1]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b10  (
    .clk(clk_pad),
    .d(ex_csr_index[10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[10]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b11  (
    .clk(clk_pad),
    .d(ex_csr_index[11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[11]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b2  (
    .clk(clk_pad),
    .d(ex_csr_index[2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[2]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b3  (
    .clk(clk_pad),
    .d(ex_csr_index[3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[3]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b4  (
    .clk(clk_pad),
    .d(ex_csr_index[4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[4]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b5  (
    .clk(clk_pad),
    .d(ex_csr_index[5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[5]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b6  (
    .clk(clk_pad),
    .d(ex_csr_index[6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[6]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b7  (
    .clk(clk_pad),
    .d(ex_csr_index[7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[7]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b8  (
    .clk(clk_pad),
    .d(ex_csr_index[8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[8]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b9  (
    .clk(clk_pad),
    .d(ex_csr_index[9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(csr_index[9]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg7_b0  (
    .clk(clk_pad),
    .d(ex_rd_index[0]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_rd_index[0]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg7_b1  (
    .clk(clk_pad),
    .d(ex_rd_index[1]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_rd_index[1]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg7_b2  (
    .clk(clk_pad),
    .d(ex_rd_index[2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_rd_index[2]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg7_b3  (
    .clk(clk_pad),
    .d(ex_rd_index[3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_rd_index[3]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg7_b4  (
    .clk(clk_pad),
    .d(ex_rd_index[4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(wb_rd_index[4]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg8_b0  (
    .clk(clk_pad),
    .d(\exu/n45 [0]),
    .en(~ex_nop),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/main_state [0]));  // ../../RTL/CPU/EX/exu.v(268)
  reg_sr_as_w1 \exu/reg8_b1  (
    .clk(clk_pad),
    .d(\exu/n45 [1]),
    .en(~ex_nop),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/main_state [1]));  // ../../RTL/CPU/EX/exu.v(268)
  reg_sr_as_w1 \exu/reg8_b2  (
    .clk(clk_pad),
    .d(\exu/n45 [2]),
    .en(~ex_nop),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/main_state [2]));  // ../../RTL/CPU/EX/exu.v(268)
  reg_sr_as_w1 \exu/reg8_b3  (
    .clk(clk_pad),
    .d(\exu/n45 [3]),
    .en(~ex_nop),
    .reset(rst_pad),
    .set(1'b0),
    .q(\exu/main_state [3]));  // ../../RTL/CPU/EX/exu.v(268)
  reg_sr_as_w1 \exu/s_ret_reg  (
    .clk(clk_pad),
    .d(ex_s_ret),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_s_ret));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/st_acc_fault_reg  (
    .clk(clk_pad),
    .d(\exu/n90 ),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_st_acc_fault));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/st_addr_mis_reg  (
    .clk(clk_pad),
    .d(\exu/n88 ),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_st_addr_mis));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/st_page_fault_reg  (
    .clk(clk_pad),
    .d(\exu/n92 ),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_st_page_fault));  // ../../RTL/CPU/EX/exu.v(448)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \exu/sub0/u0  (
    .a(\exu/shift_count [0]),
    .b(1'b1),
    .c(\exu/sub0/c0 ),
    .o({\exu/sub0/c1 ,\exu/n50 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \exu/sub0/u1  (
    .a(\exu/shift_count [1]),
    .b(1'b0),
    .c(\exu/sub0/c1 ),
    .o({\exu/sub0/c2 ,\exu/n50 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \exu/sub0/u2  (
    .a(\exu/shift_count [2]),
    .b(1'b0),
    .c(\exu/sub0/c2 ),
    .o({\exu/sub0/c3 ,\exu/n50 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \exu/sub0/u3  (
    .a(\exu/shift_count [3]),
    .b(1'b0),
    .c(\exu/sub0/c3 ),
    .o({\exu/sub0/c4 ,\exu/n50 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \exu/sub0/u4  (
    .a(\exu/shift_count [4]),
    .b(1'b0),
    .c(\exu/sub0/c4 ),
    .o({\exu/sub0/c5 ,\exu/n50 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \exu/sub0/u5  (
    .a(\exu/shift_count [5]),
    .b(1'b0),
    .c(\exu/sub0/c5 ),
    .o({\exu/sub0/c6 ,\exu/n50 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \exu/sub0/u6  (
    .a(\exu/shift_count [6]),
    .b(1'b0),
    .c(\exu/sub0/c6 ),
    .o({\exu/sub0/c7 ,\exu/n50 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \exu/sub0/u7  (
    .a(\exu/shift_count [7]),
    .b(1'b0),
    .c(\exu/sub0/c7 ),
    .o({open_n6280,\exu/n50 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \exu/sub0/ucin  (
    .a(1'b0),
    .o({\exu/sub0/c0 ,open_n6283}));
  reg_sr_as_w1 \exu/valid_reg  (
    .clk(clk_pad),
    .d(\exu/n95 ),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_valid));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \ins_dec/amo_reg  (
    .clk(clk_pad),
    .d(\ins_dec/op_amo ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(amo));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/and_clr_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n71 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(and_clr));  // ../../RTL/CPU/ID/ins_dec.v(674)
  reg_sr_as_w1 \ins_dec/cache_flush_reg  (
    .clk(clk_pad),
    .d(\ins_dec/ins_fence ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(cache_flush));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/cache_reset_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n225 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(cache_reset));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/csr_write_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n239 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_write));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/ebreak_reg  (
    .clk(clk_pad),
    .d(\ins_dec/ins_ebreak ),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ebreak));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/ecall_reg  (
    .clk(clk_pad),
    .d(\ins_dec/ins_ecall ),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ecall));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/gpr_write_reg  (
    .clk(clk_pad),
    .d(\ins_dec/dec_gpr_write ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_gpr_write));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/id_jmp_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n302 ),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_jmp));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/id_system_reg  (
    .clk(clk_pad),
    .d(id_system),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_system));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/ill_ins_reg  (
    .clk(clk_pad),
    .d(id_ill_ins),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ill_ins));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/ins_acc_fault_reg  (
    .clk(clk_pad),
    .d(id_ins_acc_fault),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_acc_fault));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/ins_addr_mis_reg  (
    .clk(clk_pad),
    .d(id_ins_addr_mis),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_addr_mis));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/ins_page_fault_reg  (
    .clk(clk_pad),
    .d(id_ins_page_fault),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_page_fault));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/int_acc_reg  (
    .clk(clk_pad),
    .d(id_int_acc),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_int_acc));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/jmp_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n59 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(jmp));  // ../../RTL/CPU/ID/ins_dec.v(674)
  reg_sr_as_w1 \ins_dec/load_reg  (
    .clk(clk_pad),
    .d(\ins_dec/op_load ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(load));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/m_ret_reg  (
    .clk(clk_pad),
    .d(1'b0),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_m_ret));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/mem_csr_data_add_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n146 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_add));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_and_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n148 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_and));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_ds2_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n145 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_ds2));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_max_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n155 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_max));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_min_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n158 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_min));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_or_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n151 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_or));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_xor_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n152 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_xor));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_add_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n132 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_add));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_and_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n134 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_and));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_ds1_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n126 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_ds1));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_or_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n135 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_or));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_slt_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n139 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_slt));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_sub_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n133 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_sub));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_xor_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n136 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_xor));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/reg0_b0  (
    .clk(clk_pad),
    .d(\ins_dec/sbyte ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_size[0]));  // ../../RTL/CPU/ID/ins_dec.v(689)
  reg_sr_as_w1 \ins_dec/reg0_b1  (
    .clk(clk_pad),
    .d(\ins_dec/dbyte ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_size[1]));  // ../../RTL/CPU/ID/ins_dec.v(689)
  reg_ar_ss_w1 \ins_dec/reg0_b2  (
    .clk(clk_pad),
    .d(\ins_dec/qbyte ),
    .en(~id_hold),
    .reset(1'b0),
    .set(\ins_dec/n107 ),
    .q(ex_size[2]));  // ../../RTL/CPU/ID/ins_dec.v(689)
  reg_sr_as_w1 \ins_dec/reg0_b3  (
    .clk(clk_pad),
    .d(\ins_dec/obyte ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_size[3]));  // ../../RTL/CPU/ID/ins_dec.v(689)
  reg_sr_as_w1 \ins_dec/reg10_b0  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[0]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b1  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[1]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b10  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[10]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b11  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[11]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b12  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[12]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b13  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[13]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b14  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[14]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b15  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[15]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b16  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[16]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b17  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[17]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b18  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[18]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b19  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[19]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b2  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[2]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b20  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[20]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b21  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[21]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b22  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[22]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b23  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[23]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b24  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[24]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b25  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[25]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b26  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[26]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b27  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[27]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b28  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[28]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b29  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[29]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b3  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[3]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b30  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[30]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b31  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[31]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b4  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[4]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b5  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[5]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b6  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[6]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b7  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[7]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b8  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[8]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b9  (
    .clk(clk_pad),
    .d(\ins_dec/n342 [9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[9]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b0  (
    .clk(clk_pad),
    .d(id_ins_pc[0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[0]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b1  (
    .clk(clk_pad),
    .d(id_ins_pc[1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[1]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b10  (
    .clk(clk_pad),
    .d(id_ins_pc[10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[10]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b11  (
    .clk(clk_pad),
    .d(id_ins_pc[11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[11]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b12  (
    .clk(clk_pad),
    .d(id_ins_pc[12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[12]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b13  (
    .clk(clk_pad),
    .d(id_ins_pc[13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[13]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b14  (
    .clk(clk_pad),
    .d(id_ins_pc[14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[14]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b15  (
    .clk(clk_pad),
    .d(id_ins_pc[15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[15]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b16  (
    .clk(clk_pad),
    .d(id_ins_pc[16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[16]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b17  (
    .clk(clk_pad),
    .d(id_ins_pc[17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[17]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b18  (
    .clk(clk_pad),
    .d(id_ins_pc[18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[18]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b19  (
    .clk(clk_pad),
    .d(id_ins_pc[19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[19]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b2  (
    .clk(clk_pad),
    .d(id_ins_pc[2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[2]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b20  (
    .clk(clk_pad),
    .d(id_ins_pc[20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[20]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b21  (
    .clk(clk_pad),
    .d(id_ins_pc[21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[21]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b22  (
    .clk(clk_pad),
    .d(id_ins_pc[22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[22]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b23  (
    .clk(clk_pad),
    .d(id_ins_pc[23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[23]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b24  (
    .clk(clk_pad),
    .d(id_ins_pc[24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[24]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b25  (
    .clk(clk_pad),
    .d(id_ins_pc[25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[25]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b26  (
    .clk(clk_pad),
    .d(id_ins_pc[26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[26]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b27  (
    .clk(clk_pad),
    .d(id_ins_pc[27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[27]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b28  (
    .clk(clk_pad),
    .d(id_ins_pc[28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[28]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b29  (
    .clk(clk_pad),
    .d(id_ins_pc[29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[29]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b3  (
    .clk(clk_pad),
    .d(id_ins_pc[3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[3]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b30  (
    .clk(clk_pad),
    .d(id_ins_pc[30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[30]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b31  (
    .clk(clk_pad),
    .d(id_ins_pc[31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[31]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b32  (
    .clk(clk_pad),
    .d(id_ins_pc[32]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[32]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b33  (
    .clk(clk_pad),
    .d(id_ins_pc[33]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[33]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b34  (
    .clk(clk_pad),
    .d(id_ins_pc[34]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[34]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b35  (
    .clk(clk_pad),
    .d(id_ins_pc[35]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[35]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b36  (
    .clk(clk_pad),
    .d(id_ins_pc[36]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[36]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b37  (
    .clk(clk_pad),
    .d(id_ins_pc[37]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[37]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b38  (
    .clk(clk_pad),
    .d(id_ins_pc[38]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[38]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b39  (
    .clk(clk_pad),
    .d(id_ins_pc[39]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[39]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b4  (
    .clk(clk_pad),
    .d(id_ins_pc[4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[4]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b40  (
    .clk(clk_pad),
    .d(id_ins_pc[40]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[40]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b41  (
    .clk(clk_pad),
    .d(id_ins_pc[41]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[41]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b42  (
    .clk(clk_pad),
    .d(id_ins_pc[42]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[42]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b43  (
    .clk(clk_pad),
    .d(id_ins_pc[43]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[43]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b44  (
    .clk(clk_pad),
    .d(id_ins_pc[44]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[44]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b45  (
    .clk(clk_pad),
    .d(id_ins_pc[45]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[45]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b46  (
    .clk(clk_pad),
    .d(id_ins_pc[46]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[46]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b47  (
    .clk(clk_pad),
    .d(id_ins_pc[47]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[47]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b48  (
    .clk(clk_pad),
    .d(id_ins_pc[48]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[48]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b49  (
    .clk(clk_pad),
    .d(id_ins_pc[49]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[49]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b5  (
    .clk(clk_pad),
    .d(id_ins_pc[5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[5]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b50  (
    .clk(clk_pad),
    .d(id_ins_pc[50]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[50]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b51  (
    .clk(clk_pad),
    .d(id_ins_pc[51]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[51]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b52  (
    .clk(clk_pad),
    .d(id_ins_pc[52]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[52]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b53  (
    .clk(clk_pad),
    .d(id_ins_pc[53]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[53]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b54  (
    .clk(clk_pad),
    .d(id_ins_pc[54]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[54]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b55  (
    .clk(clk_pad),
    .d(id_ins_pc[55]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[55]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b56  (
    .clk(clk_pad),
    .d(id_ins_pc[56]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[56]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b57  (
    .clk(clk_pad),
    .d(id_ins_pc[57]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[57]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b58  (
    .clk(clk_pad),
    .d(id_ins_pc[58]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[58]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b59  (
    .clk(clk_pad),
    .d(id_ins_pc[59]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[59]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b6  (
    .clk(clk_pad),
    .d(id_ins_pc[6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[6]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b60  (
    .clk(clk_pad),
    .d(id_ins_pc[60]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[60]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b61  (
    .clk(clk_pad),
    .d(id_ins_pc[61]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[61]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b62  (
    .clk(clk_pad),
    .d(id_ins_pc[62]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[62]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b63  (
    .clk(clk_pad),
    .d(id_ins_pc[63]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[63]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b7  (
    .clk(clk_pad),
    .d(id_ins_pc[7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[7]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b8  (
    .clk(clk_pad),
    .d(id_ins_pc[8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[8]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b9  (
    .clk(clk_pad),
    .d(id_ins_pc[9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[9]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg1_b0  (
    .clk(clk_pad),
    .d(id_ins[20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[0]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b1  (
    .clk(clk_pad),
    .d(id_ins[21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[1]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b10  (
    .clk(clk_pad),
    .d(id_ins[30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[10]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b11  (
    .clk(clk_pad),
    .d(id_ins[31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[11]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b2  (
    .clk(clk_pad),
    .d(id_ins[22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[2]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b3  (
    .clk(clk_pad),
    .d(id_ins[23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[3]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b4  (
    .clk(clk_pad),
    .d(id_ins[24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[4]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b5  (
    .clk(clk_pad),
    .d(id_ins[25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[5]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b6  (
    .clk(clk_pad),
    .d(id_ins[26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[6]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b7  (
    .clk(clk_pad),
    .d(id_ins[27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[7]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b8  (
    .clk(clk_pad),
    .d(id_ins[28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[8]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b9  (
    .clk(clk_pad),
    .d(id_ins[29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[9]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_ar_as_w1 \ins_dec/reg4_b0  (
    .clk(clk_pad),
    .d(id_ins[7]),
    .en(\ins_dec/mux13_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(ex_rd_index[0]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_ar_as_w1 \ins_dec/reg4_b1  (
    .clk(clk_pad),
    .d(id_ins[8]),
    .en(\ins_dec/mux13_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(ex_rd_index[1]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_ar_as_w1 \ins_dec/reg4_b2  (
    .clk(clk_pad),
    .d(id_ins[9]),
    .en(\ins_dec/mux13_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(ex_rd_index[2]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_ar_as_w1 \ins_dec/reg4_b3  (
    .clk(clk_pad),
    .d(id_ins[10]),
    .en(\ins_dec/mux13_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(ex_rd_index[3]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_ar_as_w1 \ins_dec/reg4_b4  (
    .clk(clk_pad),
    .d(id_ins[11]),
    .en(\ins_dec/mux13_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(ex_rd_index[4]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg5_b0  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[0]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b1  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[1]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b10  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[10]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b11  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[11]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b12  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[12]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b13  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[13]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b14  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[14]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b15  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[15]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b16  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[16]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b17  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[17]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b18  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[18]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b19  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[19]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b2  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[2]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b20  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[20]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b21  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[21]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b22  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[22]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b23  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[23]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b24  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[24]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b25  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[25]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b26  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[26]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b27  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[27]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b28  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[28]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b29  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[29]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b3  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[3]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b30  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[30]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b31  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[31]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b32  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [32]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[32]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b33  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [33]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[33]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b34  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [34]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[34]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b35  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [35]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[35]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b36  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [36]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[36]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b37  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [37]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[37]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b38  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [38]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[38]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b39  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [39]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[39]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b4  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[4]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b40  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [40]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[40]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b41  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [41]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[41]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b42  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [42]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[42]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b43  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [43]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[43]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b44  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [44]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[44]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b45  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [45]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[45]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b46  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [46]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[46]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b47  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [47]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[47]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b48  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [48]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[48]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b49  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [49]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[49]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b5  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[5]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b50  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [50]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[50]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b51  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [51]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[51]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b52  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [52]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[52]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b53  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [53]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[53]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b54  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [54]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[54]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b55  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [55]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[55]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b56  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [56]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[56]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b57  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [57]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[57]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b58  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [58]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[58]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b59  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [59]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[59]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b6  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[6]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b60  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [60]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[60]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b61  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [61]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[61]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b62  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [62]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[62]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b63  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [63]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[63]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b7  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[7]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b8  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[8]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b9  (
    .clk(clk_pad),
    .d(\ins_dec/n272 [9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[9]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b0  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[0]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b1  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[1]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b10  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[10]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b11  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[11]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b12  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[12]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b13  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[13]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b14  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[14]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b15  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[15]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b16  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[16]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b17  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[17]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b18  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[18]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b19  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[19]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b2  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[2]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b20  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[20]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b21  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[21]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b22  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[22]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b23  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[23]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b24  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[24]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b25  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[25]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b26  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[26]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b27  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[27]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b28  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[28]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b29  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[29]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b3  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[3]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b30  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[30]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b31  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[31]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b32  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [32]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[32]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b33  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [33]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[33]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b34  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [34]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[34]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b35  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [35]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[35]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b36  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [36]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[36]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b37  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [37]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[37]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b38  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [38]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[38]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b39  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [39]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[39]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b4  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[4]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b40  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [40]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[40]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b41  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [41]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[41]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b42  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [42]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[42]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b43  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [43]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[43]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b44  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [44]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[44]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b45  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [45]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[45]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b46  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [46]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[46]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b47  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [47]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[47]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b48  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [48]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[48]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b49  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [49]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[49]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b5  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[5]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b50  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [50]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[50]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b51  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [51]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[51]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b52  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [52]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[52]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b53  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [53]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[53]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b54  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [54]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[54]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b55  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [55]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[55]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b56  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [56]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[56]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b57  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [57]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[57]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b58  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [58]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[58]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b59  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [59]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[59]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b6  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[6]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b60  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [60]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[60]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b61  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [61]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[61]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b62  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [62]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[62]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b63  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [63]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[63]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b7  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[7]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b8  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[8]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b9  (
    .clk(clk_pad),
    .d(\ins_dec/n284 [9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[9]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b0  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[0]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b1  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[1]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b10  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[10]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b11  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[11]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b12  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[12]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b13  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[13]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b14  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[14]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b15  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[15]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b16  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[16]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b17  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[17]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b18  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[18]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b19  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[19]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b2  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[2]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b20  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[20]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b21  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[21]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b22  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[22]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b23  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[23]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b24  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[24]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b25  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[25]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b26  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[26]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b27  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[27]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b28  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[28]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b29  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[29]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b3  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[3]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b30  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[30]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b31  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[31]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b32  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [32]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[32]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b33  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [33]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[33]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b34  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [34]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[34]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b35  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [35]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[35]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b36  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [36]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[36]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b37  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [37]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[37]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b38  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [38]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[38]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b39  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [39]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[39]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b4  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[4]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b40  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [40]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[40]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b41  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [41]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[41]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b42  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [42]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[42]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b43  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [43]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[43]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b44  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [44]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[44]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b45  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [45]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[45]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b46  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [46]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[46]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b47  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [47]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[47]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b48  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [48]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[48]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b49  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [49]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[49]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b5  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[5]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b50  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [50]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[50]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b51  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [51]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[51]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b52  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [52]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[52]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b53  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [53]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[53]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b54  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [54]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[54]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b55  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [55]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[55]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b56  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [56]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[56]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b57  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [57]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[57]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b58  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [58]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[58]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b59  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [59]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[59]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b6  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[6]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b60  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [60]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[60]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b61  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [61]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[61]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b62  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [62]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[62]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b63  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [63]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[63]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b7  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[7]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b8  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[8]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b9  (
    .clk(clk_pad),
    .d(\ins_dec/n286 [9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[9]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b0  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[0]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b1  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[1]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b10  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[10]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b11  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[11]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b12  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[12]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b13  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[13]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b14  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[14]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b15  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[15]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b16  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[16]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b17  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[17]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b18  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[18]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b19  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[19]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b2  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[2]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b20  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[20]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b3  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[3]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b4  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[4]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b5  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[5]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b56  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [56]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[56]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b6  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[6]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b7  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[7]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b8  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[8]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b9  (
    .clk(clk_pad),
    .d(\ins_dec/n291 [9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[9]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b0  (
    .clk(clk_pad),
    .d(\ins_dec/op_count_decode [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[0]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b1  (
    .clk(clk_pad),
    .d(\ins_dec/op_count_decode [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[1]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b2  (
    .clk(clk_pad),
    .d(\ins_dec/op_count_decode [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[2]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b3  (
    .clk(clk_pad),
    .d(\ins_dec/op_count_decode [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[3]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b4  (
    .clk(clk_pad),
    .d(\ins_dec/op_count_decode [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[4]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b5  (
    .clk(clk_pad),
    .d(\ins_dec/op_count_decode [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[5]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b6  (
    .clk(clk_pad),
    .d(\ins_dec/op_count_decode [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[6]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b7  (
    .clk(clk_pad),
    .d(\ins_dec/op_count_decode [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[7]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/s_ret_reg  (
    .clk(clk_pad),
    .d(1'b0),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_s_ret));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/shift_l_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n235 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(shift_l));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/shift_r_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n232 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(shift_r));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/store_reg  (
    .clk(clk_pad),
    .d(\ins_dec/op_store ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(store));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/unsign_reg  (
    .clk(clk_pad),
    .d(\ins_dec/n206 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(unsign));  // ../../RTL/CPU/ID/ins_dec.v(674)
  reg_sr_as_w1 \ins_dec/valid_reg  (
    .clk(clk_pad),
    .d(id_valid),
    .en(~id_hold),
    .reset(~\ins_dec/u478_sel_is_0_o ),
    .set(1'b0),
    .q(ex_valid));  // ../../RTL/CPU/ID/ins_dec.v(830)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u0  (
    .a(addr_if[2]),
    .b(1'b1),
    .c(\ins_fetch/add0/c0 ),
    .o({\ins_fetch/add0/c1 ,\ins_fetch/n1 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u1  (
    .a(addr_if[3]),
    .b(1'b0),
    .c(\ins_fetch/add0/c1 ),
    .o({\ins_fetch/add0/c2 ,\ins_fetch/n1 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u10  (
    .a(addr_if[12]),
    .b(1'b0),
    .c(\ins_fetch/add0/c10 ),
    .o({\ins_fetch/add0/c11 ,\ins_fetch/n1 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u11  (
    .a(addr_if[13]),
    .b(1'b0),
    .c(\ins_fetch/add0/c11 ),
    .o({\ins_fetch/add0/c12 ,\ins_fetch/n1 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u12  (
    .a(addr_if[14]),
    .b(1'b0),
    .c(\ins_fetch/add0/c12 ),
    .o({\ins_fetch/add0/c13 ,\ins_fetch/n1 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u13  (
    .a(addr_if[15]),
    .b(1'b0),
    .c(\ins_fetch/add0/c13 ),
    .o({\ins_fetch/add0/c14 ,\ins_fetch/n1 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u14  (
    .a(addr_if[16]),
    .b(1'b0),
    .c(\ins_fetch/add0/c14 ),
    .o({\ins_fetch/add0/c15 ,\ins_fetch/n1 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u15  (
    .a(addr_if[17]),
    .b(1'b0),
    .c(\ins_fetch/add0/c15 ),
    .o({\ins_fetch/add0/c16 ,\ins_fetch/n1 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u16  (
    .a(addr_if[18]),
    .b(1'b0),
    .c(\ins_fetch/add0/c16 ),
    .o({\ins_fetch/add0/c17 ,\ins_fetch/n1 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u17  (
    .a(addr_if[19]),
    .b(1'b0),
    .c(\ins_fetch/add0/c17 ),
    .o({\ins_fetch/add0/c18 ,\ins_fetch/n1 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u18  (
    .a(addr_if[20]),
    .b(1'b0),
    .c(\ins_fetch/add0/c18 ),
    .o({\ins_fetch/add0/c19 ,\ins_fetch/n1 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u19  (
    .a(addr_if[21]),
    .b(1'b0),
    .c(\ins_fetch/add0/c19 ),
    .o({\ins_fetch/add0/c20 ,\ins_fetch/n1 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u2  (
    .a(addr_if[4]),
    .b(1'b0),
    .c(\ins_fetch/add0/c2 ),
    .o({\ins_fetch/add0/c3 ,\ins_fetch/n1 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u20  (
    .a(addr_if[22]),
    .b(1'b0),
    .c(\ins_fetch/add0/c20 ),
    .o({\ins_fetch/add0/c21 ,\ins_fetch/n1 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u21  (
    .a(addr_if[23]),
    .b(1'b0),
    .c(\ins_fetch/add0/c21 ),
    .o({\ins_fetch/add0/c22 ,\ins_fetch/n1 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u22  (
    .a(addr_if[24]),
    .b(1'b0),
    .c(\ins_fetch/add0/c22 ),
    .o({\ins_fetch/add0/c23 ,\ins_fetch/n1 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u23  (
    .a(addr_if[25]),
    .b(1'b0),
    .c(\ins_fetch/add0/c23 ),
    .o({\ins_fetch/add0/c24 ,\ins_fetch/n1 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u24  (
    .a(addr_if[26]),
    .b(1'b0),
    .c(\ins_fetch/add0/c24 ),
    .o({\ins_fetch/add0/c25 ,\ins_fetch/n1 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u25  (
    .a(addr_if[27]),
    .b(1'b0),
    .c(\ins_fetch/add0/c25 ),
    .o({\ins_fetch/add0/c26 ,\ins_fetch/n1 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u26  (
    .a(addr_if[28]),
    .b(1'b0),
    .c(\ins_fetch/add0/c26 ),
    .o({\ins_fetch/add0/c27 ,\ins_fetch/n1 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u27  (
    .a(addr_if[29]),
    .b(1'b0),
    .c(\ins_fetch/add0/c27 ),
    .o({\ins_fetch/add0/c28 ,\ins_fetch/n1 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u28  (
    .a(addr_if[30]),
    .b(1'b0),
    .c(\ins_fetch/add0/c28 ),
    .o({\ins_fetch/add0/c29 ,\ins_fetch/n1 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u29  (
    .a(addr_if[31]),
    .b(1'b0),
    .c(\ins_fetch/add0/c29 ),
    .o({\ins_fetch/add0/c30 ,\ins_fetch/n1 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u3  (
    .a(addr_if[5]),
    .b(1'b0),
    .c(\ins_fetch/add0/c3 ),
    .o({\ins_fetch/add0/c4 ,\ins_fetch/n1 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u30  (
    .a(addr_if[32]),
    .b(1'b0),
    .c(\ins_fetch/add0/c30 ),
    .o({\ins_fetch/add0/c31 ,\ins_fetch/n1 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u31  (
    .a(addr_if[33]),
    .b(1'b0),
    .c(\ins_fetch/add0/c31 ),
    .o({\ins_fetch/add0/c32 ,\ins_fetch/n1 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u32  (
    .a(addr_if[34]),
    .b(1'b0),
    .c(\ins_fetch/add0/c32 ),
    .o({\ins_fetch/add0/c33 ,\ins_fetch/n1 [32]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u33  (
    .a(addr_if[35]),
    .b(1'b0),
    .c(\ins_fetch/add0/c33 ),
    .o({\ins_fetch/add0/c34 ,\ins_fetch/n1 [33]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u34  (
    .a(addr_if[36]),
    .b(1'b0),
    .c(\ins_fetch/add0/c34 ),
    .o({\ins_fetch/add0/c35 ,\ins_fetch/n1 [34]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u35  (
    .a(addr_if[37]),
    .b(1'b0),
    .c(\ins_fetch/add0/c35 ),
    .o({\ins_fetch/add0/c36 ,\ins_fetch/n1 [35]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u36  (
    .a(addr_if[38]),
    .b(1'b0),
    .c(\ins_fetch/add0/c36 ),
    .o({\ins_fetch/add0/c37 ,\ins_fetch/n1 [36]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u37  (
    .a(addr_if[39]),
    .b(1'b0),
    .c(\ins_fetch/add0/c37 ),
    .o({\ins_fetch/add0/c38 ,\ins_fetch/n1 [37]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u38  (
    .a(addr_if[40]),
    .b(1'b0),
    .c(\ins_fetch/add0/c38 ),
    .o({\ins_fetch/add0/c39 ,\ins_fetch/n1 [38]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u39  (
    .a(addr_if[41]),
    .b(1'b0),
    .c(\ins_fetch/add0/c39 ),
    .o({\ins_fetch/add0/c40 ,\ins_fetch/n1 [39]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u4  (
    .a(addr_if[6]),
    .b(1'b0),
    .c(\ins_fetch/add0/c4 ),
    .o({\ins_fetch/add0/c5 ,\ins_fetch/n1 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u40  (
    .a(addr_if[42]),
    .b(1'b0),
    .c(\ins_fetch/add0/c40 ),
    .o({\ins_fetch/add0/c41 ,\ins_fetch/n1 [40]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u41  (
    .a(addr_if[43]),
    .b(1'b0),
    .c(\ins_fetch/add0/c41 ),
    .o({\ins_fetch/add0/c42 ,\ins_fetch/n1 [41]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u42  (
    .a(addr_if[44]),
    .b(1'b0),
    .c(\ins_fetch/add0/c42 ),
    .o({\ins_fetch/add0/c43 ,\ins_fetch/n1 [42]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u43  (
    .a(addr_if[45]),
    .b(1'b0),
    .c(\ins_fetch/add0/c43 ),
    .o({\ins_fetch/add0/c44 ,\ins_fetch/n1 [43]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u44  (
    .a(addr_if[46]),
    .b(1'b0),
    .c(\ins_fetch/add0/c44 ),
    .o({\ins_fetch/add0/c45 ,\ins_fetch/n1 [44]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u45  (
    .a(addr_if[47]),
    .b(1'b0),
    .c(\ins_fetch/add0/c45 ),
    .o({\ins_fetch/add0/c46 ,\ins_fetch/n1 [45]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u46  (
    .a(addr_if[48]),
    .b(1'b0),
    .c(\ins_fetch/add0/c46 ),
    .o({\ins_fetch/add0/c47 ,\ins_fetch/n1 [46]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u47  (
    .a(addr_if[49]),
    .b(1'b0),
    .c(\ins_fetch/add0/c47 ),
    .o({\ins_fetch/add0/c48 ,\ins_fetch/n1 [47]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u48  (
    .a(addr_if[50]),
    .b(1'b0),
    .c(\ins_fetch/add0/c48 ),
    .o({\ins_fetch/add0/c49 ,\ins_fetch/n1 [48]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u49  (
    .a(addr_if[51]),
    .b(1'b0),
    .c(\ins_fetch/add0/c49 ),
    .o({\ins_fetch/add0/c50 ,\ins_fetch/n1 [49]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u5  (
    .a(addr_if[7]),
    .b(1'b0),
    .c(\ins_fetch/add0/c5 ),
    .o({\ins_fetch/add0/c6 ,\ins_fetch/n1 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u50  (
    .a(addr_if[52]),
    .b(1'b0),
    .c(\ins_fetch/add0/c50 ),
    .o({\ins_fetch/add0/c51 ,\ins_fetch/n1 [50]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u51  (
    .a(addr_if[53]),
    .b(1'b0),
    .c(\ins_fetch/add0/c51 ),
    .o({\ins_fetch/add0/c52 ,\ins_fetch/n1 [51]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u52  (
    .a(addr_if[54]),
    .b(1'b0),
    .c(\ins_fetch/add0/c52 ),
    .o({\ins_fetch/add0/c53 ,\ins_fetch/n1 [52]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u53  (
    .a(addr_if[55]),
    .b(1'b0),
    .c(\ins_fetch/add0/c53 ),
    .o({\ins_fetch/add0/c54 ,\ins_fetch/n1 [53]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u54  (
    .a(addr_if[56]),
    .b(1'b0),
    .c(\ins_fetch/add0/c54 ),
    .o({\ins_fetch/add0/c55 ,\ins_fetch/n1 [54]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u55  (
    .a(addr_if[57]),
    .b(1'b0),
    .c(\ins_fetch/add0/c55 ),
    .o({\ins_fetch/add0/c56 ,\ins_fetch/n1 [55]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u56  (
    .a(addr_if[58]),
    .b(1'b0),
    .c(\ins_fetch/add0/c56 ),
    .o({\ins_fetch/add0/c57 ,\ins_fetch/n1 [56]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u57  (
    .a(addr_if[59]),
    .b(1'b0),
    .c(\ins_fetch/add0/c57 ),
    .o({\ins_fetch/add0/c58 ,\ins_fetch/n1 [57]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u58  (
    .a(addr_if[60]),
    .b(1'b0),
    .c(\ins_fetch/add0/c58 ),
    .o({\ins_fetch/add0/c59 ,\ins_fetch/n1 [58]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u59  (
    .a(addr_if[61]),
    .b(1'b0),
    .c(\ins_fetch/add0/c59 ),
    .o({\ins_fetch/add0/c60 ,\ins_fetch/n1 [59]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u6  (
    .a(addr_if[8]),
    .b(1'b0),
    .c(\ins_fetch/add0/c6 ),
    .o({\ins_fetch/add0/c7 ,\ins_fetch/n1 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u60  (
    .a(addr_if[62]),
    .b(1'b0),
    .c(\ins_fetch/add0/c60 ),
    .o({\ins_fetch/add0/c61 ,\ins_fetch/n1 [60]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u61  (
    .a(addr_if[63]),
    .b(1'b0),
    .c(\ins_fetch/add0/c61 ),
    .o({open_n6284,\ins_fetch/n1 [61]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u7  (
    .a(addr_if[9]),
    .b(1'b0),
    .c(\ins_fetch/add0/c7 ),
    .o({\ins_fetch/add0/c8 ,\ins_fetch/n1 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u8  (
    .a(addr_if[10]),
    .b(1'b0),
    .c(\ins_fetch/add0/c8 ),
    .o({\ins_fetch/add0/c9 ,\ins_fetch/n1 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \ins_fetch/add0/u9  (
    .a(addr_if[11]),
    .b(1'b0),
    .c(\ins_fetch/add0/c9 ),
    .o({\ins_fetch/add0/c10 ,\ins_fetch/n1 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \ins_fetch/add0/ucin  (
    .a(1'b0),
    .o({\ins_fetch/add0/c0 ,open_n6287}));
  reg_sr_as_w1 \ins_fetch/hold_reg  (
    .clk(clk_pad),
    .d(if_hold),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/hold ));  // ../../RTL/CPU/IF/ins_fetch.v(115)
  reg_sr_as_w1 \ins_fetch/ins_acc_fault_reg  (
    .clk(clk_pad),
    .d(ins_acc_fault),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_acc_fault));  // ../../RTL/CPU/IF/ins_fetch.v(137)
  reg_sr_as_w1 \ins_fetch/ins_addr_mis_reg  (
    .clk(clk_pad),
    .d(\ins_fetch/addr_mis ),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_addr_mis));  // ../../RTL/CPU/IF/ins_fetch.v(137)
  reg_sr_as_w1 \ins_fetch/ins_page_fault_reg  (
    .clk(clk_pad),
    .d(ins_page_fault),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_page_fault));  // ../../RTL/CPU/IF/ins_fetch.v(137)
  reg_sr_as_w1 \ins_fetch/int_acc_reg  (
    .clk(clk_pad),
    .d(int_req),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_int_acc));  // ../../RTL/CPU/IF/ins_fetch.v(137)
  reg_sr_as_w1 \ins_fetch/reg0_b0  (
    .clk(clk_pad),
    .d(addr_if[0]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[0]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b1  (
    .clk(clk_pad),
    .d(addr_if[1]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[1]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b10  (
    .clk(clk_pad),
    .d(addr_if[10]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[10]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b11  (
    .clk(clk_pad),
    .d(addr_if[11]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[11]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b12  (
    .clk(clk_pad),
    .d(addr_if[12]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[12]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b13  (
    .clk(clk_pad),
    .d(addr_if[13]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[13]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b14  (
    .clk(clk_pad),
    .d(addr_if[14]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[14]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b15  (
    .clk(clk_pad),
    .d(addr_if[15]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[15]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b16  (
    .clk(clk_pad),
    .d(addr_if[16]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[16]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b17  (
    .clk(clk_pad),
    .d(addr_if[17]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[17]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b18  (
    .clk(clk_pad),
    .d(addr_if[18]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[18]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b19  (
    .clk(clk_pad),
    .d(addr_if[19]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[19]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b2  (
    .clk(clk_pad),
    .d(addr_if[2]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[2]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b20  (
    .clk(clk_pad),
    .d(addr_if[20]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[20]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b21  (
    .clk(clk_pad),
    .d(addr_if[21]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[21]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b22  (
    .clk(clk_pad),
    .d(addr_if[22]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[22]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b23  (
    .clk(clk_pad),
    .d(addr_if[23]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[23]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b24  (
    .clk(clk_pad),
    .d(addr_if[24]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[24]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b25  (
    .clk(clk_pad),
    .d(addr_if[25]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[25]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b26  (
    .clk(clk_pad),
    .d(addr_if[26]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[26]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b27  (
    .clk(clk_pad),
    .d(addr_if[27]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[27]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b28  (
    .clk(clk_pad),
    .d(addr_if[28]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[28]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b29  (
    .clk(clk_pad),
    .d(addr_if[29]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[29]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b3  (
    .clk(clk_pad),
    .d(addr_if[3]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[3]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b30  (
    .clk(clk_pad),
    .d(addr_if[30]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[30]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b31  (
    .clk(clk_pad),
    .d(addr_if[31]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[31]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b32  (
    .clk(clk_pad),
    .d(addr_if[32]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[32]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b33  (
    .clk(clk_pad),
    .d(addr_if[33]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[33]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b34  (
    .clk(clk_pad),
    .d(addr_if[34]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[34]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b35  (
    .clk(clk_pad),
    .d(addr_if[35]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[35]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b36  (
    .clk(clk_pad),
    .d(addr_if[36]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[36]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b37  (
    .clk(clk_pad),
    .d(addr_if[37]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[37]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b38  (
    .clk(clk_pad),
    .d(addr_if[38]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[38]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b39  (
    .clk(clk_pad),
    .d(addr_if[39]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[39]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b4  (
    .clk(clk_pad),
    .d(addr_if[4]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[4]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b40  (
    .clk(clk_pad),
    .d(addr_if[40]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[40]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b41  (
    .clk(clk_pad),
    .d(addr_if[41]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[41]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b42  (
    .clk(clk_pad),
    .d(addr_if[42]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[42]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b43  (
    .clk(clk_pad),
    .d(addr_if[43]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[43]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b44  (
    .clk(clk_pad),
    .d(addr_if[44]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[44]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b45  (
    .clk(clk_pad),
    .d(addr_if[45]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[45]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b46  (
    .clk(clk_pad),
    .d(addr_if[46]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[46]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b47  (
    .clk(clk_pad),
    .d(addr_if[47]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[47]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b48  (
    .clk(clk_pad),
    .d(addr_if[48]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[48]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b49  (
    .clk(clk_pad),
    .d(addr_if[49]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[49]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b5  (
    .clk(clk_pad),
    .d(addr_if[5]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[5]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b50  (
    .clk(clk_pad),
    .d(addr_if[50]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[50]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b51  (
    .clk(clk_pad),
    .d(addr_if[51]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[51]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b52  (
    .clk(clk_pad),
    .d(addr_if[52]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[52]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b53  (
    .clk(clk_pad),
    .d(addr_if[53]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[53]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b54  (
    .clk(clk_pad),
    .d(addr_if[54]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[54]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b55  (
    .clk(clk_pad),
    .d(addr_if[55]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[55]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b56  (
    .clk(clk_pad),
    .d(addr_if[56]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[56]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b57  (
    .clk(clk_pad),
    .d(addr_if[57]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[57]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b58  (
    .clk(clk_pad),
    .d(addr_if[58]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[58]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b59  (
    .clk(clk_pad),
    .d(addr_if[59]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[59]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b6  (
    .clk(clk_pad),
    .d(addr_if[6]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[6]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b60  (
    .clk(clk_pad),
    .d(addr_if[60]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[60]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b61  (
    .clk(clk_pad),
    .d(addr_if[61]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[61]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b62  (
    .clk(clk_pad),
    .d(addr_if[62]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[62]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b63  (
    .clk(clk_pad),
    .d(addr_if[63]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[63]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b7  (
    .clk(clk_pad),
    .d(addr_if[7]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[7]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b8  (
    .clk(clk_pad),
    .d(addr_if[8]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[8]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b9  (
    .clk(clk_pad),
    .d(addr_if[9]),
    .en(~if_hold),
    .reset(rst_pad),
    .set(1'b0),
    .q(id_ins_pc[9]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg1_b0  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [0]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [0]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b1  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [1]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [1]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b10  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [10]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [10]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b11  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [11]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [11]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b12  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [12]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [12]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b13  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [13]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [13]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b14  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [14]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [14]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b15  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [15]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [15]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b16  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [16]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [16]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b17  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [17]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [17]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b18  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [18]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [18]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b19  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [19]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [19]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b2  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [2]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [2]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b20  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [20]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [20]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b21  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [21]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [21]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b22  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [22]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [22]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b23  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [23]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [23]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b24  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [24]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [24]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b25  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [25]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [25]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b26  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [26]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [26]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b27  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [27]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [27]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b28  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [28]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [28]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b29  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [29]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [29]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b3  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [3]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [3]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b30  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [30]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [30]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b31  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [31]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [31]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b4  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [4]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [4]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b5  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [5]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [5]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b6  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [6]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [6]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b7  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [7]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [7]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b8  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [8]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [8]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b9  (
    .clk(clk_pad),
    .d(\ins_fetch/ins_shift [9]),
    .en(\ins_fetch/n9 ),
    .reset(rst_pad),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [9]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg2_b0  (
    .clk(clk_pad),
    .d(flush_pc[0]),
    .en(pip_flush),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[0]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b1  (
    .clk(clk_pad),
    .d(flush_pc[1]),
    .en(pip_flush),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[1]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b10  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [10]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[10]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b11  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [11]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[11]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b12  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [12]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[12]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b13  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [13]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[13]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b14  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [14]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[14]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b15  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [15]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[15]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b16  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [16]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[16]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b17  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [17]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[17]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b18  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [18]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[18]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b19  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [19]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[19]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b2  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [2]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[2]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b20  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [20]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[20]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b21  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [21]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[21]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b22  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [22]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[22]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b23  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [23]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[23]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b24  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [24]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[24]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b25  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [25]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[25]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b26  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [26]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[26]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b27  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [27]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[27]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b28  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [28]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[28]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b29  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [29]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[29]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b3  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [3]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[3]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b30  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [30]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[30]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b31  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [31]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[31]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b32  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [32]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[32]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b33  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [33]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[33]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b34  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [34]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[34]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b35  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [35]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[35]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b36  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [36]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[36]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b37  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [37]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[37]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b38  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [38]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[38]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b39  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [39]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[39]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b4  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [4]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[4]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b40  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [40]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[40]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b41  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [41]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[41]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b42  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [42]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[42]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b43  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [43]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[43]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b44  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [44]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[44]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b45  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [45]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[45]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b46  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [46]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[46]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b47  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [47]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[47]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b48  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [48]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[48]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b49  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [49]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[49]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b5  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [5]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[5]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b50  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [50]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[50]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b51  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [51]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[51]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b52  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [52]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[52]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b53  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [53]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[53]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b54  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [54]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[54]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b55  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [55]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[55]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b56  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [56]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[56]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b57  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [57]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[57]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b58  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [58]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[58]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b59  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [59]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[59]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b6  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [6]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[6]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b60  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [60]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[60]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b61  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [61]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[61]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b62  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [62]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[62]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b63  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [63]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[63]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b7  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [7]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[7]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b8  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [8]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[8]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b9  (
    .clk(clk_pad),
    .d(\ins_fetch/n4 [9]),
    .en(1'b1),
    .reset(rst_pad),
    .set(1'b0),
    .q(addr_if[9]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/valid_reg  (
    .clk(clk_pad),
    .d(\ins_fetch/n27 ),
    .en(_al_n0_en),
    .reset(\ins_fetch/n25 ),
    .set(1'b0),
    .q(id_valid));  // ../../RTL/CPU/IF/ins_fetch.v(154)

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module reg_ar_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(setout),
    .reset(reset),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

