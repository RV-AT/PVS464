// Verilog netlist created by TD v4.5.12562
// Wed Apr  8 15:21:42 2020

`timescale 1ns / 1ps
module prv464_top  // ../../RTL/CPU/prv464_top.v(15)
  (
  cacheability_block,
  clk,
  hrdata,
  hready,
  hreset_n,
  hresp,
  m_ext_int,
  m_soft_int,
  m_time_int,
  mtime,
  rst,
  s_ext_int,
  haddr,
  hburst,
  hmastlock,
  hprot,
  hsize,
  htrans,
  hwdata,
  hwrite
  );

  input [31:0] cacheability_block;  // ../../RTL/CPU/prv464_top.v(17)
  input clk;  // ../../RTL/CPU/prv464_top.v(19)
  input [63:0] hrdata;  // ../../RTL/CPU/prv464_top.v(34)
  input hready;  // ../../RTL/CPU/prv464_top.v(31)
  input hreset_n;  // ../../RTL/CPU/prv464_top.v(33)
  input hresp;  // ../../RTL/CPU/prv464_top.v(32)
  input m_ext_int;  // ../../RTL/CPU/prv464_top.v(39)
  input m_soft_int;  // ../../RTL/CPU/prv464_top.v(38)
  input m_time_int;  // ../../RTL/CPU/prv464_top.v(37)
  input [63:0] mtime;  // ../../RTL/CPU/prv464_top.v(42)
  input rst;  // ../../RTL/CPU/prv464_top.v(20)
  input s_ext_int;  // ../../RTL/CPU/prv464_top.v(40)
  output [63:0] haddr;  // ../../RTL/CPU/prv464_top.v(22)
  output [2:0] hburst;  // ../../RTL/CPU/prv464_top.v(25)
  output hmastlock;  // ../../RTL/CPU/prv464_top.v(28)
  output [3:0] hprot;  // ../../RTL/CPU/prv464_top.v(26)
  output [2:0] hsize;  // ../../RTL/CPU/prv464_top.v(24)
  output [1:0] htrans;  // ../../RTL/CPU/prv464_top.v(27)
  output [63:0] hwdata;  // ../../RTL/CPU/prv464_top.v(29)
  output hwrite;  // ../../RTL/CPU/prv464_top.v(23)

  wire [63:0] addr_ex;  // ../../RTL/CPU/prv464_top.v(74)
  wire [63:0] addr_if;  // ../../RTL/CPU/prv464_top.v(65)
  wire [63:0] as1;  // ../../RTL/CPU/prv464_top.v(155)
  wire [63:0] as2;  // ../../RTL/CPU/prv464_top.v(156)
  wire [8:0] \biu/bus_unit/addr_counter ;  // ../../RTL/CPU/BIU/bus_unit.v(117)
  wire [8:0] \biu/bus_unit/last_addr ;  // ../../RTL/CPU/BIU/bus_unit.v(118)
  wire [1:0] \biu/bus_unit/mmu/i ;  // ../../RTL/CPU/BIU/mmu.v(94)
  wire [8:0] \biu/bus_unit/mmu/n28 ;
  wire [8:0] \biu/bus_unit/mmu/n29 ;
  wire [2:0] \biu/bus_unit/mmu/n33 ;
  wire [3:0] \biu/bus_unit/mmu/n36 ;
  wire [2:0] \biu/bus_unit/mmu/n38 ;
  wire [2:0] \biu/bus_unit/mmu/n39 ;
  wire [3:0] \biu/bus_unit/mmu/n40 ;
  wire [3:0] \biu/bus_unit/mmu/n43 ;
  wire [3:0] \biu/bus_unit/mmu/n44 ;
  wire [3:0] \biu/bus_unit/mmu/n46 ;
  wire [3:0] \biu/bus_unit/mmu/n49 ;
  wire [3:0] \biu/bus_unit/mmu/n50 ;
  wire [3:0] \biu/bus_unit/mmu/n51 ;
  wire [3:0] \biu/bus_unit/mmu/n52 ;
  wire [3:0] \biu/bus_unit/mmu/n53 ;
  wire [3:0] \biu/bus_unit/mmu/n54 ;
  wire [3:0] \biu/bus_unit/mmu/n55 ;
  wire [3:0] \biu/bus_unit/mmu/n56 ;
  wire [1:0] \biu/bus_unit/mmu/n59 ;
  wire [63:0] \biu/bus_unit/mmu/n63 ;
  wire [63:0] \biu/bus_unit/mmu/n64 ;
  wire [63:0] \biu/bus_unit/mmu/n65 ;
  wire [63:0] \biu/bus_unit/mmu/n66 ;
  wire [63:0] \biu/bus_unit/mmu/n68 ;
  wire [63:0] \biu/bus_unit/mmu/n70 ;
  wire [63:0] \biu/bus_unit/mmu/n71 ;
  wire [63:0] \biu/bus_unit/mmu/n75 ;
  wire [63:0] \biu/bus_unit/mmu/n76 ;
  wire [63:0] \biu/bus_unit/mmu/n78 ;
  wire [63:0] \biu/bus_unit/mmu/n79 ;
  wire [3:0] \biu/bus_unit/mmu/statu ;  // ../../RTL/CPU/BIU/mmu.v(95)
  wire [8:0] \biu/bus_unit/mmu/va_vpn ;  // ../../RTL/CPU/BIU/mmu.v(102)
  wire [1:0] \biu/bus_unit/mmu_htrans ;  // ../../RTL/CPU/BIU/bus_unit.v(104)
  wire [63:0] \biu/bus_unit/mmu_hwdata ;  // ../../RTL/CPU/BIU/bus_unit.v(106)
  wire [4:0] \biu/bus_unit/n17 ;
  wire [4:0] \biu/bus_unit/n19 ;
  wire [3:0] \biu/bus_unit/n23 ;
  wire [4:0] \biu/bus_unit/n26 ;
  wire [4:0] \biu/bus_unit/n27 ;
  wire [4:0] \biu/bus_unit/n28 ;
  wire [4:0] \biu/bus_unit/n29 ;
  wire [4:0] \biu/bus_unit/n30 ;
  wire [4:0] \biu/bus_unit/n31 ;
  wire [4:0] \biu/bus_unit/n32 ;
  wire [4:0] \biu/bus_unit/n33 ;
  wire [4:0] \biu/bus_unit/n34 ;
  wire [4:0] \biu/bus_unit/n35 ;
  wire [8:0] \biu/bus_unit/n39 ;
  wire [60:0] \biu/bus_unit/n49 ;
  wire [1:0] \biu/bus_unit/n54 ;
  wire [1:0] \biu/bus_unit/n55 ;
  wire [1:0] \biu/bus_unit/n59 ;
  wire [3:0] \biu/bus_unit/n6 ;
  wire [4:0] \biu/bus_unit/statu ;  // ../../RTL/CPU/BIU/bus_unit.v(115)
  wire [8:0] \biu/cache_counter ;  // ../../RTL/CPU/BIU/biu.v(127)
  wire [7:0] \biu/cache_ctrl_logic/ex_bsel ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(167)
  wire [127:0] \biu/cache_ctrl_logic/l1d_pa ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(143)
  wire [63:0] \biu/cache_ctrl_logic/l1d_pte ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(147)
  wire [63:0] \biu/cache_ctrl_logic/l1d_va ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(142)
  wire [127:0] \biu/cache_ctrl_logic/l1i_pa ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(141)
  wire [63:0] \biu/cache_ctrl_logic/l1i_pte ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(146)
  wire [63:0] \biu/cache_ctrl_logic/l1i_va ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(140)
  wire [4:0] \biu/cache_ctrl_logic/n100 ;
  wire [4:0] \biu/cache_ctrl_logic/n114 ;
  wire [4:0] \biu/cache_ctrl_logic/n115 ;
  wire [4:0] \biu/cache_ctrl_logic/n116 ;
  wire [4:0] \biu/cache_ctrl_logic/n117 ;
  wire [4:0] \biu/cache_ctrl_logic/n118 ;
  wire [4:0] \biu/cache_ctrl_logic/n119 ;
  wire [4:0] \biu/cache_ctrl_logic/n120 ;
  wire [4:0] \biu/cache_ctrl_logic/n121 ;
  wire [4:0] \biu/cache_ctrl_logic/n122 ;
  wire [4:0] \biu/cache_ctrl_logic/n123 ;
  wire [4:0] \biu/cache_ctrl_logic/n124 ;
  wire [4:0] \biu/cache_ctrl_logic/n125 ;
  wire [4:0] \biu/cache_ctrl_logic/n126 ;
  wire [4:0] \biu/cache_ctrl_logic/n127 ;
  wire [4:0] \biu/cache_ctrl_logic/n128 ;
  wire [4:0] \biu/cache_ctrl_logic/n129 ;
  wire [4:0] \biu/cache_ctrl_logic/n130 ;
  wire [4:0] \biu/cache_ctrl_logic/n131 ;
  wire [4:0] \biu/cache_ctrl_logic/n132 ;
  wire [63:0] \biu/cache_ctrl_logic/n147 ;
  wire [63:0] \biu/cache_ctrl_logic/n158 ;
  wire [127:0] \biu/cache_ctrl_logic/n164 ;
  wire [63:0] \biu/cache_ctrl_logic/n165 ;
  wire [127:0] \biu/cache_ctrl_logic/n166 ;
  wire [6:0] \biu/cache_ctrl_logic/n181 ;
  wire [7:0] \biu/cache_ctrl_logic/n182 ;
  wire [4:0] \biu/cache_ctrl_logic/n184 ;
  wire [6:0] \biu/cache_ctrl_logic/n185 ;
  wire [5:0] \biu/cache_ctrl_logic/n186 ;
  wire [6:0] \biu/cache_ctrl_logic/n189 ;
  wire [4:0] \biu/cache_ctrl_logic/n190 ;
  wire [5:0] \biu/cache_ctrl_logic/n192 ;
  wire [2:0] \biu/cache_ctrl_logic/n193 ;
  wire [63:0] \biu/cache_ctrl_logic/n207 ;
  wire [63:0] \biu/cache_ctrl_logic/n208 ;
  wire [63:0] \biu/cache_ctrl_logic/n209 ;
  wire [63:0] \biu/cache_ctrl_logic/n210 ;
  wire [63:0] \biu/cache_ctrl_logic/n211 ;
  wire [63:0] \biu/cache_ctrl_logic/n212 ;
  wire [63:0] \biu/cache_ctrl_logic/n213 ;
  wire [63:0] \biu/cache_ctrl_logic/n214 ;
  wire [63:0] \biu/cache_ctrl_logic/n215 ;
  wire [63:0] \biu/cache_ctrl_logic/n216 ;
  wire [63:0] \biu/cache_ctrl_logic/n217 ;
  wire [63:0] \biu/cache_ctrl_logic/n218 ;
  wire [63:0] \biu/cache_ctrl_logic/n219 ;
  wire [63:0] \biu/cache_ctrl_logic/n220 ;
  wire [63:0] \biu/cache_ctrl_logic/n221 ;
  wire [63:0] \biu/cache_ctrl_logic/n222 ;
  wire [63:0] \biu/cache_ctrl_logic/n223 ;
  wire [63:0] \biu/cache_ctrl_logic/n228 ;
  wire [63:0] \biu/cache_ctrl_logic/n229 ;
  wire [63:0] \biu/cache_ctrl_logic/n230 ;
  wire [63:0] \biu/cache_ctrl_logic/n231 ;
  wire [63:0] \biu/cache_ctrl_logic/n232 ;
  wire [63:0] \biu/cache_ctrl_logic/n233 ;
  wire [3:0] \biu/cache_ctrl_logic/n60 ;
  wire [3:0] \biu/cache_ctrl_logic/n61 ;
  wire [4:0] \biu/cache_ctrl_logic/n70 ;
  wire [4:0] \biu/cache_ctrl_logic/n71 ;
  wire [4:0] \biu/cache_ctrl_logic/n72 ;
  wire [2:0] \biu/cache_ctrl_logic/n73 ;
  wire [3:0] \biu/cache_ctrl_logic/n80 ;
  wire [3:0] \biu/cache_ctrl_logic/n81 ;
  wire [3:0] \biu/cache_ctrl_logic/n82 ;
  wire [4:0] \biu/cache_ctrl_logic/n83 ;
  wire [4:0] \biu/cache_ctrl_logic/n84 ;
  wire [4:0] \biu/cache_ctrl_logic/n87 ;
  wire [4:0] \biu/cache_ctrl_logic/n88 ;
  wire [3:0] \biu/cache_ctrl_logic/n90 ;
  wire [4:0] \biu/cache_ctrl_logic/n91 ;
  wire [4:0] \biu/cache_ctrl_logic/n92 ;
  wire [3:0] \biu/cache_ctrl_logic/n95 ;
  wire [4:0] \biu/cache_ctrl_logic/n96 ;
  wire [4:0] \biu/cache_ctrl_logic/n99 ;
  wire [11:0] \biu/cache_ctrl_logic/off ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(165)
  wire [127:0] \biu/cache_ctrl_logic/pa_temp ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(136)
  wire [63:0] \biu/cache_ctrl_logic/pte_temp ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(145)
  wire [4:0] \biu/cache_ctrl_logic/statu ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(133)
  wire [1:0] \biu/ex_data_sel ;  // ../../RTL/CPU/BIU/biu.v(81)
  wire [8:0] \biu/l1d_addr ;  // ../../RTL/CPU/BIU/biu.v(96)
  wire [7:0] \biu/l1d_bsel ;  // ../../RTL/CPU/BIU/biu.v(85)
  wire [63:0] \biu/l1d_out ;  // ../../RTL/CPU/BIU/biu.v(92)
  wire [8:0] \biu/l1i_addr ;  // ../../RTL/CPU/BIU/biu.v(95)
  wire [7:0] \biu/l1i_bsel ;  // ../../RTL/CPU/BIU/biu.v(84)
  wire [63:0] \biu/l1i_in ;  // ../../RTL/CPU/BIU/biu.v(91)
  wire [63:0] \biu/maddress ;  // ../../RTL/CPU/BIU/biu.v(119)
  wire [8:0] \biu/n0 ;
  wire [63:0] \biu/n1 ;
  wire [1:0] \biu/opc ;  // ../../RTL/CPU/BIU/biu.v(109)
  wire [127:0] \biu/paddress ;  // ../../RTL/CPU/BIU/biu.v(120)
  wire [3:0] \biu/priv ;  // ../../RTL/CPU/BIU/biu.v(110)
  wire [63:0] \biu/write_data ;  // ../../RTL/CPU/BIU/biu.v(125)
  wire [63:0] csr_data;  // ../../RTL/CPU/prv464_top.v(54)
  wire [11:0] csr_index;  // ../../RTL/CPU/prv464_top.v(180)
  wire [63:0] \cu_ru/exc_cause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(138)
  wire [63:0] \cu_ru/int_cause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(137)
  wire [63:0] \cu_ru/m_cycle_event/n2 ;
  wire [63:0] \cu_ru/m_cycle_event/n3 ;
  wire [63:0] \cu_ru/m_cycle_event/n4 ;
  wire [63:0] \cu_ru/m_cycle_event/n9 ;
  wire [63:0] \cu_ru/m_s_cause/n4 ;
  wire [63:0] \cu_ru/m_s_cause/n5 ;
  wire [63:0] \cu_ru/m_s_cause/n6 ;
  wire [63:0] \cu_ru/m_s_cause/n7 ;
  wire [61:0] \cu_ru/m_s_epc/n0 ;
  wire [63:0] \cu_ru/m_s_epc/n1 ;
  wire [63:0] \cu_ru/m_s_epc/n10 ;
  wire [63:0] \cu_ru/m_s_epc/n2 ;
  wire [63:0] \cu_ru/m_s_epc/n7 ;
  wire [63:0] \cu_ru/m_s_epc/n8 ;
  wire [63:0] \cu_ru/m_s_epc/n9 ;
  wire [1:0] \cu_ru/m_s_status/n21 ;
  wire [1:0] \cu_ru/m_s_status/n24 ;
  wire [1:0] \cu_ru/m_s_status/n35 ;
  wire [1:0] \cu_ru/m_s_status/n4 ;
  wire [1:0] \cu_ru/m_s_status/n47 ;
  wire [1:0] \cu_ru/m_s_status/n5 ;
  wire [1:0] \cu_ru/m_s_status/n6 ;
  wire [1:0] \cu_ru/m_s_status/n60 ;
  wire [3:0] \cu_ru/m_s_status/n61 ;
  wire [1:0] \cu_ru/m_s_status/n62 ;
  wire [3:0] \cu_ru/m_s_status/n63 ;
  wire [3:0] \cu_ru/m_s_status/n64 ;
  wire [63:0] \cu_ru/m_s_tval/n10 ;
  wire [63:0] \cu_ru/m_s_tval/n11 ;
  wire [63:0] \cu_ru/m_s_tval/n3 ;
  wire [63:0] \cu_ru/m_s_tval/n8 ;
  wire [63:0] \cu_ru/m_s_tval/n9 ;
  wire [63:0] \cu_ru/m_s_tvec/n7 ;
  wire [63:0] \cu_ru/m_sie ;  // ../../RTL/CPU/CU&RU/cu_ru.v(157)
  wire [63:0] \cu_ru/m_sip ;  // ../../RTL/CPU/CU&RU/cu_ru.v(158)
  wire [63:0] \cu_ru/mcause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(161)
  wire [63:0] \cu_ru/mcycle ;  // ../../RTL/CPU/CU&RU/cu_ru.v(170)
  wire [63:0] \cu_ru/medeleg ;  // ../../RTL/CPU/CU&RU/cu_ru.v(156)
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n91 ;
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n93 ;
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n94 ;
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n95 ;
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n97 ;
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n98 ;
  wire [3:0] \cu_ru/medeleg_exc_ctrl/n99 ;
  wire [63:0] \cu_ru/mepc ;  // ../../RTL/CPU/CU&RU/cu_ru.v(163)
  wire [63:0] \cu_ru/mideleg ;  // ../../RTL/CPU/CU&RU/cu_ru.v(155)
  wire [63:0] \cu_ru/mideleg_int_ctrl/n37 ;
  wire [63:0] \cu_ru/mideleg_int_ctrl/n38 ;
  wire [63:0] \cu_ru/minstret ;  // ../../RTL/CPU/CU&RU/cu_ru.v(171)
  wire [63:0] \cu_ru/mscratch ;  // ../../RTL/CPU/CU&RU/cu_ru.v(172)
  wire [63:0] \cu_ru/mstatus ;  // ../../RTL/CPU/CU&RU/cu_ru.v(153)
  wire [63:0] \cu_ru/mtval ;  // ../../RTL/CPU/CU&RU/cu_ru.v(165)
  wire [63:0] \cu_ru/mtvec ;  // ../../RTL/CPU/CU&RU/cu_ru.v(167)
  wire [63:0] \cu_ru/n100 ;
  wire [63:0] \cu_ru/n101 ;
  wire [63:0] \cu_ru/n102 ;
  wire [63:0] \cu_ru/n103 ;
  wire [63:0] \cu_ru/n104 ;
  wire [63:0] \cu_ru/n105 ;
  wire [63:0] \cu_ru/n106 ;
  wire [63:0] \cu_ru/n107 ;
  wire [63:0] \cu_ru/n108 ;
  wire [63:0] \cu_ru/n109 ;
  wire [63:0] \cu_ru/n110 ;
  wire [63:0] \cu_ru/n111 ;
  wire [63:0] \cu_ru/n112 ;
  wire [63:0] \cu_ru/n113 ;
  wire [63:0] \cu_ru/n114 ;
  wire [63:0] \cu_ru/n115 ;
  wire [61:0] \cu_ru/n43 ;
  wire [4:0] \cu_ru/n46 ;
  wire [63:0] \cu_ru/n47 ;
  wire [4:0] \cu_ru/n49 ;
  wire [63:0] \cu_ru/n50 ;
  wire [4:0] \cu_ru/n52 ;
  wire [63:0] \cu_ru/n57 ;
  wire [63:0] \cu_ru/n58 ;
  wire [63:0] \cu_ru/n59 ;
  wire [63:0] \cu_ru/n60 ;
  wire [63:0] \cu_ru/n61 ;
  wire [63:0] \cu_ru/n62 ;
  wire [63:0] \cu_ru/n63 ;
  wire [63:0] \cu_ru/n64 ;
  wire [63:0] \cu_ru/n65 ;
  wire [63:0] \cu_ru/n67 ;
  wire [63:0] \cu_ru/n68 ;
  wire [63:0] \cu_ru/n69 ;
  wire [63:0] \cu_ru/n70 ;
  wire [63:0] \cu_ru/n71 ;
  wire [63:0] \cu_ru/n72 ;
  wire [63:0] \cu_ru/n73 ;
  wire [63:0] \cu_ru/n74 ;
  wire [63:0] \cu_ru/n75 ;
  wire [63:0] \cu_ru/n76 ;
  wire [63:0] \cu_ru/n77 ;
  wire [63:0] \cu_ru/n78 ;
  wire [63:0] \cu_ru/n79 ;
  wire [63:0] \cu_ru/n80 ;
  wire [63:0] \cu_ru/n81 ;
  wire [63:0] \cu_ru/n82 ;
  wire [63:0] \cu_ru/n83 ;
  wire [63:0] \cu_ru/n84 ;
  wire [63:0] \cu_ru/n85 ;
  wire [63:0] \cu_ru/n86 ;
  wire [63:0] \cu_ru/n87 ;
  wire [63:0] \cu_ru/n90 ;
  wire [63:0] \cu_ru/n91 ;
  wire [63:0] \cu_ru/n94 ;
  wire [63:0] \cu_ru/n95 ;
  wire [63:0] \cu_ru/n96 ;
  wire [63:0] \cu_ru/n97 ;
  wire [63:0] \cu_ru/n99 ;
  wire [63:0] \cu_ru/scause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(162)
  wire [63:0] \cu_ru/sepc ;  // ../../RTL/CPU/CU&RU/cu_ru.v(164)
  wire [63:0] \cu_ru/sscratch ;  // ../../RTL/CPU/CU&RU/cu_ru.v(173)
  wire [63:0] \cu_ru/stval ;  // ../../RTL/CPU/CU&RU/cu_ru.v(166)
  wire [63:0] \cu_ru/stvec ;  // ../../RTL/CPU/CU&RU/cu_ru.v(168)
  wire [63:0] \cu_ru/trap_cause ;  // ../../RTL/CPU/CU&RU/cu_ru.v(131)
  wire [63:0] \cu_ru/tvec ;  // ../../RTL/CPU/CU&RU/cu_ru.v(133)
  wire [63:0] \cu_ru/vec_pc ;  // ../../RTL/CPU/CU&RU/cu_ru.v(135)
  wire [63:0] data_csr;  // ../../RTL/CPU/prv464_top.v(182)
  wire [63:0] data_rd;  // ../../RTL/CPU/prv464_top.v(183)
  wire [63:0] data_read;  // ../../RTL/CPU/prv464_top.v(75)
  wire [63:0] ds1;  // ../../RTL/CPU/prv464_top.v(153)
  wire [63:0] ds2;  // ../../RTL/CPU/prv464_top.v(154)
  wire [11:0] ex_csr_index;  // ../../RTL/CPU/prv464_top.v(147)
  wire [63:0] ex_exc_code;  // ../../RTL/CPU/prv464_top.v(99)
  wire [63:0] ex_ins_pc;  // ../../RTL/CPU/prv464_top.v(100)
  wire [3:0] ex_priv;  // ../../RTL/CPU/prv464_top.v(73)
  wire [4:0] ex_rd_index;  // ../../RTL/CPU/prv464_top.v(150)
  wire [3:0] ex_size;  // ../../RTL/CPU/prv464_top.v(133)
  wire [63:0] \exu/alu_au/add_64 ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(55)
  wire [63:0] \exu/alu_au/alu_add ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(54)
  wire [63:0] \exu/alu_au/alu_and ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(58)
  wire [63:0] \exu/alu_au/alu_max ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(64)
  wire [63:0] \exu/alu_au/alu_min ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(65)
  wire [63:0] \exu/alu_au/alu_or ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(59)
  wire [63:0] \exu/alu_au/alu_sub ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(57)
  wire [63:0] \exu/alu_au/alu_xor ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(60)
  wire [63:0] \exu/alu_au/n16 ;
  wire [63:0] \exu/alu_au/n17 ;
  wire [63:0] \exu/alu_au/n18 ;
  wire [63:0] \exu/alu_au/n28 ;
  wire [63:0] \exu/alu_au/n29 ;
  wire [63:0] \exu/alu_au/n30 ;
  wire [63:0] \exu/alu_au/n31 ;
  wire [63:0] \exu/alu_au/n32 ;
  wire [63:0] \exu/alu_au/n33 ;
  wire [63:0] \exu/alu_au/n34 ;
  wire [63:0] \exu/alu_au/n35 ;
  wire [63:0] \exu/alu_au/n36 ;
  wire [63:0] \exu/alu_au/n37 ;
  wire [63:0] \exu/alu_au/n38 ;
  wire [63:0] \exu/alu_au/n39 ;
  wire [63:0] \exu/alu_au/n40 ;
  wire [63:0] \exu/alu_au/n43 ;
  wire [63:0] \exu/alu_au/n45 ;
  wire [63:0] \exu/alu_au/n46 ;
  wire [63:0] \exu/alu_au/n47 ;
  wire [63:0] \exu/alu_au/n48 ;
  wire [63:0] \exu/alu_au/n49 ;
  wire [63:0] \exu/alu_au/n50 ;
  wire [63:0] \exu/alu_au/n51 ;
  wire [63:0] \exu/alu_au/n52 ;
  wire [63:0] \exu/alu_au/n53 ;
  wire [63:0] \exu/alu_au/n54 ;
  wire [63:0] \exu/alu_au/n55 ;
  wire [63:0] \exu/alu_au/sub_64 ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(56)
  wire [63:0] \exu/alu_data_mem_csr ;  // ../../RTL/CPU/EX/exu.v(193)
  wire [63:0] \exu/data_lsu_cache ;  // ../../RTL/CPU/EX/exu.v(197)
  wire [63:0] \exu/data_lsu_uncache ;  // ../../RTL/CPU/EX/exu.v(198)
  wire [63:0] \exu/lsu/data_lsu_cache_shift ;  // ../../RTL/CPU/EX/LSU/lsu.v(28)
  wire [63:0] \exu/lsu/data_lsu_uncache_shift ;  // ../../RTL/CPU/EX/LSU/lsu.v(29)
  wire [63:0] \exu/lsu/n1 ;
  wire [63:0] \exu/lsu/n10 ;
  wire [63:0] \exu/lsu/n22 ;
  wire [55:0] \exu/lsu/n23 ;
  wire [63:0] \exu/lsu/n24 ;
  wire [47:0] \exu/lsu/n25 ;
  wire [63:0] \exu/lsu/n26 ;
  wire [39:0] \exu/lsu/n27 ;
  wire [63:0] \exu/lsu/n28 ;
  wire [63:0] \exu/lsu/n3 ;
  wire [63:0] \exu/lsu/n36 ;
  wire [55:0] \exu/lsu/n37 ;
  wire [63:0] \exu/lsu/n38 ;
  wire [47:0] \exu/lsu/n39 ;
  wire [63:0] \exu/lsu/n4 ;
  wire [63:0] \exu/lsu/n40 ;
  wire [39:0] \exu/lsu/n41 ;
  wire [63:0] \exu/lsu/n42 ;
  wire [63:0] \exu/lsu/n52 ;
  wire [63:0] \exu/lsu/n54 ;
  wire [63:0] \exu/lsu/n55 ;
  wire [63:0] \exu/lsu/n57 ;
  wire [63:0] \exu/lsu/n58 ;
  wire [63:0] \exu/lsu/n59 ;
  wire [63:0] \exu/lsu/n6 ;
  wire [63:0] \exu/lsu/n60 ;
  wire [63:0] \exu/lsu/n61 ;
  wire [63:0] \exu/lsu/n62 ;
  wire [63:0] \exu/lsu/n63 ;
  wire [63:0] \exu/lsu/n64 ;
  wire [63:0] \exu/lsu/n65 ;
  wire [63:0] \exu/lsu/n7 ;
  wire [63:0] \exu/lsu/n9 ;
  wire [3:0] \exu/main_state ;  // ../../RTL/CPU/EX/exu.v(184)
  wire [3:0] \exu/n22 ;
  wire [3:0] \exu/n23 ;
  wire [3:0] \exu/n24 ;
  wire [3:0] \exu/n25 ;
  wire [3:0] \exu/n26 ;
  wire [1:0] \exu/n27 ;
  wire [2:0] \exu/n29 ;
  wire [3:0] \exu/n33 ;
  wire [3:0] \exu/n36 ;
  wire [3:0] \exu/n37 ;
  wire [3:0] \exu/n38 ;
  wire [3:0] \exu/n39 ;
  wire [3:0] \exu/n40 ;
  wire [3:0] \exu/n41 ;
  wire [3:0] \exu/n42 ;
  wire [3:0] \exu/n43 ;
  wire [3:0] \exu/n44 ;
  wire [3:0] \exu/n45 ;
  wire [7:0] \exu/n50 ;
  wire [7:0] \exu/n51 ;
  wire [7:0] \exu/n52 ;
  wire [31:0] \exu/n54 ;
  wire [64:0] \exu/n55 ;
  wire [32:0] \exu/n56 ;
  wire [63:0] \exu/n57 ;
  wire [63:0] \exu/n58 ;
  wire [63:0] \exu/n61 ;
  wire [63:0] \exu/n62 ;
  wire [63:0] \exu/n63 ;
  wire [63:0] \exu/n64 ;
  wire [63:0] \exu/n71 ;
  wire [7:0] \exu/shift_count ;  // ../../RTL/CPU/EX/exu.v(185)
  wire [63:0] flush_pc;  // ../../RTL/CPU/prv464_top.v(61)
  wire [31:0] id_ins;  // ../../RTL/CPU/prv464_top.v(90)
  wire [63:0] id_ins_pc;  // ../../RTL/CPU/prv464_top.v(91)
  wire [4:0] id_rs1_index;  // ../../RTL/CPU/prv464_top.v(57)
  wire [4:0] id_rs2_index;  // ../../RTL/CPU/prv464_top.v(59)
  wire [63:0] \ins_dec/n270 ;
  wire [63:0] \ins_dec/n271 ;
  wire [63:0] \ins_dec/n272 ;
  wire [63:0] \ins_dec/n280 ;
  wire [63:0] \ins_dec/n281 ;
  wire [63:0] \ins_dec/n282 ;
  wire [63:0] \ins_dec/n283 ;
  wire [63:0] \ins_dec/n284 ;
  wire [63:0] \ins_dec/n286 ;
  wire [63:0] \ins_dec/n287 ;
  wire [63:0] \ins_dec/n288 ;
  wire [63:0] \ins_dec/n289 ;
  wire [63:0] \ins_dec/n290 ;
  wire [63:0] \ins_dec/n291 ;
  wire [31:0] \ins_dec/n342 ;
  wire [7:0] \ins_dec/n58 ;
  wire [7:0] \ins_dec/op_count_decode ;  // ../../RTL/CPU/ID/ins_dec.v(239)
  wire [31:0] \ins_fetch/ins_hold ;  // ../../RTL/CPU/IF/ins_fetch.v(55)
  wire [31:0] \ins_fetch/ins_shift ;  // ../../RTL/CPU/IF/ins_fetch.v(59)
  wire [61:0] \ins_fetch/n1 ;
  wire [61:0] \ins_fetch/n3 ;
  wire [63:0] \ins_fetch/n4 ;
  wire [63:0] ins_read;  // ../../RTL/CPU/prv464_top.v(67)
  wire [3:0] mod_priv;  // ../../RTL/CPU/prv464_top.v(48)
  wire [63:0] new_pc;  // ../../RTL/CPU/prv464_top.v(184)
  wire [7:0] op_count;  // ../../RTL/CPU/prv464_top.v(157)
  wire [3:0] priv;  // ../../RTL/CPU/prv464_top.v(47)
  wire [63:0] rs1_data;  // ../../RTL/CPU/prv464_top.v(56)
  wire [63:0] rs2_data;  // ../../RTL/CPU/prv464_top.v(58)
  wire [63:0] satp;  // ../../RTL/CPU/prv464_top.v(46)
  wire [63:0] uncache_data;  // ../../RTL/CPU/prv464_top.v(77)
  wire [63:0] wb_exc_code;  // ../../RTL/CPU/prv464_top.v(185)
  wire [63:0] wb_ins_pc;  // ../../RTL/CPU/prv464_top.v(186)
  wire [4:0] wb_rd_index;  // ../../RTL/CPU/prv464_top.v(181)
  wire amo;  // ../../RTL/CPU/prv464_top.v(138)
  wire amo_neg;
  wire and_clr;  // ../../RTL/CPU/prv464_top.v(129)
  wire \biu/bus_error ;  // ../../RTL/CPU/BIU/biu.v(117)
  wire \biu/bus_error_neg ;
  wire \biu/bus_unit/mmu/leaf_page ;  // ../../RTL/CPU/BIU/mmu.v(99)
  wire \biu/bus_unit/mmu/mux10_b0_sel_is_2_o ;
  wire \biu/bus_unit/mmu/mux16_b2_sel_is_0_o ;
  wire \biu/bus_unit/mmu/mux17_b3_sel_is_0_o ;
  wire \biu/bus_unit/mmu/mux18_b3_sel_is_2_o ;
  wire \biu/bus_unit/mmu/mux20_b0_sel_is_3_o ;
  wire \biu/bus_unit/mmu/mux23_b0_sel_is_3_o ;
  wire \biu/bus_unit/mmu/mux23_b0_sel_is_3_o_neg ;
  wire \biu/bus_unit/mmu/mux24_b0_sel_is_1_o ;
  wire \biu/bus_unit/mmu/mux34_b0_sel_is_3_o ;
  wire \biu/bus_unit/mmu/mux6_b1_sel_is_0_o ;
  wire \biu/bus_unit/mmu/mux9_b0_sel_is_0_o ;
  wire \biu/bus_unit/mmu/n0 ;
  wire \biu/bus_unit/mmu/n1 ;
  wire \biu/bus_unit/mmu/n10 ;
  wire \biu/bus_unit/mmu/n11 ;
  wire \biu/bus_unit/mmu/n12 ;
  wire \biu/bus_unit/mmu/n13 ;
  wire \biu/bus_unit/mmu/n14 ;
  wire \biu/bus_unit/mmu/n15 ;
  wire \biu/bus_unit/mmu/n16 ;
  wire \biu/bus_unit/mmu/n17 ;
  wire \biu/bus_unit/mmu/n18 ;
  wire \biu/bus_unit/mmu/n19 ;
  wire \biu/bus_unit/mmu/n2 ;
  wire \biu/bus_unit/mmu/n20 ;
  wire \biu/bus_unit/mmu/n21 ;
  wire \biu/bus_unit/mmu/n22 ;
  wire \biu/bus_unit/mmu/n23 ;
  wire \biu/bus_unit/mmu/n24 ;
  wire \biu/bus_unit/mmu/n25 ;
  wire \biu/bus_unit/mmu/n26 ;
  wire \biu/bus_unit/mmu/n27 ;
  wire \biu/bus_unit/mmu/n3 ;
  wire \biu/bus_unit/mmu/n30 ;
  wire \biu/bus_unit/mmu/n30_neg ;
  wire \biu/bus_unit/mmu/n31 ;
  wire \biu/bus_unit/mmu/n32 ;
  wire \biu/bus_unit/mmu/n34 ;
  wire \biu/bus_unit/mmu/n34_neg ;
  wire \biu/bus_unit/mmu/n35 ;
  wire \biu/bus_unit/mmu/n35_neg ;
  wire \biu/bus_unit/mmu/n37 ;
  wire \biu/bus_unit/mmu/n4 ;
  wire \biu/bus_unit/mmu/n41 ;
  wire \biu/bus_unit/mmu/n42 ;
  wire \biu/bus_unit/mmu/n45 ;
  wire \biu/bus_unit/mmu/n5 ;
  wire \biu/bus_unit/mmu/n58 ;
  wire \biu/bus_unit/mmu/n6 ;
  wire \biu/bus_unit/mmu/n7 ;
  wire \biu/bus_unit/mmu/n73 ;
  wire \biu/bus_unit/mmu/n74 ;
  wire \biu/bus_unit/mmu/n77 ;
  wire \biu/bus_unit/mmu/n8 ;
  wire \biu/bus_unit/mmu/n81 ;
  wire \biu/bus_unit/mmu/n9 ;
  wire \biu/bus_unit/mmu/page_chk_ok ;  // ../../RTL/CPU/BIU/mmu.v(100)
  wire \biu/bus_unit/mmu/page_unvalid ;  // ../../RTL/CPU/BIU/mmu.v(97)
  wire \biu/bus_unit/mmu/page_unvalid_neg ;
  wire \biu/bus_unit/mmu/pointer_page ;  // ../../RTL/CPU/BIU/mmu.v(98)
  wire \biu/bus_unit/mmu/pointer_page_neg ;
  wire \biu/bus_unit/mmu_acc_fault ;  // ../../RTL/CPU/BIU/bus_unit.v(110)
  wire \biu/bus_unit/mmu_acc_fault_neg ;
  wire \biu/bus_unit/mmu_hwrite ;  // ../../RTL/CPU/BIU/bus_unit.v(100)
  wire \biu/bus_unit/mmu_page_fault ;  // ../../RTL/CPU/BIU/bus_unit.v(111)
  wire \biu/bus_unit/mmu_page_fault_neg ;
  wire \biu/bus_unit/mmu_trans_rdy ;  // ../../RTL/CPU/BIU/bus_unit.v(109)
  wire \biu/bus_unit/mmu_trans_rdy_neg ;
  wire \biu/bus_unit/mux10_b0_sel_is_2_o ;
  wire \biu/bus_unit/mux10_b3_sel_is_0_o ;
  wire \biu/bus_unit/mux11_b2_sel_is_0_o ;
  wire \biu/bus_unit/mux11_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux13_b0_sel_is_0_o ;
  wire \biu/bus_unit/mux14_b1_sel_is_0_o ;
  wire \biu/bus_unit/mux14_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux15_b2_sel_is_2_o ;
  wire \biu/bus_unit/mux15_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux16_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux17_b4_sel_is_2_o ;
  wire \biu/bus_unit/mux19_b0_sel_is_3_o ;
  wire \biu/bus_unit/mux1_b1_sel_is_0_o ;
  wire \biu/bus_unit/mux1_b2_sel_is_2_o ;
  wire \biu/bus_unit/mux24_b1_sel_is_0_o ;
  wire \biu/bus_unit/mux24_b1_sel_is_0_o_neg ;
  wire \biu/bus_unit/mux25_b1_sel_is_0_o ;
  wire \biu/bus_unit/mux26_b0_sel_is_0_o ;
  wire \biu/bus_unit/mux28_b0_sel_is_0_o ;
  wire \biu/bus_unit/mux2_b0_sel_is_0_o ;
  wire \biu/bus_unit/mux2_b1_sel_is_2_o ;
  wire \biu/bus_unit/mux2_b2_sel_is_2_o ;
  wire \biu/bus_unit/mux2_b3_sel_is_2_o ;
  wire \biu/bus_unit/mux9_b0_sel_is_0_o ;
  wire \biu/bus_unit/n0 ;
  wire \biu/bus_unit/n0_neg ;
  wire \biu/bus_unit/n1 ;
  wire \biu/bus_unit/n10 ;
  wire \biu/bus_unit/n11 ;
  wire \biu/bus_unit/n11_neg ;
  wire \biu/bus_unit/n12 ;
  wire \biu/bus_unit/n12_neg ;
  wire \biu/bus_unit/n13 ;
  wire \biu/bus_unit/n13_neg ;
  wire \biu/bus_unit/n14 ;
  wire \biu/bus_unit/n14_neg ;
  wire \biu/bus_unit/n15 ;
  wire \biu/bus_unit/n16 ;
  wire \biu/bus_unit/n18 ;
  wire \biu/bus_unit/n18_neg ;
  wire \biu/bus_unit/n1_neg ;
  wire \biu/bus_unit/n2 ;
  wire \biu/bus_unit/n20 ;
  wire \biu/bus_unit/n20_neg ;
  wire \biu/bus_unit/n22 ;
  wire \biu/bus_unit/n22_neg ;
  wire \biu/bus_unit/n25 ;
  wire \biu/bus_unit/n2_neg ;
  wire \biu/bus_unit/n3 ;
  wire \biu/bus_unit/n37 ;
  wire \biu/bus_unit/n38 ;
  wire \biu/bus_unit/n44 ;
  wire \biu/bus_unit/n45 ;
  wire \biu/bus_unit/n46 ;
  wire \biu/bus_unit/n47 ;
  wire \biu/bus_unit/n48 ;
  wire \biu/bus_unit/n50 ;
  wire \biu/bus_unit/n50_neg ;
  wire \biu/bus_unit/n51 ;
  wire \biu/bus_unit/n51_neg ;
  wire \biu/bus_unit/n52 ;
  wire \biu/bus_unit/n53 ;
  wire \biu/bus_unit/n56 ;
  wire \biu/bus_unit/n56_neg ;
  wire \biu/bus_unit/n58 ;
  wire \biu/bus_unit/n58_neg ;
  wire \biu/bus_unit/n60 ;
  wire \biu/bus_unit/n7 ;
  wire \biu/bus_unit/n7_neg ;
  wire \biu/bus_unit/n8 ;
  wire \biu/bus_unit/n9 ;
  wire \biu/cache/n1 ;
  wire \biu/cache/n11 ;
  wire \biu/cache/n13 ;
  wire \biu/cache/n15 ;
  wire \biu/cache/n17 ;
  wire \biu/cache/n19 ;
  wire \biu/cache/n21 ;
  wire \biu/cache/n23 ;
  wire \biu/cache/n25 ;
  wire \biu/cache/n27 ;
  wire \biu/cache/n29 ;
  wire \biu/cache/n3 ;
  wire \biu/cache/n31 ;
  wire \biu/cache/n5 ;
  wire \biu/cache/n7 ;
  wire \biu/cache/n9 ;
  wire \biu/cache_addr_sel ;  // ../../RTL/CPU/BIU/biu.v(79)
  wire \biu/cache_ctrl_logic/ex_l1d_chkok ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(158)
  wire \biu/cache_ctrl_logic/ex_l1d_hit ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(154)
  wire \biu/cache_ctrl_logic/ex_l1i_chkok ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(157)
  wire \biu/cache_ctrl_logic/ex_l1i_hit ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(155)
  wire \biu/cache_ctrl_logic/if_l1i_chkok ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(159)
  wire \biu/cache_ctrl_logic/if_l1i_hit ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(156)
  wire \biu/cache_ctrl_logic/l1d_miss ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(162)
  wire \biu/cache_ctrl_logic/l1d_value ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(138)
  wire \biu/cache_ctrl_logic/l1d_wr_sel ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(435)
  wire \biu/cache_ctrl_logic/l1d_write_burst ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(170)
  wire \biu/cache_ctrl_logic/l1d_write_through ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(178)
  wire \biu/cache_ctrl_logic/l1i_miss ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(161)
  wire \biu/cache_ctrl_logic/l1i_value ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(137)
  wire \biu/cache_ctrl_logic/l1i_wr_sel ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(434)
  wire \biu/cache_ctrl_logic/l1i_wr_sel_neg ;
  wire \biu/cache_ctrl_logic/l1i_write_burst ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(169)
  wire \biu/cache_ctrl_logic/l1i_write_through ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(177)
  wire \biu/cache_ctrl_logic/mux11_b2_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux20_b0_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux21_b0_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux22_b0_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux23_b0_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux24_b0_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux26_b2_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux2_b1_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux30_b4_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux31_b4_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux35_b3_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux36_b3_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux37_b4_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux39_b0_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux40_b2_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux41_b1_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux41_b2_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux42_b4_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux43_b1_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux43_b4_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux44_b4_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux6_b2_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux7_b1_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/mux7_b2_sel_is_2_o ;
  wire \biu/cache_ctrl_logic/mux9_b2_sel_is_0_o ;
  wire \biu/cache_ctrl_logic/n0 ;
  wire \biu/cache_ctrl_logic/n1 ;
  wire \biu/cache_ctrl_logic/n10 ;
  wire \biu/cache_ctrl_logic/n101 ;
  wire \biu/cache_ctrl_logic/n102 ;
  wire \biu/cache_ctrl_logic/n102_neg ;
  wire \biu/cache_ctrl_logic/n104 ;
  wire \biu/cache_ctrl_logic/n104_neg ;
  wire \biu/cache_ctrl_logic/n106 ;
  wire \biu/cache_ctrl_logic/n106_neg ;
  wire \biu/cache_ctrl_logic/n107 ;
  wire \biu/cache_ctrl_logic/n107_neg ;
  wire \biu/cache_ctrl_logic/n108 ;
  wire \biu/cache_ctrl_logic/n108_neg ;
  wire \biu/cache_ctrl_logic/n11 ;
  wire \biu/cache_ctrl_logic/n12 ;
  wire \biu/cache_ctrl_logic/n13 ;
  wire \biu/cache_ctrl_logic/n135 ;
  wire \biu/cache_ctrl_logic/n138 ;
  wire \biu/cache_ctrl_logic/n139 ;
  wire \biu/cache_ctrl_logic/n14 ;
  wire \biu/cache_ctrl_logic/n140 ;
  wire \biu/cache_ctrl_logic/n146 ;
  wire \biu/cache_ctrl_logic/n149 ;
  wire \biu/cache_ctrl_logic/n15 ;
  wire \biu/cache_ctrl_logic/n157 ;
  wire \biu/cache_ctrl_logic/n16 ;
  wire \biu/cache_ctrl_logic/n160 ;
  wire \biu/cache_ctrl_logic/n161 ;
  wire \biu/cache_ctrl_logic/n161_neg ;
  wire \biu/cache_ctrl_logic/n162 ;
  wire \biu/cache_ctrl_logic/n163 ;
  wire \biu/cache_ctrl_logic/n17 ;
  wire \biu/cache_ctrl_logic/n170 ;
  wire \biu/cache_ctrl_logic/n171 ;
  wire \biu/cache_ctrl_logic/n172 ;
  wire \biu/cache_ctrl_logic/n173 ;
  wire \biu/cache_ctrl_logic/n174 ;
  wire \biu/cache_ctrl_logic/n175 ;
  wire \biu/cache_ctrl_logic/n176 ;
  wire \biu/cache_ctrl_logic/n177 ;
  wire \biu/cache_ctrl_logic/n178 ;
  wire \biu/cache_ctrl_logic/n179 ;
  wire \biu/cache_ctrl_logic/n18 ;
  wire \biu/cache_ctrl_logic/n183 ;
  wire \biu/cache_ctrl_logic/n187 ;
  wire \biu/cache_ctrl_logic/n188 ;
  wire \biu/cache_ctrl_logic/n19 ;
  wire \biu/cache_ctrl_logic/n191 ;
  wire \biu/cache_ctrl_logic/n194 ;
  wire \biu/cache_ctrl_logic/n195 ;
  wire \biu/cache_ctrl_logic/n196 ;
  wire \biu/cache_ctrl_logic/n197 ;
  wire \biu/cache_ctrl_logic/n198 ;
  wire \biu/cache_ctrl_logic/n199 ;
  wire \biu/cache_ctrl_logic/n2 ;
  wire \biu/cache_ctrl_logic/n20 ;
  wire \biu/cache_ctrl_logic/n200 ;
  wire \biu/cache_ctrl_logic/n201 ;
  wire \biu/cache_ctrl_logic/n202 ;
  wire \biu/cache_ctrl_logic/n203 ;
  wire \biu/cache_ctrl_logic/n204 ;
  wire \biu/cache_ctrl_logic/n205 ;
  wire \biu/cache_ctrl_logic/n206 ;
  wire \biu/cache_ctrl_logic/n21 ;
  wire \biu/cache_ctrl_logic/n22 ;
  wire \biu/cache_ctrl_logic/n224 ;
  wire \biu/cache_ctrl_logic/n225 ;
  wire \biu/cache_ctrl_logic/n226 ;
  wire \biu/cache_ctrl_logic/n227 ;
  wire \biu/cache_ctrl_logic/n23 ;
  wire \biu/cache_ctrl_logic/n234 ;
  wire \biu/cache_ctrl_logic/n235 ;
  wire \biu/cache_ctrl_logic/n236 ;
  wire \biu/cache_ctrl_logic/n237 ;
  wire \biu/cache_ctrl_logic/n238 ;
  wire \biu/cache_ctrl_logic/n239 ;
  wire \biu/cache_ctrl_logic/n24 ;
  wire \biu/cache_ctrl_logic/n240 ;
  wire \biu/cache_ctrl_logic/n241 ;
  wire \biu/cache_ctrl_logic/n242 ;
  wire \biu/cache_ctrl_logic/n243 ;
  wire \biu/cache_ctrl_logic/n244 ;
  wire \biu/cache_ctrl_logic/n245 ;
  wire \biu/cache_ctrl_logic/n246 ;
  wire \biu/cache_ctrl_logic/n247 ;
  wire \biu/cache_ctrl_logic/n248 ;
  wire \biu/cache_ctrl_logic/n249 ;
  wire \biu/cache_ctrl_logic/n25 ;
  wire \biu/cache_ctrl_logic/n250 ;
  wire \biu/cache_ctrl_logic/n251 ;
  wire \biu/cache_ctrl_logic/n252 ;
  wire \biu/cache_ctrl_logic/n253 ;
  wire \biu/cache_ctrl_logic/n26 ;
  wire \biu/cache_ctrl_logic/n27 ;
  wire \biu/cache_ctrl_logic/n28 ;
  wire \biu/cache_ctrl_logic/n29 ;
  wire \biu/cache_ctrl_logic/n3 ;
  wire \biu/cache_ctrl_logic/n30 ;
  wire \biu/cache_ctrl_logic/n31 ;
  wire \biu/cache_ctrl_logic/n32 ;
  wire \biu/cache_ctrl_logic/n33 ;
  wire \biu/cache_ctrl_logic/n34 ;
  wire \biu/cache_ctrl_logic/n35 ;
  wire \biu/cache_ctrl_logic/n36 ;
  wire \biu/cache_ctrl_logic/n37 ;
  wire \biu/cache_ctrl_logic/n38 ;
  wire \biu/cache_ctrl_logic/n39 ;
  wire \biu/cache_ctrl_logic/n4 ;
  wire \biu/cache_ctrl_logic/n40 ;
  wire \biu/cache_ctrl_logic/n41 ;
  wire \biu/cache_ctrl_logic/n42 ;
  wire \biu/cache_ctrl_logic/n43 ;
  wire \biu/cache_ctrl_logic/n44 ;
  wire \biu/cache_ctrl_logic/n45 ;
  wire \biu/cache_ctrl_logic/n46 ;
  wire \biu/cache_ctrl_logic/n47 ;
  wire \biu/cache_ctrl_logic/n48 ;
  wire \biu/cache_ctrl_logic/n49 ;
  wire \biu/cache_ctrl_logic/n5 ;
  wire \biu/cache_ctrl_logic/n50 ;
  wire \biu/cache_ctrl_logic/n51 ;
  wire \biu/cache_ctrl_logic/n52 ;
  wire \biu/cache_ctrl_logic/n53 ;
  wire \biu/cache_ctrl_logic/n54 ;
  wire \biu/cache_ctrl_logic/n55 ;
  wire \biu/cache_ctrl_logic/n56 ;
  wire \biu/cache_ctrl_logic/n56_neg ;
  wire \biu/cache_ctrl_logic/n57 ;
  wire \biu/cache_ctrl_logic/n57_neg ;
  wire \biu/cache_ctrl_logic/n58 ;
  wire \biu/cache_ctrl_logic/n59 ;
  wire \biu/cache_ctrl_logic/n6 ;
  wire \biu/cache_ctrl_logic/n62 ;
  wire \biu/cache_ctrl_logic/n62_neg ;
  wire \biu/cache_ctrl_logic/n63 ;
  wire \biu/cache_ctrl_logic/n63_neg ;
  wire \biu/cache_ctrl_logic/n64 ;
  wire \biu/cache_ctrl_logic/n64_neg ;
  wire \biu/cache_ctrl_logic/n65 ;
  wire \biu/cache_ctrl_logic/n65_neg ;
  wire \biu/cache_ctrl_logic/n66 ;
  wire \biu/cache_ctrl_logic/n66_neg ;
  wire \biu/cache_ctrl_logic/n67 ;
  wire \biu/cache_ctrl_logic/n67_neg ;
  wire \biu/cache_ctrl_logic/n68 ;
  wire \biu/cache_ctrl_logic/n68_neg ;
  wire \biu/cache_ctrl_logic/n69 ;
  wire \biu/cache_ctrl_logic/n7 ;
  wire \biu/cache_ctrl_logic/n75 ;
  wire \biu/cache_ctrl_logic/n76 ;
  wire \biu/cache_ctrl_logic/n76_neg ;
  wire \biu/cache_ctrl_logic/n77 ;
  wire \biu/cache_ctrl_logic/n77_neg ;
  wire \biu/cache_ctrl_logic/n78 ;
  wire \biu/cache_ctrl_logic/n79 ;
  wire \biu/cache_ctrl_logic/n8 ;
  wire \biu/cache_ctrl_logic/n85 ;
  wire \biu/cache_ctrl_logic/n85_neg ;
  wire \biu/cache_ctrl_logic/n86 ;
  wire \biu/cache_ctrl_logic/n86_neg ;
  wire \biu/cache_ctrl_logic/n89 ;
  wire \biu/cache_ctrl_logic/n89_neg ;
  wire \biu/cache_ctrl_logic/n9 ;
  wire \biu/cache_ctrl_logic/n93 ;
  wire \biu/cache_ctrl_logic/n93_neg ;
  wire \biu/cache_ctrl_logic/n94 ;
  wire \biu/cache_ctrl_logic/n97 ;
  wire \biu/cache_ctrl_logic/n98 ;
  wire \biu/cache_ctrl_logic/pte_l1d_upd ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(174)
  wire \biu/cache_ctrl_logic/pte_l1i_upd ;  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(173)
  wire \biu/cache_ctrl_logic/u128_sel_is_0_o ;
  wire \biu/cache_write ;  // ../../RTL/CPU/BIU/biu.v(115)
  wire \biu/cacheable ;  // ../../RTL/CPU/BIU/biu.v(113)
  wire \biu/ex_data_sel[1]_neg ;
  wire \biu/l1d_write ;  // ../../RTL/CPU/BIU/biu.v(82)
  wire \biu/l1i_write ;  // ../../RTL/CPU/BIU/biu.v(83)
  wire \biu/new_pte_update ;  // ../../RTL/CPU/BIU/biu.v(107)
  wire \biu/opc[1]_neg ;
  wire \biu/pa_cov ;  // ../../RTL/CPU/BIU/biu.v(102)
  wire \biu/pa_cov_neg ;
  wire \biu/paddr ;  // ../../RTL/CPU/BIU/biu.v(99)
  wire \biu/page_fault ;  // ../../RTL/CPU/BIU/biu.v(116)
  wire \biu/page_fault_neg ;
  wire \biu/rd ;  // ../../RTL/CPU/BIU/biu.v(101)
  wire \biu/trans_rdy ;  // ../../RTL/CPU/BIU/biu.v(114)
  wire \biu/wr ;  // ../../RTL/CPU/BIU/biu.v(100)
  wire \biu/wr_neg ;
  wire cache_flush;  // ../../RTL/CPU/prv464_top.v(139)
  wire cache_flush_biu;  // ../../RTL/CPU/prv464_top.v(79)
  wire cache_ready_ex;  // ../../RTL/CPU/prv464_top.v(87)
  wire cache_ready_if;  // ../../RTL/CPU/prv464_top.v(70)
  wire cache_reset;  // ../../RTL/CPU/prv464_top.v(140)
  wire \cu_ru/add0_2_co ;
  wire \cu_ru/csr_satp/n0 ;
  wire \cu_ru/exc_target_m ;  // ../../RTL/CPU/CU&RU/cu_ru.v(146)
  wire \cu_ru/exc_target_s ;  // ../../RTL/CPU/CU&RU/cu_ru.v(145)
  wire \cu_ru/exception ;  // ../../RTL/CPU/CU&RU/cu_ru.v(140)
  wire \cu_ru/exception_neg ;
  wire \cu_ru/int_target_m ;  // ../../RTL/CPU/CU&RU/cu_ru.v(144)
  wire \cu_ru/int_target_s ;  // ../../RTL/CPU/CU&RU/cu_ru.v(143)
  wire \cu_ru/m_cycle_event/mcountinhibit[2] ;  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(16)
  wire \cu_ru/m_cycle_event/mcountinhibit[2]_neg ;
  wire \cu_ru/m_cycle_event/mux2_b0_sel_is_2_o ;
  wire \cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ;
  wire \cu_ru/m_cycle_event/n0 ;
  wire \cu_ru/m_cycle_event/n0_neg ;
  wire \cu_ru/m_cycle_event/n13 ;
  wire \cu_ru/m_s_cause/mux2_b0_sel_is_2_o ;
  wire \cu_ru/m_s_cause/mux4_b0_sel_is_2_o ;
  wire \cu_ru/m_s_cause/mux7_b10_sel_is_0_o ;
  wire \cu_ru/m_s_cause/n0 ;
  wire \cu_ru/m_s_cause/n0_neg ;
  wire \cu_ru/m_s_cause/n1 ;
  wire \cu_ru/m_s_epc/mux1_b0_sel_is_3_o ;
  wire \cu_ru/m_s_epc/mux4_b0_sel_is_2_o ;
  wire \cu_ru/m_s_epc/mux6_b0_sel_is_2_o ;
  wire \cu_ru/m_s_epc/n3 ;
  wire \cu_ru/m_s_epc/n3_neg ;
  wire \cu_ru/m_s_epc/n4 ;
  wire \cu_ru/m_s_ie/n0 ;
  wire \cu_ru/m_s_ie/n0_neg ;
  wire \cu_ru/m_s_ie/n1 ;
  wire \cu_ru/m_s_ie/n1_neg ;
  wire \cu_ru/m_s_ie/u11_sel_is_0_o ;
  wire \cu_ru/m_s_ip/n0 ;
  wire \cu_ru/m_s_ip/n0_neg ;
  wire \cu_ru/m_s_ip/n1 ;
  wire \cu_ru/m_s_ip/n2 ;
  wire \cu_ru/m_s_ip/n2_neg ;
  wire \cu_ru/m_s_ip/seip ;  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(28)
  wire \cu_ru/m_s_ip/u11_sel_is_0_o ;
  wire \cu_ru/m_s_ip/u12_sel_is_2_o ;
  wire \cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ;
  wire \cu_ru/m_s_scratch/n0 ;
  wire \cu_ru/m_s_scratch/n0_neg ;
  wire \cu_ru/m_s_scratch/n1 ;
  wire \cu_ru/m_s_status/mux1_b0_sel_is_0_o ;
  wire \cu_ru/m_s_status/mux3_b0_sel_is_2_o ;
  wire \cu_ru/m_s_status/n0 ;
  wire \cu_ru/m_s_status/n0_neg ;
  wire \cu_ru/m_s_status/n1 ;
  wire \cu_ru/m_s_status/n13 ;
  wire \cu_ru/m_s_status/n14 ;
  wire \cu_ru/m_s_status/n15 ;
  wire \cu_ru/m_s_status/n16 ;
  wire \cu_ru/m_s_status/n17 ;
  wire \cu_ru/m_s_status/n18 ;
  wire \cu_ru/m_s_status/n19 ;
  wire \cu_ru/m_s_status/n1_neg ;
  wire \cu_ru/m_s_status/n2 ;
  wire \cu_ru/m_s_status/n20 ;
  wire \cu_ru/m_s_status/n22 ;
  wire \cu_ru/m_s_status/n23 ;
  wire \cu_ru/m_s_status/n25 ;
  wire \cu_ru/m_s_status/n26 ;
  wire \cu_ru/m_s_status/n27 ;
  wire \cu_ru/m_s_status/n3 ;
  wire \cu_ru/m_s_status/n33 ;
  wire \cu_ru/m_s_status/n34 ;
  wire \cu_ru/m_s_status/n36 ;
  wire \cu_ru/m_s_status/n37 ;
  wire \cu_ru/m_s_status/n3_neg ;
  wire \cu_ru/m_s_status/n44 ;
  wire \cu_ru/m_s_status/n45 ;
  wire \cu_ru/m_s_status/n46 ;
  wire \cu_ru/m_s_status/u14_sel_is_2_o ;
  wire \cu_ru/m_s_status/u34_sel_is_0_o ;
  wire \cu_ru/m_s_tval/mux3_b0_sel_is_2_o ;
  wire \cu_ru/m_s_tval/mux5_b0_sel_is_2_o ;
  wire \cu_ru/m_s_tval/n0 ;
  wire \cu_ru/m_s_tval/n1 ;
  wire \cu_ru/m_s_tval/n2 ;
  wire \cu_ru/m_s_tval/n4 ;
  wire \cu_ru/m_s_tval/n4_neg ;
  wire \cu_ru/m_s_tval/n5 ;
  wire \cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ;
  wire \cu_ru/m_s_tvec/n0 ;
  wire \cu_ru/m_s_tvec/n0_neg ;
  wire \cu_ru/m_s_tvec/n1 ;
  wire \cu_ru/mcountinhibit ;  // ../../RTL/CPU/CU&RU/cu_ru.v(639)
  wire \cu_ru/medeleg_exc_ctrl/bk_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(73)
  wire \cu_ru/medeleg_exc_ctrl/bk_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(87)
  wire \cu_ru/medeleg_exc_ctrl/ecs_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(79)
  wire \cu_ru/medeleg_exc_ctrl/ecs_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(93)
  wire \cu_ru/medeleg_exc_ctrl/ecu_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(78)
  wire \cu_ru/medeleg_exc_ctrl/ecu_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(92)
  wire \cu_ru/medeleg_exc_ctrl/iaf_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(71)
  wire \cu_ru/medeleg_exc_ctrl/iaf_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(85)
  wire \cu_ru/medeleg_exc_ctrl/iam_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(70)
  wire \cu_ru/medeleg_exc_ctrl/iam_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(84)
  wire \cu_ru/medeleg_exc_ctrl/ii_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(72)
  wire \cu_ru/medeleg_exc_ctrl/ii_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(86)
  wire \cu_ru/medeleg_exc_ctrl/ipf_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(80)
  wire \cu_ru/medeleg_exc_ctrl/ipf_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(94)
  wire \cu_ru/medeleg_exc_ctrl/laf_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(75)
  wire \cu_ru/medeleg_exc_ctrl/laf_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(89)
  wire \cu_ru/medeleg_exc_ctrl/lam_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(74)
  wire \cu_ru/medeleg_exc_ctrl/lam_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(88)
  wire \cu_ru/medeleg_exc_ctrl/lpf_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(81)
  wire \cu_ru/medeleg_exc_ctrl/lpf_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(95)
  wire \cu_ru/medeleg_exc_ctrl/mux10_b1_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux10_b1_sel_is_2_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux10_b3_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux10_b3_sel_is_0_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux11_b1_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux11_b3_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux1_b0_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux1_b1_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux1_b1_sel_is_2_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux2_b0_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux2_b1_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux2_b1_sel_is_0_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux2_b3_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux2_b3_sel_is_0_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux3_b1_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux3_b1_sel_is_0_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux3_b3_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux4_b0_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux4_b1_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux4_b1_sel_is_0_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux4_b3_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux4_b3_sel_is_2_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux5_b0_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux5_b1_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux5_b3_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux6_b1_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux6_b2_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux6_b3_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux6_b3_sel_is_2_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux7_b1_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux7_b1_sel_is_2_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux7_b2_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux7_b3_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux8_b1_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux8_b1_sel_is_0_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/mux8_b2_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux8_b3_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux9_b1_sel_is_0_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux9_b2_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux9_b3_sel_is_2_o ;
  wire \cu_ru/medeleg_exc_ctrl/mux9_b3_sel_is_2_o_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n0 ;
  wire \cu_ru/medeleg_exc_ctrl/n100 ;
  wire \cu_ru/medeleg_exc_ctrl/n101 ;
  wire \cu_ru/medeleg_exc_ctrl/n102 ;
  wire \cu_ru/medeleg_exc_ctrl/n103 ;
  wire \cu_ru/medeleg_exc_ctrl/n104 ;
  wire \cu_ru/medeleg_exc_ctrl/n105 ;
  wire \cu_ru/medeleg_exc_ctrl/n106 ;
  wire \cu_ru/medeleg_exc_ctrl/n107 ;
  wire \cu_ru/medeleg_exc_ctrl/n108 ;
  wire \cu_ru/medeleg_exc_ctrl/n109 ;
  wire \cu_ru/medeleg_exc_ctrl/n110 ;
  wire \cu_ru/medeleg_exc_ctrl/n111 ;
  wire \cu_ru/medeleg_exc_ctrl/n112 ;
  wire \cu_ru/medeleg_exc_ctrl/n113 ;
  wire \cu_ru/medeleg_exc_ctrl/n114 ;
  wire \cu_ru/medeleg_exc_ctrl/n115 ;
  wire \cu_ru/medeleg_exc_ctrl/n116 ;
  wire \cu_ru/medeleg_exc_ctrl/n117 ;
  wire \cu_ru/medeleg_exc_ctrl/n118 ;
  wire \cu_ru/medeleg_exc_ctrl/n119 ;
  wire \cu_ru/medeleg_exc_ctrl/n120 ;
  wire \cu_ru/medeleg_exc_ctrl/n121 ;
  wire \cu_ru/medeleg_exc_ctrl/n122 ;
  wire \cu_ru/medeleg_exc_ctrl/n123 ;
  wire \cu_ru/medeleg_exc_ctrl/n27 ;
  wire \cu_ru/medeleg_exc_ctrl/n28 ;
  wire \cu_ru/medeleg_exc_ctrl/n29 ;
  wire \cu_ru/medeleg_exc_ctrl/n30 ;
  wire \cu_ru/medeleg_exc_ctrl/n31 ;
  wire \cu_ru/medeleg_exc_ctrl/n32 ;
  wire \cu_ru/medeleg_exc_ctrl/n33 ;
  wire \cu_ru/medeleg_exc_ctrl/n34 ;
  wire \cu_ru/medeleg_exc_ctrl/n35 ;
  wire \cu_ru/medeleg_exc_ctrl/n36 ;
  wire \cu_ru/medeleg_exc_ctrl/n37 ;
  wire \cu_ru/medeleg_exc_ctrl/n38 ;
  wire \cu_ru/medeleg_exc_ctrl/n39 ;
  wire \cu_ru/medeleg_exc_ctrl/n40 ;
  wire \cu_ru/medeleg_exc_ctrl/n41 ;
  wire \cu_ru/medeleg_exc_ctrl/n42 ;
  wire \cu_ru/medeleg_exc_ctrl/n43 ;
  wire \cu_ru/medeleg_exc_ctrl/n44 ;
  wire \cu_ru/medeleg_exc_ctrl/n45 ;
  wire \cu_ru/medeleg_exc_ctrl/n46 ;
  wire \cu_ru/medeleg_exc_ctrl/n47 ;
  wire \cu_ru/medeleg_exc_ctrl/n48 ;
  wire \cu_ru/medeleg_exc_ctrl/n49 ;
  wire \cu_ru/medeleg_exc_ctrl/n50 ;
  wire \cu_ru/medeleg_exc_ctrl/n51 ;
  wire \cu_ru/medeleg_exc_ctrl/n52 ;
  wire \cu_ru/medeleg_exc_ctrl/n53 ;
  wire \cu_ru/medeleg_exc_ctrl/n54 ;
  wire \cu_ru/medeleg_exc_ctrl/n55 ;
  wire \cu_ru/medeleg_exc_ctrl/n56 ;
  wire \cu_ru/medeleg_exc_ctrl/n57 ;
  wire \cu_ru/medeleg_exc_ctrl/n58 ;
  wire \cu_ru/medeleg_exc_ctrl/n59 ;
  wire \cu_ru/medeleg_exc_ctrl/n60 ;
  wire \cu_ru/medeleg_exc_ctrl/n61 ;
  wire \cu_ru/medeleg_exc_ctrl/n62 ;
  wire \cu_ru/medeleg_exc_ctrl/n63 ;
  wire \cu_ru/medeleg_exc_ctrl/n64 ;
  wire \cu_ru/medeleg_exc_ctrl/n65 ;
  wire \cu_ru/medeleg_exc_ctrl/n66 ;
  wire \cu_ru/medeleg_exc_ctrl/n67 ;
  wire \cu_ru/medeleg_exc_ctrl/n68 ;
  wire \cu_ru/medeleg_exc_ctrl/n69 ;
  wire \cu_ru/medeleg_exc_ctrl/n70 ;
  wire \cu_ru/medeleg_exc_ctrl/n71 ;
  wire \cu_ru/medeleg_exc_ctrl/n72 ;
  wire \cu_ru/medeleg_exc_ctrl/n73 ;
  wire \cu_ru/medeleg_exc_ctrl/n74 ;
  wire \cu_ru/medeleg_exc_ctrl/n75 ;
  wire \cu_ru/medeleg_exc_ctrl/n76 ;
  wire \cu_ru/medeleg_exc_ctrl/n76_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n77 ;
  wire \cu_ru/medeleg_exc_ctrl/n77_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n78 ;
  wire \cu_ru/medeleg_exc_ctrl/n78_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n79 ;
  wire \cu_ru/medeleg_exc_ctrl/n79_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n80 ;
  wire \cu_ru/medeleg_exc_ctrl/n80_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n81 ;
  wire \cu_ru/medeleg_exc_ctrl/n81_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n82 ;
  wire \cu_ru/medeleg_exc_ctrl/n82_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n83 ;
  wire \cu_ru/medeleg_exc_ctrl/n83_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n84 ;
  wire \cu_ru/medeleg_exc_ctrl/n84_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n85 ;
  wire \cu_ru/medeleg_exc_ctrl/n85_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n86 ;
  wire \cu_ru/medeleg_exc_ctrl/n86_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n87 ;
  wire \cu_ru/medeleg_exc_ctrl/n87_neg ;
  wire \cu_ru/medeleg_exc_ctrl/n88 ;
  wire \cu_ru/medeleg_exc_ctrl/saf_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(77)
  wire \cu_ru/medeleg_exc_ctrl/saf_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(91)
  wire \cu_ru/medeleg_exc_ctrl/sam_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(76)
  wire \cu_ru/medeleg_exc_ctrl/sam_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(90)
  wire \cu_ru/medeleg_exc_ctrl/spf_target_m ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(82)
  wire \cu_ru/medeleg_exc_ctrl/spf_target_s ;  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(96)
  wire \cu_ru/mideleg_int_ctrl/mei_ack_m ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(58)
  wire \cu_ru/mideleg_int_ctrl/mei_ack_m_neg ;
  wire \cu_ru/mideleg_int_ctrl/msi_ack_m ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(59)
  wire \cu_ru/mideleg_int_ctrl/msi_ack_m_neg ;
  wire \cu_ru/mideleg_int_ctrl/mti_ack_m ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(60)
  wire \cu_ru/mideleg_int_ctrl/mti_ack_m_neg ;
  wire \cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o ;
  wire \cu_ru/mideleg_int_ctrl/mux2_b0_sel_is_2_o ;
  wire \cu_ru/mideleg_int_ctrl/mux2_b3_sel_is_2_o ;
  wire \cu_ru/mideleg_int_ctrl/mux3_b0_sel_is_2_o ;
  wire \cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o ;
  wire \cu_ru/mideleg_int_ctrl/mux3_b3_sel_is_2_o ;
  wire \cu_ru/mideleg_int_ctrl/mux3_b3_sel_is_2_o_neg ;
  wire \cu_ru/mideleg_int_ctrl/mux4_b0_sel_is_2_o ;
  wire \cu_ru/mideleg_int_ctrl/mux4_b1_sel_is_2_o ;
  wire \cu_ru/mideleg_int_ctrl/mux4_b2_sel_is_0_o ;
  wire \cu_ru/mideleg_int_ctrl/mux4_b3_sel_is_0_o ;
  wire \cu_ru/mideleg_int_ctrl/n0 ;
  wire \cu_ru/mideleg_int_ctrl/n10 ;
  wire \cu_ru/mideleg_int_ctrl/n11 ;
  wire \cu_ru/mideleg_int_ctrl/n12 ;
  wire \cu_ru/mideleg_int_ctrl/n13 ;
  wire \cu_ru/mideleg_int_ctrl/n14 ;
  wire \cu_ru/mideleg_int_ctrl/n15 ;
  wire \cu_ru/mideleg_int_ctrl/n16 ;
  wire \cu_ru/mideleg_int_ctrl/n18 ;
  wire \cu_ru/mideleg_int_ctrl/n19 ;
  wire \cu_ru/mideleg_int_ctrl/n20 ;
  wire \cu_ru/mideleg_int_ctrl/n21 ;
  wire \cu_ru/mideleg_int_ctrl/n22 ;
  wire \cu_ru/mideleg_int_ctrl/n23 ;
  wire \cu_ru/mideleg_int_ctrl/n24 ;
  wire \cu_ru/mideleg_int_ctrl/n25 ;
  wire \cu_ru/mideleg_int_ctrl/n26 ;
  wire \cu_ru/mideleg_int_ctrl/n27 ;
  wire \cu_ru/mideleg_int_ctrl/n28 ;
  wire \cu_ru/mideleg_int_ctrl/n29 ;
  wire \cu_ru/mideleg_int_ctrl/n30 ;
  wire \cu_ru/mideleg_int_ctrl/n31 ;
  wire \cu_ru/mideleg_int_ctrl/n32 ;
  wire \cu_ru/mideleg_int_ctrl/n33 ;
  wire \cu_ru/mideleg_int_ctrl/n33_neg ;
  wire \cu_ru/mideleg_int_ctrl/n34 ;
  wire \cu_ru/mideleg_int_ctrl/n34_neg ;
  wire \cu_ru/mideleg_int_ctrl/n35 ;
  wire \cu_ru/mideleg_int_ctrl/n7 ;
  wire \cu_ru/mideleg_int_ctrl/n8 ;
  wire \cu_ru/mideleg_int_ctrl/n9 ;
  wire \cu_ru/mideleg_int_ctrl/sei_ack_m ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(61)
  wire \cu_ru/mideleg_int_ctrl/sei_ack_s ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(65)
  wire \cu_ru/mideleg_int_ctrl/ssi_ack_m ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(62)
  wire \cu_ru/mideleg_int_ctrl/ssi_ack_s ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(66)
  wire \cu_ru/mideleg_int_ctrl/sti_ack_m ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(63)
  wire \cu_ru/mideleg_int_ctrl/sti_ack_s ;  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(67)
  wire \cu_ru/mie ;  // ../../RTL/CPU/CU&RU/cu_ru.v(381)
  wire \cu_ru/mrw_mcause_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(207)
  wire \cu_ru/mrw_mcounterinhibit_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(217)
  wire \cu_ru/mrw_mcycle_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(213)
  wire \cu_ru/mrw_medeleg_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(200)
  wire \cu_ru/mrw_mepc_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(206)
  wire \cu_ru/mrw_mideleg_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(201)
  wire \cu_ru/mrw_mie_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(202)
  wire \cu_ru/mrw_mip_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(209)
  wire \cu_ru/mrw_mscratch_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(205)
  wire \cu_ru/mrw_mstatus_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(198)
  wire \cu_ru/mrw_mtval_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(208)
  wire \cu_ru/mrw_mtvec_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(203)
  wire \cu_ru/mux34_b0_sel_is_2_o ;
  wire \cu_ru/n0 ;
  wire \cu_ru/n1 ;
  wire \cu_ru/n10 ;
  wire \cu_ru/n11 ;
  wire \cu_ru/n116 ;
  wire \cu_ru/n12 ;
  wire \cu_ru/n13 ;
  wire \cu_ru/n14 ;
  wire \cu_ru/n15 ;
  wire \cu_ru/n16 ;
  wire \cu_ru/n17 ;
  wire \cu_ru/n18 ;
  wire \cu_ru/n19 ;
  wire \cu_ru/n2 ;
  wire \cu_ru/n20 ;
  wire \cu_ru/n23 ;
  wire \cu_ru/n24 ;
  wire \cu_ru/n25 ;
  wire \cu_ru/n26 ;
  wire \cu_ru/n27 ;
  wire \cu_ru/n28 ;
  wire \cu_ru/n29 ;
  wire \cu_ru/n3 ;
  wire \cu_ru/n30 ;
  wire \cu_ru/n31 ;
  wire \cu_ru/n33 ;
  wire \cu_ru/n34 ;
  wire \cu_ru/n35 ;
  wire \cu_ru/n36 ;
  wire \cu_ru/n37 ;
  wire \cu_ru/n38 ;
  wire \cu_ru/n39 ;
  wire \cu_ru/n4 ;
  wire \cu_ru/n40 ;
  wire \cu_ru/n41 ;
  wire \cu_ru/n42 ;
  wire \cu_ru/n45 ;
  wire \cu_ru/n48 ;
  wire \cu_ru/n5 ;
  wire \cu_ru/n51 ;
  wire \cu_ru/n53 ;
  wire \cu_ru/n56 ;
  wire \cu_ru/n6 ;
  wire \cu_ru/n66 ;
  wire \cu_ru/n7 ;
  wire \cu_ru/n8 ;
  wire \cu_ru/n9 ;
  wire \cu_ru/n98 ;
  wire \cu_ru/next_pc ;  // ../../RTL/CPU/CU&RU/cu_ru.v(150)
  wire \cu_ru/read_cycle_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(220)
  wire \cu_ru/read_instret_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(222)
  wire \cu_ru/read_marchid_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(236)
  wire \cu_ru/read_mcause_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(248)
  wire \cu_ru/read_mcounterinhibit_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(258)
  wire \cu_ru/read_mcycle_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(254)
  wire \cu_ru/read_medeleg_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(241)
  wire \cu_ru/read_mepc_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(247)
  wire \cu_ru/read_mideleg_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(242)
  wire \cu_ru/read_mie_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(243)
  wire \cu_ru/read_mimp_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(237)
  wire \cu_ru/read_minstret_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(255)
  wire \cu_ru/read_mip_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(250)
  wire \cu_ru/read_mscratch_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(246)
  wire \cu_ru/read_mstatus_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(239)
  wire \cu_ru/read_mtval_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(249)
  wire \cu_ru/read_mtvec_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(244)
  wire \cu_ru/read_mvendorid_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(235)
  wire \cu_ru/read_satp_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(234)
  wire \cu_ru/read_scause_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(231)
  wire \cu_ru/read_sepc_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(230)
  wire \cu_ru/read_sie_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(226)
  wire \cu_ru/read_sip_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(233)
  wire \cu_ru/read_sscratch_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(229)
  wire \cu_ru/read_sstatus_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(225)
  wire \cu_ru/read_stval_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(232)
  wire \cu_ru/read_stvec_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(227)
  wire \cu_ru/read_time_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(221)
  wire \cu_ru/srw_satp_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(193)
  wire \cu_ru/srw_scause_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(190)
  wire \cu_ru/srw_sepc_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(189)
  wire \cu_ru/srw_sie_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(185)
  wire \cu_ru/srw_sip_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(192)
  wire \cu_ru/srw_sscratch_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(188)
  wire \cu_ru/srw_sstatus_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(184)
  wire \cu_ru/srw_stval_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(191)
  wire \cu_ru/srw_stvec_sel ;  // ../../RTL/CPU/CU&RU/cu_ru.v(186)
  wire \cu_ru/trap_target_m ;  // ../../RTL/CPU/CU&RU/cu_ru.v(148)
  wire \cu_ru/trap_target_m_neg ;
  wire \cu_ru/trap_target_s ;  // ../../RTL/CPU/CU&RU/cu_ru.v(149)
  wire \cu_ru/trap_target_s_neg ;
  wire ex_csr_write;  // ../../RTL/CPU/prv464_top.v(145)
  wire ex_ebreak;  // ../../RTL/CPU/prv464_top.v(171)
  wire ex_ecall;  // ../../RTL/CPU/prv464_top.v(170)
  wire ex_gpr_write;  // ../../RTL/CPU/prv464_top.v(146)
  wire ex_ill_ins;  // ../../RTL/CPU/prv464_top.v(167)
  wire ex_ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(162)
  wire ex_ins_addr_mis;  // ../../RTL/CPU/prv464_top.v(163)
  wire ex_ins_page_fault;  // ../../RTL/CPU/prv464_top.v(164)
  wire ex_int_acc;  // ../../RTL/CPU/prv464_top.v(165)
  wire ex_jmp;  // ../../RTL/CPU/prv464_top.v(161)
  wire ex_m_ret;  // ../../RTL/CPU/prv464_top.v(168)
  wire ex_more_exception;  // ../../RTL/CPU/prv464_top.v(576)
  wire ex_more_exception_neg;
  wire ex_nop;  // ../../RTL/CPU/prv464_top.v(580)
  wire ex_ready;  // ../../RTL/CPU/prv464_top.v(577)
  wire ex_s_ret;  // ../../RTL/CPU/prv464_top.v(169)
  wire \ex_size[2]_neg ;
  wire ex_system;  // ../../RTL/CPU/prv464_top.v(160)
  wire ex_valid;  // ../../RTL/CPU/prv464_top.v(166)
  wire \exu/alu_au/ds1_great_than_ds2 ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(68)
  wire \exu/alu_au/ds1_light_than_ds2 ;  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(67)
  wire \exu/alu_au/n0 ;
  wire \exu/alu_au/n10 ;
  wire \exu/alu_au/n11 ;
  wire \exu/alu_au/n12 ;
  wire \exu/alu_au/n13 ;
  wire \exu/alu_au/n14 ;
  wire \exu/alu_au/n15 ;
  wire \exu/alu_au/n2 ;
  wire \exu/alu_au/n4 ;
  wire \exu/alu_au/n5 ;
  wire \exu/alu_au/n6 ;
  wire \exu/alu_au/n7 ;
  wire \exu/alu_au/n8 ;
  wire \exu/alu_au/n9 ;
  wire \exu/amo_ready ;  // ../../RTL/CPU/EX/exu.v(208)
  wire \exu/c_amo_mem0 ;  // ../../RTL/CPU/EX/exu.v(178)
  wire \exu/c_amo_mem01 ;  // ../../RTL/CPU/EX/exu.v(179)
  wire \exu/c_amo_mem01_neg ;
  wire \exu/c_amo_mem0_neg ;
  wire \exu/c_amo_mem1 ;  // ../../RTL/CPU/EX/exu.v(181)
  wire \exu/c_amo_mem1_neg ;
  wire \exu/c_fence ;  // ../../RTL/CPU/EX/exu.v(182)
  wire \exu/c_load ;  // ../../RTL/CPU/EX/exu.v(175)
  wire \exu/c_load_1 ;  // ../../RTL/CPU/EX/exu.v(176)
  wire \exu/c_load_neg ;
  wire \exu/c_shift ;  // ../../RTL/CPU/EX/exu.v(174)
  wire \exu/c_shift_neg ;
  wire \exu/c_stb ;  // ../../RTL/CPU/EX/exu.v(173)
  wire \exu/c_store ;  // ../../RTL/CPU/EX/exu.v(177)
  wire \exu/c_store_neg ;
  wire \exu/exception_id ;  // ../../RTL/CPU/EX/exu.v(199)
  wire \exu/fence_ready ;  // ../../RTL/CPU/EX/exu.v(207)
  wire \exu/load_addr_mis ;  // ../../RTL/CPU/EX/exu.v(202)
  wire \exu/load_ready ;  // ../../RTL/CPU/EX/exu.v(205)
  wire \exu/lsu/mux27_b56_sel_is_3_o ;
  wire \exu/lsu/n0 ;
  wire \exu/lsu/n2 ;
  wire \exu/lsu/n5 ;
  wire \exu/lsu/n51 ;
  wire \exu/lsu/n53 ;
  wire \exu/lsu/n56 ;
  wire \exu/lsu/n8 ;
  wire \exu/mux12_b2_sel_is_0_o ;
  wire \exu/mux13_b1_sel_is_0_o ;
  wire \exu/mux13_b2_sel_is_2_o ;
  wire \exu/mux16_b2_sel_is_0_o ;
  wire \exu/mux17_b1_sel_is_0_o ;
  wire \exu/mux18_b3_sel_is_2_o ;
  wire \exu/mux1_b0_sel_is_0_o ;
  wire \exu/mux27_b32_sel_is_1_o ;
  wire \exu/mux27_b63_sel_is_3_o ;
  wire \exu/mux2_b1_sel_is_2_o ;
  wire \exu/mux2_b2_sel_is_0_o ;
  wire \exu/mux3_b1_sel_is_2_o ;
  wire \exu/mux3_b3_sel_is_0_o ;
  wire \exu/mux48_b32_sel_is_1_o ;
  wire \exu/mux4_b0_sel_is_0_o ;
  wire \exu/mux4_b3_sel_is_2_o ;
  wire \exu/mux8_b1_sel_is_2_o ;
  wire \exu/n0 ;
  wire \exu/n10 ;
  wire \exu/n11 ;
  wire \exu/n12 ;
  wire \exu/n13 ;
  wire \exu/n132 ;
  wire \exu/n133 ;
  wire \exu/n134 ;
  wire \exu/n135 ;
  wire \exu/n136 ;
  wire \exu/n137 ;
  wire \exu/n138 ;
  wire \exu/n139 ;
  wire \exu/n14 ;
  wire \exu/n140 ;
  wire \exu/n141 ;
  wire \exu/n142 ;
  wire \exu/n143 ;
  wire \exu/n144 ;
  wire \exu/n145 ;
  wire \exu/n146 ;
  wire \exu/n147 ;
  wire \exu/n148 ;
  wire \exu/n149 ;
  wire \exu/n15 ;
  wire \exu/n16 ;
  wire \exu/n17 ;
  wire \exu/n18 ;
  wire \exu/n19 ;
  wire \exu/n2 ;
  wire \exu/n20 ;
  wire \exu/n20_neg ;
  wire \exu/n21 ;
  wire \exu/n21_neg ;
  wire \exu/n28 ;
  wire \exu/n3 ;
  wire \exu/n31 ;
  wire \exu/n35 ;
  wire \exu/n35_neg ;
  wire \exu/n4 ;
  wire \exu/n48 ;
  wire \exu/n49 ;
  wire \exu/n5 ;
  wire \exu/n59 ;
  wire \exu/n6 ;
  wire \exu/n60 ;
  wire \exu/n7 ;
  wire \exu/n8 ;
  wire \exu/n86 ;
  wire \exu/n87 ;
  wire \exu/n88 ;
  wire \exu/n89 ;
  wire \exu/n9 ;
  wire \exu/n90 ;
  wire \exu/n91 ;
  wire \exu/n92 ;
  wire \exu/n93 ;
  wire \exu/n94 ;
  wire \exu/n95 ;
  wire \exu/shift_multi_ready ;  // ../../RTL/CPU/EX/exu.v(209)
  wire \exu/shift_ready ;  // ../../RTL/CPU/EX/exu.v(188)
  wire \exu/store_addr_mis ;  // ../../RTL/CPU/EX/exu.v(203)
  wire \exu/store_ready ;  // ../../RTL/CPU/EX/exu.v(206)
  wire id_branch;  // ../../RTL/CPU/prv464_top.v(174)
  wire id_hold;  // ../../RTL/CPU/prv464_top.v(177)
  wire id_hold_neg;
  wire id_ill_ins;  // ../../RTL/CPU/prv464_top.v(176)
  wire id_ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(92)
  wire id_ins_addr_mis;  // ../../RTL/CPU/prv464_top.v(93)
  wire id_ins_page_fault;  // ../../RTL/CPU/prv464_top.v(94)
  wire id_int_acc;  // ../../RTL/CPU/prv464_top.v(95)
  wire id_nop;  // ../../RTL/CPU/prv464_top.v(178)
  wire id_nop_neg;
  wire id_system;  // ../../RTL/CPU/prv464_top.v(175)
  wire id_valid;  // ../../RTL/CPU/prv464_top.v(96)
  wire if_hold;  // ../../RTL/CPU/prv464_top.v(263)
  wire if_nop;  // ../../RTL/CPU/prv464_top.v(262)
  wire ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(68)
  wire ins_acc_fault_neg;
  wire \ins_dec/dbyte ;  // ../../RTL/CPU/ID/ins_dec.v(235)
  wire \ins_dec/dec_csr_acc_fault ;  // ../../RTL/CPU/ID/ins_dec.v(334)
  wire \ins_dec/dec_gpr_write ;  // ../../RTL/CPU/ID/ins_dec.v(119)
  wire \ins_dec/dec_ins_dec_fault ;  // ../../RTL/CPU/ID/ins_dec.v(336)
  wire \ins_dec/dec_ins_unpermit ;  // ../../RTL/CPU/ID/ins_dec.v(335)
  wire \ins_dec/ds1_mem_iden ;  // ../../RTL/CPU/ID/ins_dec.v(339)
  wire \ins_dec/funct12_0 ;  // ../../RTL/CPU/ID/ins_dec.v(223)
  wire \ins_dec/funct12_1 ;  // ../../RTL/CPU/ID/ins_dec.v(224)
  wire \ins_dec/funct3_0 ;  // ../../RTL/CPU/ID/ins_dec.v(172)
  wire \ins_dec/funct3_1 ;  // ../../RTL/CPU/ID/ins_dec.v(173)
  wire \ins_dec/funct3_2 ;  // ../../RTL/CPU/ID/ins_dec.v(174)
  wire \ins_dec/funct3_3 ;  // ../../RTL/CPU/ID/ins_dec.v(175)
  wire \ins_dec/funct3_4 ;  // ../../RTL/CPU/ID/ins_dec.v(176)
  wire \ins_dec/funct3_5 ;  // ../../RTL/CPU/ID/ins_dec.v(177)
  wire \ins_dec/funct3_6 ;  // ../../RTL/CPU/ID/ins_dec.v(178)
  wire \ins_dec/funct3_7 ;  // ../../RTL/CPU/ID/ins_dec.v(179)
  wire \ins_dec/funct5_0 ;  // ../../RTL/CPU/ID/ins_dec.v(181)
  wire \ins_dec/funct5_1 ;  // ../../RTL/CPU/ID/ins_dec.v(182)
  wire \ins_dec/funct5_12 ;  // ../../RTL/CPU/ID/ins_dec.v(193)
  wire \ins_dec/funct5_16 ;  // ../../RTL/CPU/ID/ins_dec.v(197)
  wire \ins_dec/funct5_2 ;  // ../../RTL/CPU/ID/ins_dec.v(183)
  wire \ins_dec/funct5_20 ;  // ../../RTL/CPU/ID/ins_dec.v(201)
  wire \ins_dec/funct5_24 ;  // ../../RTL/CPU/ID/ins_dec.v(205)
  wire \ins_dec/funct5_28 ;  // ../../RTL/CPU/ID/ins_dec.v(209)
  wire \ins_dec/funct5_3 ;  // ../../RTL/CPU/ID/ins_dec.v(184)
  wire \ins_dec/funct5_4 ;  // ../../RTL/CPU/ID/ins_dec.v(185)
  wire \ins_dec/funct5_8 ;  // ../../RTL/CPU/ID/ins_dec.v(189)
  wire \ins_dec/funct6_0 ;  // ../../RTL/CPU/ID/ins_dec.v(214)
  wire \ins_dec/funct6_16 ;  // ../../RTL/CPU/ID/ins_dec.v(215)
  wire \ins_dec/funct7_0 ;  // ../../RTL/CPU/ID/ins_dec.v(220)
  wire \ins_dec/funct7_24 ;  // ../../RTL/CPU/ID/ins_dec.v(218)
  wire \ins_dec/funct7_32 ;  // ../../RTL/CPU/ID/ins_dec.v(217)
  wire \ins_dec/funct7_8 ;  // ../../RTL/CPU/ID/ins_dec.v(219)
  wire \ins_dec/funct7_9 ;  // ../../RTL/CPU/ID/ins_dec.v(410)
  wire \ins_dec/ins_add ;  // ../../RTL/CPU/ID/ins_dec.v(272)
  wire \ins_dec/ins_addi ;  // ../../RTL/CPU/ID/ins_dec.v(262)
  wire \ins_dec/ins_addiw ;  // ../../RTL/CPU/ID/ins_dec.v(295)
  wire \ins_dec/ins_addw ;  // ../../RTL/CPU/ID/ins_dec.v(299)
  wire \ins_dec/ins_amoaddd ;  // ../../RTL/CPU/ID/ins_dec.v(320)
  wire \ins_dec/ins_amoaddw ;  // ../../RTL/CPU/ID/ins_dec.v(308)
  wire \ins_dec/ins_amoandd ;  // ../../RTL/CPU/ID/ins_dec.v(322)
  wire \ins_dec/ins_amoandw ;  // ../../RTL/CPU/ID/ins_dec.v(310)
  wire \ins_dec/ins_amomaxd ;  // ../../RTL/CPU/ID/ins_dec.v(325)
  wire \ins_dec/ins_amomaxud ;  // ../../RTL/CPU/ID/ins_dec.v(327)
  wire \ins_dec/ins_amomaxuw ;  // ../../RTL/CPU/ID/ins_dec.v(315)
  wire \ins_dec/ins_amomaxw ;  // ../../RTL/CPU/ID/ins_dec.v(313)
  wire \ins_dec/ins_amomind ;  // ../../RTL/CPU/ID/ins_dec.v(324)
  wire \ins_dec/ins_amominud ;  // ../../RTL/CPU/ID/ins_dec.v(326)
  wire \ins_dec/ins_amominuw ;  // ../../RTL/CPU/ID/ins_dec.v(314)
  wire \ins_dec/ins_amominw ;  // ../../RTL/CPU/ID/ins_dec.v(312)
  wire \ins_dec/ins_amoord ;  // ../../RTL/CPU/ID/ins_dec.v(323)
  wire \ins_dec/ins_amoorw ;  // ../../RTL/CPU/ID/ins_dec.v(311)
  wire \ins_dec/ins_amoswapd ;  // ../../RTL/CPU/ID/ins_dec.v(319)
  wire \ins_dec/ins_amoswapw ;  // ../../RTL/CPU/ID/ins_dec.v(307)
  wire \ins_dec/ins_amoxord ;  // ../../RTL/CPU/ID/ins_dec.v(321)
  wire \ins_dec/ins_amoxorw ;  // ../../RTL/CPU/ID/ins_dec.v(309)
  wire \ins_dec/ins_and ;  // ../../RTL/CPU/ID/ins_dec.v(281)
  wire \ins_dec/ins_andi ;  // ../../RTL/CPU/ID/ins_dec.v(268)
  wire \ins_dec/ins_bgeu ;  // ../../RTL/CPU/ID/ins_dec.v(251)
  wire \ins_dec/ins_bltu ;  // ../../RTL/CPU/ID/ins_dec.v(250)
  wire \ins_dec/ins_csrrc ;  // ../../RTL/CPU/ID/ins_dec.v(287)
  wire \ins_dec/ins_csrrci ;  // ../../RTL/CPU/ID/ins_dec.v(290)
  wire \ins_dec/ins_csrrs ;  // ../../RTL/CPU/ID/ins_dec.v(286)
  wire \ins_dec/ins_csrrsi ;  // ../../RTL/CPU/ID/ins_dec.v(289)
  wire \ins_dec/ins_csrrw ;  // ../../RTL/CPU/ID/ins_dec.v(285)
  wire \ins_dec/ins_csrrwi ;  // ../../RTL/CPU/ID/ins_dec.v(288)
  wire \ins_dec/ins_ebreak ;  // ../../RTL/CPU/ID/ins_dec.v(284)
  wire \ins_dec/ins_ecall ;  // ../../RTL/CPU/ID/ins_dec.v(283)
  wire \ins_dec/ins_fence ;  // ../../RTL/CPU/ID/ins_dec.v(282)
  wire \ins_dec/ins_lb ;  // ../../RTL/CPU/ID/ins_dec.v(252)
  wire \ins_dec/ins_lbu ;  // ../../RTL/CPU/ID/ins_dec.v(253)
  wire \ins_dec/ins_ld ;  // ../../RTL/CPU/ID/ins_dec.v(293)
  wire \ins_dec/ins_lh ;  // ../../RTL/CPU/ID/ins_dec.v(254)
  wire \ins_dec/ins_lhu ;  // ../../RTL/CPU/ID/ins_dec.v(255)
  wire \ins_dec/ins_lrd ;  // ../../RTL/CPU/ID/ins_dec.v(317)
  wire \ins_dec/ins_lrw ;  // ../../RTL/CPU/ID/ins_dec.v(305)
  wire \ins_dec/ins_lw ;  // ../../RTL/CPU/ID/ins_dec.v(256)
  wire \ins_dec/ins_lwu ;  // ../../RTL/CPU/ID/ins_dec.v(292)
  wire \ins_dec/ins_mret ;  // ../../RTL/CPU/ID/ins_dec.v(329)
  wire \ins_dec/ins_or ;  // ../../RTL/CPU/ID/ins_dec.v(280)
  wire \ins_dec/ins_ori ;  // ../../RTL/CPU/ID/ins_dec.v(267)
  wire \ins_dec/ins_sb ;  // ../../RTL/CPU/ID/ins_dec.v(258)
  wire \ins_dec/ins_scd ;  // ../../RTL/CPU/ID/ins_dec.v(318)
  wire \ins_dec/ins_scw ;  // ../../RTL/CPU/ID/ins_dec.v(306)
  wire \ins_dec/ins_sfencevma ;  // ../../RTL/CPU/ID/ins_dec.v(331)
  wire \ins_dec/ins_sh ;  // ../../RTL/CPU/ID/ins_dec.v(259)
  wire \ins_dec/ins_sll ;  // ../../RTL/CPU/ID/ins_dec.v(274)
  wire \ins_dec/ins_slli ;  // ../../RTL/CPU/ID/ins_dec.v(269)
  wire \ins_dec/ins_slliw ;  // ../../RTL/CPU/ID/ins_dec.v(296)
  wire \ins_dec/ins_sllw ;  // ../../RTL/CPU/ID/ins_dec.v(301)
  wire \ins_dec/ins_slt ;  // ../../RTL/CPU/ID/ins_dec.v(275)
  wire \ins_dec/ins_slti ;  // ../../RTL/CPU/ID/ins_dec.v(264)
  wire \ins_dec/ins_sltiu ;  // ../../RTL/CPU/ID/ins_dec.v(265)
  wire \ins_dec/ins_sltu ;  // ../../RTL/CPU/ID/ins_dec.v(276)
  wire \ins_dec/ins_sra ;  // ../../RTL/CPU/ID/ins_dec.v(279)
  wire \ins_dec/ins_srai ;  // ../../RTL/CPU/ID/ins_dec.v(271)
  wire \ins_dec/ins_sraiw ;  // ../../RTL/CPU/ID/ins_dec.v(298)
  wire \ins_dec/ins_sraw ;  // ../../RTL/CPU/ID/ins_dec.v(303)
  wire \ins_dec/ins_sret ;  // ../../RTL/CPU/ID/ins_dec.v(330)
  wire \ins_dec/ins_srl ;  // ../../RTL/CPU/ID/ins_dec.v(278)
  wire \ins_dec/ins_srli ;  // ../../RTL/CPU/ID/ins_dec.v(270)
  wire \ins_dec/ins_srliw ;  // ../../RTL/CPU/ID/ins_dec.v(297)
  wire \ins_dec/ins_srlw ;  // ../../RTL/CPU/ID/ins_dec.v(302)
  wire \ins_dec/ins_sub ;  // ../../RTL/CPU/ID/ins_dec.v(273)
  wire \ins_dec/ins_subw ;  // ../../RTL/CPU/ID/ins_dec.v(300)
  wire \ins_dec/ins_sw ;  // ../../RTL/CPU/ID/ins_dec.v(260)
  wire \ins_dec/ins_wfi ;  // ../../RTL/CPU/ID/ins_dec.v(505)
  wire \ins_dec/ins_xor ;  // ../../RTL/CPU/ID/ins_dec.v(277)
  wire \ins_dec/ins_xori ;  // ../../RTL/CPU/ID/ins_dec.v(266)
  wire \ins_dec/mux13_b0_sel_is_0_o ;
  wire \ins_dec/mux19_b10_sel_is_2_o ;
  wire \ins_dec/mux1_b6_sel_is_0_o ;
  wire \ins_dec/mux20_b56_sel_is_0_o ;
  wire \ins_dec/mux24_b10_sel_is_0_o ;
  wire \ins_dec/mux25_b56_sel_is_0_o ;
  wire \ins_dec/mux25_b56_sel_is_0_o_neg ;
  wire \ins_dec/mux26_b20_sel_is_0_o ;
  wire \ins_dec/mux26_b56_sel_is_0_o ;
  wire \ins_dec/mux26_b56_sel_is_0_o_neg ;
  wire \ins_dec/mux27_b12_sel_is_0_o ;
  wire \ins_dec/mux27_b20_sel_is_2_o ;
  wire \ins_dec/mux27_b56_sel_is_0_o ;
  wire \ins_dec/n0 ;
  wire \ins_dec/n1 ;
  wire \ins_dec/n10 ;
  wire \ins_dec/n100 ;
  wire \ins_dec/n101 ;
  wire \ins_dec/n102 ;
  wire \ins_dec/n103 ;
  wire \ins_dec/n104 ;
  wire \ins_dec/n105 ;
  wire \ins_dec/n106 ;
  wire \ins_dec/n107 ;
  wire \ins_dec/n107_neg ;
  wire \ins_dec/n108 ;
  wire \ins_dec/n109 ;
  wire \ins_dec/n11 ;
  wire \ins_dec/n110 ;
  wire \ins_dec/n111 ;
  wire \ins_dec/n112 ;
  wire \ins_dec/n113 ;
  wire \ins_dec/n114 ;
  wire \ins_dec/n115 ;
  wire \ins_dec/n116 ;
  wire \ins_dec/n117 ;
  wire \ins_dec/n118 ;
  wire \ins_dec/n119 ;
  wire \ins_dec/n12 ;
  wire \ins_dec/n120 ;
  wire \ins_dec/n121 ;
  wire \ins_dec/n122 ;
  wire \ins_dec/n123 ;
  wire \ins_dec/n124 ;
  wire \ins_dec/n125 ;
  wire \ins_dec/n126 ;
  wire \ins_dec/n127 ;
  wire \ins_dec/n128 ;
  wire \ins_dec/n129 ;
  wire \ins_dec/n13 ;
  wire \ins_dec/n130 ;
  wire \ins_dec/n131 ;
  wire \ins_dec/n132 ;
  wire \ins_dec/n133 ;
  wire \ins_dec/n134 ;
  wire \ins_dec/n135 ;
  wire \ins_dec/n136 ;
  wire \ins_dec/n137 ;
  wire \ins_dec/n138 ;
  wire \ins_dec/n139 ;
  wire \ins_dec/n14 ;
  wire \ins_dec/n141 ;
  wire \ins_dec/n142 ;
  wire \ins_dec/n143 ;
  wire \ins_dec/n144 ;
  wire \ins_dec/n145 ;
  wire \ins_dec/n146 ;
  wire \ins_dec/n147 ;
  wire \ins_dec/n148 ;
  wire \ins_dec/n149 ;
  wire \ins_dec/n15 ;
  wire \ins_dec/n150 ;
  wire \ins_dec/n151 ;
  wire \ins_dec/n152 ;
  wire \ins_dec/n153 ;
  wire \ins_dec/n154 ;
  wire \ins_dec/n155 ;
  wire \ins_dec/n156 ;
  wire \ins_dec/n157 ;
  wire \ins_dec/n158 ;
  wire \ins_dec/n16 ;
  wire \ins_dec/n17 ;
  wire \ins_dec/n18 ;
  wire \ins_dec/n19 ;
  wire \ins_dec/n195 ;
  wire \ins_dec/n196 ;
  wire \ins_dec/n197 ;
  wire \ins_dec/n198 ;
  wire \ins_dec/n199 ;
  wire \ins_dec/n2 ;
  wire \ins_dec/n20 ;
  wire \ins_dec/n200 ;
  wire \ins_dec/n201 ;
  wire \ins_dec/n202 ;
  wire \ins_dec/n203 ;
  wire \ins_dec/n204 ;
  wire \ins_dec/n205 ;
  wire \ins_dec/n206 ;
  wire \ins_dec/n21 ;
  wire \ins_dec/n22 ;
  wire \ins_dec/n225 ;
  wire \ins_dec/n226 ;
  wire \ins_dec/n227 ;
  wire \ins_dec/n228 ;
  wire \ins_dec/n229 ;
  wire \ins_dec/n23 ;
  wire \ins_dec/n230 ;
  wire \ins_dec/n231 ;
  wire \ins_dec/n232 ;
  wire \ins_dec/n233 ;
  wire \ins_dec/n234 ;
  wire \ins_dec/n235 ;
  wire \ins_dec/n236 ;
  wire \ins_dec/n237 ;
  wire \ins_dec/n238 ;
  wire \ins_dec/n239 ;
  wire \ins_dec/n24 ;
  wire \ins_dec/n25 ;
  wire \ins_dec/n26 ;
  wire \ins_dec/n266 ;
  wire \ins_dec/n267 ;
  wire \ins_dec/n268 ;
  wire \ins_dec/n269 ;
  wire \ins_dec/n27 ;
  wire \ins_dec/n273 ;
  wire \ins_dec/n274 ;
  wire \ins_dec/n275 ;
  wire \ins_dec/n275_neg ;
  wire \ins_dec/n276 ;
  wire \ins_dec/n277 ;
  wire \ins_dec/n277_neg ;
  wire \ins_dec/n278 ;
  wire \ins_dec/n279 ;
  wire \ins_dec/n28 ;
  wire \ins_dec/n285 ;
  wire \ins_dec/n29 ;
  wire \ins_dec/n3 ;
  wire \ins_dec/n30 ;
  wire \ins_dec/n302 ;
  wire \ins_dec/n303 ;
  wire \ins_dec/n304 ;
  wire \ins_dec/n305 ;
  wire \ins_dec/n31 ;
  wire \ins_dec/n32 ;
  wire \ins_dec/n33 ;
  wire \ins_dec/n34 ;
  wire \ins_dec/n35 ;
  wire \ins_dec/n36 ;
  wire \ins_dec/n37 ;
  wire \ins_dec/n38 ;
  wire \ins_dec/n39 ;
  wire \ins_dec/n4 ;
  wire \ins_dec/n40 ;
  wire \ins_dec/n41 ;
  wire \ins_dec/n42 ;
  wire \ins_dec/n43 ;
  wire \ins_dec/n44 ;
  wire \ins_dec/n45 ;
  wire \ins_dec/n46 ;
  wire \ins_dec/n47 ;
  wire \ins_dec/n48 ;
  wire \ins_dec/n49 ;
  wire \ins_dec/n5 ;
  wire \ins_dec/n50 ;
  wire \ins_dec/n51 ;
  wire \ins_dec/n52 ;
  wire \ins_dec/n53 ;
  wire \ins_dec/n54 ;
  wire \ins_dec/n55 ;
  wire \ins_dec/n55_neg ;
  wire \ins_dec/n56 ;
  wire \ins_dec/n57 ;
  wire \ins_dec/n57_neg ;
  wire \ins_dec/n59 ;
  wire \ins_dec/n6 ;
  wire \ins_dec/n60 ;
  wire \ins_dec/n61 ;
  wire \ins_dec/n62 ;
  wire \ins_dec/n63 ;
  wire \ins_dec/n64 ;
  wire \ins_dec/n65 ;
  wire \ins_dec/n66 ;
  wire \ins_dec/n67 ;
  wire \ins_dec/n68 ;
  wire \ins_dec/n69 ;
  wire \ins_dec/n7 ;
  wire \ins_dec/n70 ;
  wire \ins_dec/n71 ;
  wire \ins_dec/n72 ;
  wire \ins_dec/n73 ;
  wire \ins_dec/n74 ;
  wire \ins_dec/n75 ;
  wire \ins_dec/n78 ;
  wire \ins_dec/n8 ;
  wire \ins_dec/n80 ;
  wire \ins_dec/n81 ;
  wire \ins_dec/n82 ;
  wire \ins_dec/n83 ;
  wire \ins_dec/n84 ;
  wire \ins_dec/n86 ;
  wire \ins_dec/n87 ;
  wire \ins_dec/n88 ;
  wire \ins_dec/n89 ;
  wire \ins_dec/n9 ;
  wire \ins_dec/n90 ;
  wire \ins_dec/n91 ;
  wire \ins_dec/n92 ;
  wire \ins_dec/n93 ;
  wire \ins_dec/n94 ;
  wire \ins_dec/n95 ;
  wire \ins_dec/n96 ;
  wire \ins_dec/n97 ;
  wire \ins_dec/n98 ;
  wire \ins_dec/n99 ;
  wire \ins_dec/obyte ;  // ../../RTL/CPU/ID/ins_dec.v(237)
  wire \ins_dec/op_32_imm ;  // ../../RTL/CPU/ID/ins_dec.v(158)
  wire \ins_dec/op_32_reg ;  // ../../RTL/CPU/ID/ins_dec.v(167)
  wire \ins_dec/op_amo ;  // ../../RTL/CPU/ID/ins_dec.v(168)
  wire \ins_dec/op_auipc ;  // ../../RTL/CPU/ID/ins_dec.v(160)
  wire \ins_dec/op_branch ;  // ../../RTL/CPU/ID/ins_dec.v(163)
  wire \ins_dec/op_branch_neg ;
  wire \ins_dec/op_imm ;  // ../../RTL/CPU/ID/ins_dec.v(157)
  wire \ins_dec/op_jal ;  // ../../RTL/CPU/ID/ins_dec.v(161)
  wire \ins_dec/op_jal_neg ;
  wire \ins_dec/op_jalr ;  // ../../RTL/CPU/ID/ins_dec.v(162)
  wire \ins_dec/op_jalr_neg ;
  wire \ins_dec/op_load ;  // ../../RTL/CPU/ID/ins_dec.v(165)
  wire \ins_dec/op_load_neg ;
  wire \ins_dec/op_lui ;  // ../../RTL/CPU/ID/ins_dec.v(159)
  wire \ins_dec/op_reg ;  // ../../RTL/CPU/ID/ins_dec.v(166)
  wire \ins_dec/op_store ;  // ../../RTL/CPU/ID/ins_dec.v(164)
  wire \ins_dec/op_store_neg ;
  wire \ins_dec/qbyte ;  // ../../RTL/CPU/ID/ins_dec.v(236)
  wire \ins_dec/sbyte ;  // ../../RTL/CPU/ID/ins_dec.v(234)
  wire \ins_dec/u461_sel_is_0_o ;
  wire \ins_dec/u478_sel_is_0_o ;
  wire \ins_fetch/addr_mis ;  // ../../RTL/CPU/IF/ins_fetch.v(57)
  wire \ins_fetch/hold ;  // ../../RTL/CPU/IF/ins_fetch.v(53)
  wire \ins_fetch/hold_neg ;
  wire \ins_fetch/mux8_b0_sel_is_2_o ;
  wire \ins_fetch/n0 ;
  wire \ins_fetch/n0_neg ;
  wire \ins_fetch/n23 ;
  wire \ins_fetch/n24 ;
  wire \ins_fetch/n25 ;
  wire \ins_fetch/n26 ;
  wire \ins_fetch/n27 ;
  wire \ins_fetch/n31 ;
  wire \ins_fetch/n9 ;
  wire \ins_fetch/u72_sel_is_1_o ;
  wire ins_page_fault;  // ../../RTL/CPU/prv464_top.v(69)
  wire int_req;  // ../../RTL/CPU/prv464_top.v(259)
  wire jmp;  // ../../RTL/CPU/prv464_top.v(127)
  wire load;  // ../../RTL/CPU/prv464_top.v(136)
  wire load_acc_fault;  // ../../RTL/CPU/prv464_top.v(83)
  wire load_acc_fault_neg;
  wire load_neg;
  wire load_page_fault;  // ../../RTL/CPU/prv464_top.v(84)
  wire mem_csr_data_add;  // ../../RTL/CPU/prv464_top.v(116)
  wire mem_csr_data_and;  // ../../RTL/CPU/prv464_top.v(117)
  wire mem_csr_data_ds2;  // ../../RTL/CPU/prv464_top.v(115)
  wire mem_csr_data_max;  // ../../RTL/CPU/prv464_top.v(120)
  wire mem_csr_data_min;  // ../../RTL/CPU/prv464_top.v(121)
  wire mem_csr_data_or;  // ../../RTL/CPU/prv464_top.v(118)
  wire mem_csr_data_xor;  // ../../RTL/CPU/prv464_top.v(119)
  wire mprv;  // ../../RTL/CPU/prv464_top.v(53)
  wire mxr;  // ../../RTL/CPU/prv464_top.v(52)
  wire pc_jmp;  // ../../RTL/CPU/prv464_top.v(522)
  wire \pip_ctrl/ex_exception ;  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(80)
  wire \pip_ctrl/id_ex_war ;  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(83)
  wire \pip_ctrl/id_exception ;  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(79)
  wire \pip_ctrl/id_wb_war ;  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(84)
  wire \pip_ctrl/n0 ;
  wire \pip_ctrl/n1 ;
  wire \pip_ctrl/n10 ;
  wire \pip_ctrl/n11 ;
  wire \pip_ctrl/n12 ;
  wire \pip_ctrl/n13 ;
  wire \pip_ctrl/n14 ;
  wire \pip_ctrl/n15 ;
  wire \pip_ctrl/n16 ;
  wire \pip_ctrl/n17 ;
  wire \pip_ctrl/n18 ;
  wire \pip_ctrl/n19 ;
  wire \pip_ctrl/n2 ;
  wire \pip_ctrl/n20 ;
  wire \pip_ctrl/n21 ;
  wire \pip_ctrl/n22 ;
  wire \pip_ctrl/n23 ;
  wire \pip_ctrl/n24 ;
  wire \pip_ctrl/n25 ;
  wire \pip_ctrl/n26 ;
  wire \pip_ctrl/n27 ;
  wire \pip_ctrl/n28 ;
  wire \pip_ctrl/n29 ;
  wire \pip_ctrl/n3 ;
  wire \pip_ctrl/n30 ;
  wire \pip_ctrl/n31 ;
  wire \pip_ctrl/n32 ;
  wire \pip_ctrl/n33 ;
  wire \pip_ctrl/n34 ;
  wire \pip_ctrl/n35 ;
  wire \pip_ctrl/n36 ;
  wire \pip_ctrl/n37 ;
  wire \pip_ctrl/n38 ;
  wire \pip_ctrl/n39 ;
  wire \pip_ctrl/n4 ;
  wire \pip_ctrl/n40 ;
  wire \pip_ctrl/n41 ;
  wire \pip_ctrl/n42 ;
  wire \pip_ctrl/n43 ;
  wire \pip_ctrl/n44 ;
  wire \pip_ctrl/n45 ;
  wire \pip_ctrl/n46 ;
  wire \pip_ctrl/n47 ;
  wire \pip_ctrl/n48 ;
  wire \pip_ctrl/n49 ;
  wire \pip_ctrl/n5 ;
  wire \pip_ctrl/n50 ;
  wire \pip_ctrl/n51 ;
  wire \pip_ctrl/n52 ;
  wire \pip_ctrl/n53 ;
  wire \pip_ctrl/n55 ;
  wire \pip_ctrl/n56 ;
  wire \pip_ctrl/n57 ;
  wire \pip_ctrl/n58 ;
  wire \pip_ctrl/n59 ;
  wire \pip_ctrl/n6 ;
  wire \pip_ctrl/n7 ;
  wire \pip_ctrl/n8 ;
  wire \pip_ctrl/n9 ;
  wire pip_flush;  // ../../RTL/CPU/prv464_top.v(265)
  wire \priv[1]_neg ;
  wire \priv[3]_neg ;
  wire rd_data_add;  // ../../RTL/CPU/prv464_top.v(104)
  wire rd_data_and;  // ../../RTL/CPU/prv464_top.v(106)
  wire rd_data_ds1;  // ../../RTL/CPU/prv464_top.v(103)
  wire rd_data_or;  // ../../RTL/CPU/prv464_top.v(107)
  wire rd_data_slt;  // ../../RTL/CPU/prv464_top.v(109)
  wire rd_data_sub;  // ../../RTL/CPU/prv464_top.v(105)
  wire rd_data_xor;  // ../../RTL/CPU/prv464_top.v(108)
  wire rd_ins;  // ../../RTL/CPU/prv464_top.v(66)
  wire read;  // ../../RTL/CPU/prv464_top.v(81)
  wire rst_neg;
  wire shift_l;  // ../../RTL/CPU/prv464_top.v(142)
  wire shift_r;  // ../../RTL/CPU/prv464_top.v(141)
  wire store;  // ../../RTL/CPU/prv464_top.v(137)
  wire store_acc_fault;  // ../../RTL/CPU/prv464_top.v(85)
  wire store_acc_fault_neg;
  wire store_neg;
  wire store_page_fault;  // ../../RTL/CPU/prv464_top.v(86)
  wire sum;  // ../../RTL/CPU/prv464_top.v(51)
  wire tsr;  // ../../RTL/CPU/prv464_top.v(50)
  wire tvm;  // ../../RTL/CPU/prv464_top.v(49)
  wire tw;  // ../../RTL/CPU/prv464_top.v(309)
  wire uncache_data_rdy;  // ../../RTL/CPU/prv464_top.v(88)
  wire unpage;  // ../../RTL/CPU/prv464_top.v(72)
  wire unsign;  // ../../RTL/CPU/prv464_top.v(128)
  wire wb_csr_write;  // ../../RTL/CPU/prv464_top.v(520)
  wire wb_ebreak;  // ../../RTL/CPU/prv464_top.v(547)
  wire wb_ecall;  // ../../RTL/CPU/prv464_top.v(546)
  wire wb_gpr_write;  // ../../RTL/CPU/prv464_top.v(521)
  wire wb_ill_ins;  // ../../RTL/CPU/prv464_top.v(543)
  wire wb_ins_acc_fault;  // ../../RTL/CPU/prv464_top.v(532)
  wire wb_ins_addr_mis;  // ../../RTL/CPU/prv464_top.v(533)
  wire wb_ins_page_fault;  // ../../RTL/CPU/prv464_top.v(534)
  wire wb_int_acc;  // ../../RTL/CPU/prv464_top.v(541)
  wire wb_jmp;  // ../../RTL/CPU/prv464_top.v(531)
  wire wb_ld_acc_fault;  // ../../RTL/CPU/prv464_top.v(537)
  wire wb_ld_addr_mis;  // ../../RTL/CPU/prv464_top.v(535)
  wire wb_ld_page_fault;  // ../../RTL/CPU/prv464_top.v(539)
  wire wb_m_ret;  // ../../RTL/CPU/prv464_top.v(544)
  wire wb_s_ret;  // ../../RTL/CPU/prv464_top.v(545)
  wire wb_st_acc_fault;  // ../../RTL/CPU/prv464_top.v(538)
  wire wb_st_addr_mis;  // ../../RTL/CPU/prv464_top.v(536)
  wire wb_st_page_fault;  // ../../RTL/CPU/prv464_top.v(540)
  wire wb_system;  // ../../RTL/CPU/prv464_top.v(530)
  wire wb_valid;  // ../../RTL/CPU/prv464_top.v(542)
  wire write;  // ../../RTL/CPU/prv464_top.v(82)

  assign hburst[2] = 1'b0;
  assign hburst[1] = 1'b0;
  assign hmastlock = 1'b0;
  assign hprot[3] = 1'b0;
  assign hprot[2] = 1'b0;
  assign hprot[1] = 1'b1;
  assign hprot[0] = 1'b1;
  assign hsize[2] = 1'b0;
  not amo_inv (amo_neg, amo);
  not \biu/bus_error_inv  (\biu/bus_error_neg , \biu/bus_error );
  add_pu9_pu9_o9 \biu/bus_unit/add0  (
    .i0(\biu/bus_unit/addr_counter ),
    .i1(9'b000000001),
    .o(\biu/bus_unit/n39 ));  // ../../RTL/CPU/BIU/bus_unit.v(175)
  add_pu61_pu61_o61 \biu/bus_unit/add1  (
    .i0({52'b0000000000000000000000000000000000000000000000000000,\biu/bus_unit/addr_counter }),
    .i1(\biu/maddress [63:3]),
    .o(\biu/bus_unit/n49 ));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  eq_w5 \biu/bus_unit/eq0  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b00000),
    .o(\biu/bus_unit/n0 ));  // ../../RTL/CPU/BIU/bus_unit.v(126)
  eq_w5 \biu/bus_unit/eq1  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b00001),
    .o(\biu/bus_unit/n7 ));  // ../../RTL/CPU/BIU/bus_unit.v(130)
  eq_w5 \biu/bus_unit/eq10  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b11111),
    .o(\biu/bus_unit/n25 ));  // ../../RTL/CPU/BIU/bus_unit.v(160)
  eq_w5 \biu/bus_unit/eq11  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b01000),
    .o(\biu/bus_unit/n45 ));  // ../../RTL/CPU/BIU/bus_unit.v(181)
  eq_w5 \biu/bus_unit/eq2  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b01001),
    .o(\biu/bus_unit/n11 ));  // ../../RTL/CPU/BIU/bus_unit.v(134)
  eq_w5 \biu/bus_unit/eq3  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b00010),
    .o(\biu/bus_unit/n12 ));  // ../../RTL/CPU/BIU/bus_unit.v(137)
  eq_w5 \biu/bus_unit/eq4  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b00100),
    .o(\biu/bus_unit/n13 ));  // ../../RTL/CPU/BIU/bus_unit.v(140)
  eq_w5 \biu/bus_unit/eq5  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b01010),
    .o(\biu/bus_unit/n14 ));  // ../../RTL/CPU/BIU/bus_unit.v(145)
  eq_w9 \biu/bus_unit/eq6  (
    .i0(\biu/bus_unit/addr_counter ),
    .i1(9'b111111111),
    .o(\biu/bus_unit/n15 ));  // ../../RTL/CPU/BIU/bus_unit.v(146)
  eq_w5 \biu/bus_unit/eq7  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b00011),
    .o(\biu/bus_unit/n18 ));  // ../../RTL/CPU/BIU/bus_unit.v(148)
  eq_w5 \biu/bus_unit/eq8  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b00101),
    .o(\biu/bus_unit/n20 ));  // ../../RTL/CPU/BIU/bus_unit.v(151)
  eq_w5 \biu/bus_unit/eq9  (
    .i0(\biu/bus_unit/statu ),
    .i1(5'b01011),
    .o(\biu/bus_unit/n22 ));  // ../../RTL/CPU/BIU/bus_unit.v(156)
  eq_w2 \biu/bus_unit/mmu/eq0  (
    .i0(\biu/bus_unit/mmu/i ),
    .i1(2'b00),
    .o(\biu/bus_unit/mmu/n1 ));  // ../../RTL/CPU/BIU/mmu.v(105)
  eq_w3 \biu/bus_unit/mmu/eq1  (
    .i0({\biu/priv [3],\biu/priv [1:0]}),
    .i1(3'b001),
    .o(\biu/bus_unit/mmu/n7 ));  // ../../RTL/CPU/BIU/mmu.v(110)
  eq_w4 \biu/bus_unit/mmu/eq10  (
    .i0(satp[63:60]),
    .i1(4'b1000),
    .o(\biu/bus_unit/mmu/n31 ));  // ../../RTL/CPU/BIU/mmu.v(125)
  eq_w4 \biu/bus_unit/mmu/eq11  (
    .i0(\biu/bus_unit/mmu/statu ),
    .i1(4'b0001),
    .o(\biu/bus_unit/mmu/n34 ));  // ../../RTL/CPU/BIU/mmu.v(127)
  eq_w4 \biu/bus_unit/mmu/eq12  (
    .i0(\biu/bus_unit/mmu/statu ),
    .i1(4'b0010),
    .o(\biu/bus_unit/mmu/n35 ));  // ../../RTL/CPU/BIU/mmu.v(130)
  eq_w4 \biu/bus_unit/mmu/eq13  (
    .i0(\biu/bus_unit/mmu/statu ),
    .i1(4'b0011),
    .o(\biu/bus_unit/mmu/n37 ));  // ../../RTL/CPU/BIU/mmu.v(133)
  eq_w4 \biu/bus_unit/mmu/eq14  (
    .i0(\biu/bus_unit/mmu/statu ),
    .i1(4'b0100),
    .o(\biu/bus_unit/mmu/n41 ));  // ../../RTL/CPU/BIU/mmu.v(136)
  eq_w4 \biu/bus_unit/mmu/eq15  (
    .i0(\biu/bus_unit/mmu/statu ),
    .i1(4'b0101),
    .o(\biu/bus_unit/mmu_hwrite ));  // ../../RTL/CPU/BIU/mmu.v(139)
  eq_w4 \biu/bus_unit/mmu/eq16  (
    .i0(\biu/bus_unit/mmu/statu ),
    .i1(4'b0110),
    .o(\biu/bus_unit/mmu/n45 ));  // ../../RTL/CPU/BIU/mmu.v(142)
  eq_w4 \biu/bus_unit/mmu/eq17  (
    .i0(\biu/bus_unit/mmu/statu ),
    .i1(4'b0111),
    .o(\biu/bus_unit/mmu_trans_rdy ));  // ../../RTL/CPU/BIU/mmu.v(145)
  eq_w4 \biu/bus_unit/mmu/eq18  (
    .i0(\biu/bus_unit/mmu/statu ),
    .i1(4'b1000),
    .o(\biu/bus_unit/mmu_page_fault ));  // ../../RTL/CPU/BIU/mmu.v(148)
  eq_w4 \biu/bus_unit/mmu/eq19  (
    .i0(\biu/bus_unit/mmu/statu ),
    .i1(4'b1001),
    .o(\biu/bus_unit/mmu_acc_fault ));  // ../../RTL/CPU/BIU/mmu.v(151)
  eq_w3 \biu/bus_unit/mmu/eq2  (
    .i0({\biu/priv [3],\biu/priv [1:0]}),
    .i1(3'b010),
    .o(\biu/bus_unit/mmu/n8 ));  // ../../RTL/CPU/BIU/mmu.v(110)
  eq_w32 \biu/bus_unit/mmu/eq20  (
    .i0(\biu/paddress [63:32]),
    .i1(cacheability_block),
    .o(\biu/bus_unit/mmu/n81 ));  // ../../RTL/CPU/BIU/mmu.v(221)
  eq_w2 \biu/bus_unit/mmu/eq3  (
    .i0(\biu/opc ),
    .i1(2'b01),
    .o(\biu/bus_unit/mmu/n12 ));  // ../../RTL/CPU/BIU/mmu.v(111)
  eq_w2 \biu/bus_unit/mmu/eq4  (
    .i0(\biu/opc ),
    .i1(2'b00),
    .o(\biu/bus_unit/mmu/n14 ));  // ../../RTL/CPU/BIU/mmu.v(111)
  eq_w2 \biu/bus_unit/mmu/eq5  (
    .i0(\biu/opc ),
    .i1(2'b10),
    .o(\biu/bus_unit/mmu/n19 ));  // ../../RTL/CPU/BIU/mmu.v(111)
  eq_w3 \biu/bus_unit/mmu/eq6  (
    .i0({\biu/priv [3],\biu/priv [1:0]}),
    .i1(3'b100),
    .o(\biu/bus_unit/mmu/n25 ));  // ../../RTL/CPU/BIU/mmu.v(113)
  eq_w2 \biu/bus_unit/mmu/eq7  (
    .i0(\biu/bus_unit/mmu/i ),
    .i1(2'b10),
    .o(\biu/bus_unit/mmu/n26 ));  // ../../RTL/CPU/BIU/mmu.v(115)
  eq_w2 \biu/bus_unit/mmu/eq8  (
    .i0(\biu/bus_unit/mmu/i ),
    .i1(2'b01),
    .o(\biu/bus_unit/mmu/n27 ));  // ../../RTL/CPU/BIU/mmu.v(115)
  eq_w4 \biu/bus_unit/mmu/eq9  (
    .i0(\biu/bus_unit/mmu/statu ),
    .i1(4'b0000),
    .o(\biu/bus_unit/mmu/n30 ));  // ../../RTL/CPU/BIU/mmu.v(124)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux0_b0  (
    .i0(1'b0),
    .i1(\biu/maddress [30]),
    .sel(\biu/bus_unit/mmu/n1 ),
    .o(\biu/bus_unit/mmu/n28 [0]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux0_b1  (
    .i0(1'b0),
    .i1(\biu/maddress [31]),
    .sel(\biu/bus_unit/mmu/n1 ),
    .o(\biu/bus_unit/mmu/n28 [1]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux0_b2  (
    .i0(1'b0),
    .i1(\biu/maddress [32]),
    .sel(\biu/bus_unit/mmu/n1 ),
    .o(\biu/bus_unit/mmu/n28 [2]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux0_b3  (
    .i0(1'b0),
    .i1(\biu/maddress [33]),
    .sel(\biu/bus_unit/mmu/n1 ),
    .o(\biu/bus_unit/mmu/n28 [3]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux0_b4  (
    .i0(1'b0),
    .i1(\biu/maddress [34]),
    .sel(\biu/bus_unit/mmu/n1 ),
    .o(\biu/bus_unit/mmu/n28 [4]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux0_b5  (
    .i0(1'b0),
    .i1(\biu/maddress [35]),
    .sel(\biu/bus_unit/mmu/n1 ),
    .o(\biu/bus_unit/mmu/n28 [5]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux0_b6  (
    .i0(1'b0),
    .i1(\biu/maddress [36]),
    .sel(\biu/bus_unit/mmu/n1 ),
    .o(\biu/bus_unit/mmu/n28 [6]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux0_b7  (
    .i0(1'b0),
    .i1(\biu/maddress [37]),
    .sel(\biu/bus_unit/mmu/n1 ),
    .o(\biu/bus_unit/mmu/n28 [7]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux0_b8  (
    .i0(1'b0),
    .i1(\biu/maddress [38]),
    .sel(\biu/bus_unit/mmu/n1 ),
    .o(\biu/bus_unit/mmu/n28 [8]));  // ../../RTL/CPU/BIU/mmu.v(115)
  AL_MUX \biu/bus_unit/mmu/mux10_b0  (
    .i0(1'b0),
    .i1(\biu/bus_unit/mmu/statu [0]),
    .sel(\biu/bus_unit/mmu/mux10_b0_sel_is_2_o ),
    .o(\biu/bus_unit/mmu/n49 [0]));
  and \biu/bus_unit/mmu/mux10_b0_sel_is_2  (\biu/bus_unit/mmu/mux10_b0_sel_is_2_o , \biu/bus_unit/mmu_trans_rdy_neg , \biu/bus_unit/mmu/mux9_b0_sel_is_0_o );
  AL_MUX \biu/bus_unit/mmu/mux10_b1  (
    .i0(1'b0),
    .i1(\biu/bus_unit/mmu/statu [1]),
    .sel(\biu/bus_unit/mmu/mux10_b0_sel_is_2_o ),
    .o(\biu/bus_unit/mmu/n49 [1]));
  AL_MUX \biu/bus_unit/mmu/mux10_b2  (
    .i0(1'b0),
    .i1(\biu/bus_unit/mmu/statu [2]),
    .sel(\biu/bus_unit/mmu/mux10_b0_sel_is_2_o ),
    .o(\biu/bus_unit/mmu/n49 [2]));
  AL_MUX \biu/bus_unit/mmu/mux10_b3  (
    .i0(1'b0),
    .i1(\biu/bus_unit/mmu/statu [3]),
    .sel(\biu/bus_unit/mmu/mux10_b0_sel_is_2_o ),
    .o(\biu/bus_unit/mmu/n49 [3]));
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux11_b0  (
    .i0(\biu/bus_unit/mmu/n49 [0]),
    .i1(\biu/bus_unit/mmu/n46 [1]),
    .sel(\biu/bus_unit/mmu/n45 ),
    .o(\biu/bus_unit/mmu/n50 [0]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux11_b1  (
    .i0(\biu/bus_unit/mmu/n49 [1]),
    .i1(\biu/bus_unit/mmu/n46 [1]),
    .sel(\biu/bus_unit/mmu/n45 ),
    .o(\biu/bus_unit/mmu/n50 [1]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux11_b2  (
    .i0(\biu/bus_unit/mmu/n49 [2]),
    .i1(\biu/bus_unit/mmu/n46 [1]),
    .sel(\biu/bus_unit/mmu/n45 ),
    .o(\biu/bus_unit/mmu/n50 [2]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux11_b3  (
    .i0(\biu/bus_unit/mmu/n49 [3]),
    .i1(hresp),
    .sel(\biu/bus_unit/mmu/n45 ),
    .o(\biu/bus_unit/mmu/n50 [3]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux12_b0  (
    .i0(\biu/bus_unit/mmu/n50 [0]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu_hwrite ),
    .o(\biu/bus_unit/mmu/n51 [0]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux12_b1  (
    .i0(\biu/bus_unit/mmu/n50 [1]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu_hwrite ),
    .o(\biu/bus_unit/mmu/n51 [1]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux12_b2  (
    .i0(\biu/bus_unit/mmu/n50 [2]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu_hwrite ),
    .o(\biu/bus_unit/mmu/n51 [2]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux12_b3  (
    .i0(\biu/bus_unit/mmu/n50 [3]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu_hwrite ),
    .o(\biu/bus_unit/mmu/n51 [3]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux13_b0  (
    .i0(\biu/bus_unit/mmu/n51 [0]),
    .i1(\biu/bus_unit/mmu/n44 [0]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n52 [0]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux13_b1  (
    .i0(\biu/bus_unit/mmu/n51 [1]),
    .i1(\biu/bus_unit/mmu/n44 [1]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n52 [1]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux13_b2  (
    .i0(\biu/bus_unit/mmu/n51 [2]),
    .i1(\biu/bus_unit/mmu/n44 [0]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n52 [2]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux13_b3  (
    .i0(\biu/bus_unit/mmu/n51 [3]),
    .i1(\biu/bus_unit/mmu/n44 [3]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n52 [3]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux14_b0  (
    .i0(\biu/bus_unit/mmu/n52 [0]),
    .i1(\biu/bus_unit/mmu/n40 [0]),
    .sel(\biu/bus_unit/mmu/n37 ),
    .o(\biu/bus_unit/mmu/n53 [0]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux14_b1  (
    .i0(\biu/bus_unit/mmu/n52 [1]),
    .i1(\biu/bus_unit/mmu/n40 [1]),
    .sel(\biu/bus_unit/mmu/n37 ),
    .o(\biu/bus_unit/mmu/n53 [1]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux14_b2  (
    .i0(\biu/bus_unit/mmu/n52 [2]),
    .i1(\biu/bus_unit/mmu/n40 [2]),
    .sel(\biu/bus_unit/mmu/n37 ),
    .o(\biu/bus_unit/mmu/n53 [2]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux14_b3  (
    .i0(\biu/bus_unit/mmu/n52 [3]),
    .i1(\biu/bus_unit/mmu/n40 [3]),
    .sel(\biu/bus_unit/mmu/n37 ),
    .o(\biu/bus_unit/mmu/n53 [3]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux15_b0  (
    .i0(\biu/bus_unit/mmu/n53 [0]),
    .i1(\biu/bus_unit/mmu/n36 [0]),
    .sel(\biu/bus_unit/mmu/n35 ),
    .o(\biu/bus_unit/mmu/n54 [0]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux15_b1  (
    .i0(\biu/bus_unit/mmu/n53 [1]),
    .i1(\biu/bus_unit/mmu/n36 [1]),
    .sel(\biu/bus_unit/mmu/n35 ),
    .o(\biu/bus_unit/mmu/n54 [1]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux15_b3  (
    .i0(\biu/bus_unit/mmu/n53 [3]),
    .i1(\biu/bus_unit/mmu/n36 [3]),
    .sel(\biu/bus_unit/mmu/n35 ),
    .o(\biu/bus_unit/mmu/n54 [3]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux16_b0  (
    .i0(\biu/bus_unit/mmu/n54 [0]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n34 ),
    .o(\biu/bus_unit/mmu/n55 [0]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux16_b1  (
    .i0(\biu/bus_unit/mmu/n54 [1]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n34 ),
    .o(\biu/bus_unit/mmu/n55 [1]));  // ../../RTL/CPU/BIU/mmu.v(153)
  AL_MUX \biu/bus_unit/mmu/mux16_b2  (
    .i0(1'b0),
    .i1(\biu/bus_unit/mmu/n53 [2]),
    .sel(\biu/bus_unit/mmu/mux16_b2_sel_is_0_o ),
    .o(\biu/bus_unit/mmu/n55 [2]));
  and \biu/bus_unit/mmu/mux16_b2_sel_is_0  (\biu/bus_unit/mmu/mux16_b2_sel_is_0_o , \biu/bus_unit/mmu/n34_neg , \biu/bus_unit/mmu/n35_neg );
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux17_b0  (
    .i0(\biu/bus_unit/mmu/n55 [0]),
    .i1(\biu/bus_unit/mmu/n33 [0]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n56 [0]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux17_b1  (
    .i0(\biu/bus_unit/mmu/n55 [1]),
    .i1(\biu/bus_unit/mmu/n33 [1]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n56 [1]));  // ../../RTL/CPU/BIU/mmu.v(153)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux17_b2  (
    .i0(\biu/bus_unit/mmu/n55 [2]),
    .i1(\biu/bus_unit/mmu/n33 [1]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n56 [2]));  // ../../RTL/CPU/BIU/mmu.v(153)
  and \biu/bus_unit/mmu/mux17_b3_sel_is_0  (\biu/bus_unit/mmu/mux17_b3_sel_is_0_o , \biu/bus_unit/mmu/n30_neg , \biu/bus_unit/mmu/n34_neg );
  and \biu/bus_unit/mmu/mux18_b3_sel_is_2  (\biu/bus_unit/mmu/mux18_b3_sel_is_2_o , rst_neg, \biu/bus_unit/mmu/mux17_b3_sel_is_0_o );
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux1_b0  (
    .i0(\biu/bus_unit/mmu/n28 [0]),
    .i1(\biu/maddress [21]),
    .sel(\biu/bus_unit/mmu/n27 ),
    .o(\biu/bus_unit/mmu/n29 [0]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux1_b1  (
    .i0(\biu/bus_unit/mmu/n28 [1]),
    .i1(\biu/maddress [22]),
    .sel(\biu/bus_unit/mmu/n27 ),
    .o(\biu/bus_unit/mmu/n29 [1]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux1_b2  (
    .i0(\biu/bus_unit/mmu/n28 [2]),
    .i1(\biu/maddress [23]),
    .sel(\biu/bus_unit/mmu/n27 ),
    .o(\biu/bus_unit/mmu/n29 [2]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux1_b3  (
    .i0(\biu/bus_unit/mmu/n28 [3]),
    .i1(\biu/maddress [24]),
    .sel(\biu/bus_unit/mmu/n27 ),
    .o(\biu/bus_unit/mmu/n29 [3]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux1_b4  (
    .i0(\biu/bus_unit/mmu/n28 [4]),
    .i1(\biu/maddress [25]),
    .sel(\biu/bus_unit/mmu/n27 ),
    .o(\biu/bus_unit/mmu/n29 [4]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux1_b5  (
    .i0(\biu/bus_unit/mmu/n28 [5]),
    .i1(\biu/maddress [26]),
    .sel(\biu/bus_unit/mmu/n27 ),
    .o(\biu/bus_unit/mmu/n29 [5]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux1_b6  (
    .i0(\biu/bus_unit/mmu/n28 [6]),
    .i1(\biu/maddress [27]),
    .sel(\biu/bus_unit/mmu/n27 ),
    .o(\biu/bus_unit/mmu/n29 [6]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux1_b7  (
    .i0(\biu/bus_unit/mmu/n28 [7]),
    .i1(\biu/maddress [28]),
    .sel(\biu/bus_unit/mmu/n27 ),
    .o(\biu/bus_unit/mmu/n29 [7]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux1_b8  (
    .i0(\biu/bus_unit/mmu/n28 [8]),
    .i1(\biu/maddress [29]),
    .sel(\biu/bus_unit/mmu/n27 ),
    .o(\biu/bus_unit/mmu/n29 [8]));  // ../../RTL/CPU/BIU/mmu.v(115)
  and \biu/bus_unit/mmu/mux20_b0_sel_is_3  (\biu/bus_unit/mmu/mux20_b0_sel_is_3_o , \biu/bus_unit/mmu/n37 , \biu/bus_unit/mmu/pointer_page );
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b0  (
    .i0(\biu/paddress [0]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [0]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b1  (
    .i0(\biu/paddress [1]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [1]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b10  (
    .i0(\biu/paddress [10]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [10]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b11  (
    .i0(\biu/paddress [11]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [11]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b12  (
    .i0(\biu/paddress [12]),
    .i1(\biu/maddress [12]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [12]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b13  (
    .i0(\biu/paddress [13]),
    .i1(\biu/maddress [13]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [13]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b14  (
    .i0(\biu/paddress [14]),
    .i1(\biu/maddress [14]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [14]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b15  (
    .i0(\biu/paddress [15]),
    .i1(\biu/maddress [15]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [15]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b16  (
    .i0(\biu/paddress [16]),
    .i1(\biu/maddress [16]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [16]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b17  (
    .i0(\biu/paddress [17]),
    .i1(\biu/maddress [17]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [17]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b18  (
    .i0(\biu/paddress [18]),
    .i1(\biu/maddress [18]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [18]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b19  (
    .i0(\biu/paddress [19]),
    .i1(\biu/maddress [19]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [19]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b2  (
    .i0(\biu/paddress [2]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [2]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b20  (
    .i0(\biu/paddress [20]),
    .i1(\biu/maddress [20]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [20]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b21  (
    .i0(\biu/paddress [21]),
    .i1(\biu/maddress [21]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [21]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b22  (
    .i0(\biu/paddress [22]),
    .i1(\biu/maddress [22]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [22]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b23  (
    .i0(\biu/paddress [23]),
    .i1(\biu/maddress [23]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [23]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b24  (
    .i0(\biu/paddress [24]),
    .i1(\biu/maddress [24]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [24]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b25  (
    .i0(\biu/paddress [25]),
    .i1(\biu/maddress [25]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [25]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b26  (
    .i0(\biu/paddress [26]),
    .i1(\biu/maddress [26]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [26]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b27  (
    .i0(\biu/paddress [27]),
    .i1(\biu/maddress [27]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [27]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b28  (
    .i0(\biu/paddress [28]),
    .i1(\biu/maddress [28]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [28]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b29  (
    .i0(\biu/paddress [29]),
    .i1(\biu/maddress [29]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [29]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b3  (
    .i0(\biu/paddress [3]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [3]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b30  (
    .i0(\biu/paddress [30]),
    .i1(\biu/maddress [30]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [30]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b31  (
    .i0(\biu/paddress [31]),
    .i1(\biu/maddress [31]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [31]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b32  (
    .i0(\biu/paddress [32]),
    .i1(\biu/maddress [32]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [32]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b33  (
    .i0(\biu/paddress [33]),
    .i1(\biu/maddress [33]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [33]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b34  (
    .i0(\biu/paddress [34]),
    .i1(\biu/maddress [34]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [34]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b35  (
    .i0(\biu/paddress [35]),
    .i1(\biu/maddress [35]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [35]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b36  (
    .i0(\biu/paddress [36]),
    .i1(\biu/maddress [36]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [36]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b37  (
    .i0(\biu/paddress [37]),
    .i1(\biu/maddress [37]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [37]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b38  (
    .i0(\biu/paddress [38]),
    .i1(\biu/maddress [38]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [38]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b39  (
    .i0(\biu/paddress [39]),
    .i1(\biu/maddress [39]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [39]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b4  (
    .i0(\biu/paddress [4]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [4]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b40  (
    .i0(\biu/paddress [40]),
    .i1(\biu/maddress [40]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [40]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b41  (
    .i0(\biu/paddress [41]),
    .i1(\biu/maddress [41]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [41]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b42  (
    .i0(\biu/paddress [42]),
    .i1(\biu/maddress [42]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [42]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b43  (
    .i0(\biu/paddress [43]),
    .i1(\biu/maddress [43]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [43]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b44  (
    .i0(\biu/paddress [44]),
    .i1(\biu/maddress [44]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [44]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b45  (
    .i0(\biu/paddress [45]),
    .i1(\biu/maddress [45]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [45]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b46  (
    .i0(\biu/paddress [46]),
    .i1(\biu/maddress [46]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [46]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b47  (
    .i0(\biu/paddress [47]),
    .i1(\biu/maddress [47]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [47]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b48  (
    .i0(\biu/paddress [48]),
    .i1(\biu/maddress [48]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [48]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b49  (
    .i0(\biu/paddress [49]),
    .i1(\biu/maddress [49]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [49]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b5  (
    .i0(\biu/paddress [5]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [5]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b50  (
    .i0(\biu/paddress [50]),
    .i1(\biu/maddress [50]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [50]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b51  (
    .i0(\biu/paddress [51]),
    .i1(\biu/maddress [51]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [51]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b52  (
    .i0(\biu/paddress [52]),
    .i1(\biu/maddress [52]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [52]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b53  (
    .i0(\biu/paddress [53]),
    .i1(\biu/maddress [53]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [53]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b54  (
    .i0(\biu/paddress [54]),
    .i1(\biu/maddress [54]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [54]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b55  (
    .i0(\biu/paddress [55]),
    .i1(\biu/maddress [55]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [55]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b56  (
    .i0(\biu/paddress [56]),
    .i1(\biu/maddress [56]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [56]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b57  (
    .i0(\biu/paddress [57]),
    .i1(\biu/maddress [57]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [57]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b58  (
    .i0(\biu/paddress [58]),
    .i1(\biu/maddress [58]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [58]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b59  (
    .i0(\biu/paddress [59]),
    .i1(\biu/maddress [59]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [59]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b6  (
    .i0(\biu/paddress [6]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [6]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b60  (
    .i0(\biu/paddress [60]),
    .i1(\biu/maddress [60]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [60]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b61  (
    .i0(\biu/paddress [61]),
    .i1(\biu/maddress [61]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [61]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b62  (
    .i0(\biu/paddress [62]),
    .i1(\biu/maddress [62]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [62]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b63  (
    .i0(\biu/paddress [63]),
    .i1(\biu/maddress [63]),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [63]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b7  (
    .i0(\biu/paddress [7]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [7]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b8  (
    .i0(\biu/paddress [8]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [8]));  // ../../RTL/CPU/BIU/mmu.v(174)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux22_b9  (
    .i0(\biu/paddress [9]),
    .i1(1'b0),
    .sel(\biu/pa_cov ),
    .o(\biu/bus_unit/mmu/n63 [9]));  // ../../RTL/CPU/BIU/mmu.v(174)
  and \biu/bus_unit/mmu/mux23_b0_sel_is_3  (\biu/bus_unit/mmu/mux23_b0_sel_is_3_o , \biu/bus_unit/mmu/i [0], \biu/bus_unit/mmu/i [1]);
  not \biu/bus_unit/mmu/mux23_b0_sel_is_3_o_inv  (\biu/bus_unit/mmu/mux23_b0_sel_is_3_o_neg , \biu/bus_unit/mmu/mux23_b0_sel_is_3_o );
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b12  (
    .i0(\biu/bus_unit/mmu_hwdata [10]),
    .i1(\biu/maddress [12]),
    .i2(\biu/maddress [12]),
    .i3(\biu/paddress [12]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [12]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b13  (
    .i0(\biu/bus_unit/mmu_hwdata [11]),
    .i1(\biu/maddress [13]),
    .i2(\biu/maddress [13]),
    .i3(\biu/paddress [13]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [13]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b14  (
    .i0(\biu/bus_unit/mmu_hwdata [12]),
    .i1(\biu/maddress [14]),
    .i2(\biu/maddress [14]),
    .i3(\biu/paddress [14]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [14]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b15  (
    .i0(\biu/bus_unit/mmu_hwdata [13]),
    .i1(\biu/maddress [15]),
    .i2(\biu/maddress [15]),
    .i3(\biu/paddress [15]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [15]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b16  (
    .i0(\biu/bus_unit/mmu_hwdata [14]),
    .i1(\biu/maddress [16]),
    .i2(\biu/maddress [16]),
    .i3(\biu/paddress [16]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [16]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b17  (
    .i0(\biu/bus_unit/mmu_hwdata [15]),
    .i1(\biu/maddress [17]),
    .i2(\biu/maddress [17]),
    .i3(\biu/paddress [17]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [17]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b18  (
    .i0(\biu/bus_unit/mmu_hwdata [16]),
    .i1(\biu/maddress [18]),
    .i2(\biu/maddress [18]),
    .i3(\biu/paddress [18]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [18]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b19  (
    .i0(\biu/bus_unit/mmu_hwdata [17]),
    .i1(\biu/maddress [19]),
    .i2(\biu/maddress [19]),
    .i3(\biu/paddress [19]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [19]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b20  (
    .i0(\biu/bus_unit/mmu_hwdata [18]),
    .i1(\biu/maddress [20]),
    .i2(\biu/maddress [20]),
    .i3(\biu/paddress [20]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [20]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b21  (
    .i0(\biu/bus_unit/mmu_hwdata [19]),
    .i1(\biu/bus_unit/mmu_hwdata [19]),
    .i2(\biu/maddress [21]),
    .i3(\biu/paddress [21]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [21]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b22  (
    .i0(\biu/bus_unit/mmu_hwdata [20]),
    .i1(\biu/bus_unit/mmu_hwdata [20]),
    .i2(\biu/maddress [22]),
    .i3(\biu/paddress [22]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [22]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b23  (
    .i0(\biu/bus_unit/mmu_hwdata [21]),
    .i1(\biu/bus_unit/mmu_hwdata [21]),
    .i2(\biu/maddress [23]),
    .i3(\biu/paddress [23]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [23]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b24  (
    .i0(\biu/bus_unit/mmu_hwdata [22]),
    .i1(\biu/bus_unit/mmu_hwdata [22]),
    .i2(\biu/maddress [24]),
    .i3(\biu/paddress [24]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [24]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b25  (
    .i0(\biu/bus_unit/mmu_hwdata [23]),
    .i1(\biu/bus_unit/mmu_hwdata [23]),
    .i2(\biu/maddress [25]),
    .i3(\biu/paddress [25]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [25]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b26  (
    .i0(\biu/bus_unit/mmu_hwdata [24]),
    .i1(\biu/bus_unit/mmu_hwdata [24]),
    .i2(\biu/maddress [26]),
    .i3(\biu/paddress [26]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [26]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b27  (
    .i0(\biu/bus_unit/mmu_hwdata [25]),
    .i1(\biu/bus_unit/mmu_hwdata [25]),
    .i2(\biu/maddress [27]),
    .i3(\biu/paddress [27]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [27]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b28  (
    .i0(\biu/bus_unit/mmu_hwdata [26]),
    .i1(\biu/bus_unit/mmu_hwdata [26]),
    .i2(\biu/maddress [28]),
    .i3(\biu/paddress [28]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [28]));  // ../../RTL/CPU/BIU/mmu.v(181)
  binary_mux_s2_w1 \biu/bus_unit/mmu/mux23_b29  (
    .i0(\biu/bus_unit/mmu_hwdata [27]),
    .i1(\biu/bus_unit/mmu_hwdata [27]),
    .i2(\biu/maddress [29]),
    .i3(\biu/paddress [29]),
    .sel(\biu/bus_unit/mmu/i ),
    .o(\biu/bus_unit/mmu/n64 [29]));  // ../../RTL/CPU/BIU/mmu.v(181)
  AL_MUX \biu/bus_unit/mmu/mux24_b0  (
    .i0(\biu/paddress [0]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [0]));
  and \biu/bus_unit/mmu/mux24_b0_sel_is_1  (\biu/bus_unit/mmu/mux24_b0_sel_is_1_o , \biu/bus_unit/mmu/n41 , \biu/bus_unit/mmu/mux23_b0_sel_is_3_o_neg );
  AL_MUX \biu/bus_unit/mmu/mux24_b1  (
    .i0(\biu/paddress [1]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [1]));
  AL_MUX \biu/bus_unit/mmu/mux24_b10  (
    .i0(\biu/paddress [10]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [10]));
  AL_MUX \biu/bus_unit/mmu/mux24_b11  (
    .i0(\biu/paddress [11]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [11]));
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b12  (
    .i0(\biu/paddress [12]),
    .i1(\biu/bus_unit/mmu/n64 [12]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [12]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b13  (
    .i0(\biu/paddress [13]),
    .i1(\biu/bus_unit/mmu/n64 [13]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [13]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b14  (
    .i0(\biu/paddress [14]),
    .i1(\biu/bus_unit/mmu/n64 [14]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [14]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b15  (
    .i0(\biu/paddress [15]),
    .i1(\biu/bus_unit/mmu/n64 [15]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [15]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b16  (
    .i0(\biu/paddress [16]),
    .i1(\biu/bus_unit/mmu/n64 [16]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [16]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b17  (
    .i0(\biu/paddress [17]),
    .i1(\biu/bus_unit/mmu/n64 [17]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [17]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b18  (
    .i0(\biu/paddress [18]),
    .i1(\biu/bus_unit/mmu/n64 [18]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [18]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b19  (
    .i0(\biu/paddress [19]),
    .i1(\biu/bus_unit/mmu/n64 [19]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [19]));  // ../../RTL/CPU/BIU/mmu.v(182)
  AL_MUX \biu/bus_unit/mmu/mux24_b2  (
    .i0(\biu/paddress [2]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [2]));
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b20  (
    .i0(\biu/paddress [20]),
    .i1(\biu/bus_unit/mmu/n64 [20]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [20]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b21  (
    .i0(\biu/paddress [21]),
    .i1(\biu/bus_unit/mmu/n64 [21]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [21]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b22  (
    .i0(\biu/paddress [22]),
    .i1(\biu/bus_unit/mmu/n64 [22]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [22]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b23  (
    .i0(\biu/paddress [23]),
    .i1(\biu/bus_unit/mmu/n64 [23]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [23]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b24  (
    .i0(\biu/paddress [24]),
    .i1(\biu/bus_unit/mmu/n64 [24]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [24]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b25  (
    .i0(\biu/paddress [25]),
    .i1(\biu/bus_unit/mmu/n64 [25]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [25]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b26  (
    .i0(\biu/paddress [26]),
    .i1(\biu/bus_unit/mmu/n64 [26]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [26]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b27  (
    .i0(\biu/paddress [27]),
    .i1(\biu/bus_unit/mmu/n64 [27]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [27]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b28  (
    .i0(\biu/paddress [28]),
    .i1(\biu/bus_unit/mmu/n64 [28]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [28]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux24_b29  (
    .i0(\biu/paddress [29]),
    .i1(\biu/bus_unit/mmu/n64 [29]),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n65 [29]));  // ../../RTL/CPU/BIU/mmu.v(182)
  AL_MUX \biu/bus_unit/mmu/mux24_b3  (
    .i0(\biu/paddress [3]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [3]));
  AL_MUX \biu/bus_unit/mmu/mux24_b30  (
    .i0(\biu/paddress [30]),
    .i1(\biu/bus_unit/mmu_hwdata [28]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [30]));
  AL_MUX \biu/bus_unit/mmu/mux24_b31  (
    .i0(\biu/paddress [31]),
    .i1(\biu/bus_unit/mmu_hwdata [29]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [31]));
  AL_MUX \biu/bus_unit/mmu/mux24_b32  (
    .i0(\biu/paddress [32]),
    .i1(\biu/bus_unit/mmu_hwdata [30]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [32]));
  AL_MUX \biu/bus_unit/mmu/mux24_b33  (
    .i0(\biu/paddress [33]),
    .i1(\biu/bus_unit/mmu_hwdata [31]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [33]));
  AL_MUX \biu/bus_unit/mmu/mux24_b34  (
    .i0(\biu/paddress [34]),
    .i1(\biu/bus_unit/mmu_hwdata [32]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [34]));
  AL_MUX \biu/bus_unit/mmu/mux24_b35  (
    .i0(\biu/paddress [35]),
    .i1(\biu/bus_unit/mmu_hwdata [33]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [35]));
  AL_MUX \biu/bus_unit/mmu/mux24_b36  (
    .i0(\biu/paddress [36]),
    .i1(\biu/bus_unit/mmu_hwdata [34]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [36]));
  AL_MUX \biu/bus_unit/mmu/mux24_b37  (
    .i0(\biu/paddress [37]),
    .i1(\biu/bus_unit/mmu_hwdata [35]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [37]));
  AL_MUX \biu/bus_unit/mmu/mux24_b38  (
    .i0(\biu/paddress [38]),
    .i1(\biu/bus_unit/mmu_hwdata [36]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [38]));
  AL_MUX \biu/bus_unit/mmu/mux24_b39  (
    .i0(\biu/paddress [39]),
    .i1(\biu/bus_unit/mmu_hwdata [37]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [39]));
  AL_MUX \biu/bus_unit/mmu/mux24_b4  (
    .i0(\biu/paddress [4]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [4]));
  AL_MUX \biu/bus_unit/mmu/mux24_b40  (
    .i0(\biu/paddress [40]),
    .i1(\biu/bus_unit/mmu_hwdata [38]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [40]));
  AL_MUX \biu/bus_unit/mmu/mux24_b41  (
    .i0(\biu/paddress [41]),
    .i1(\biu/bus_unit/mmu_hwdata [39]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [41]));
  AL_MUX \biu/bus_unit/mmu/mux24_b42  (
    .i0(\biu/paddress [42]),
    .i1(\biu/bus_unit/mmu_hwdata [40]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [42]));
  AL_MUX \biu/bus_unit/mmu/mux24_b43  (
    .i0(\biu/paddress [43]),
    .i1(\biu/bus_unit/mmu_hwdata [41]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [43]));
  AL_MUX \biu/bus_unit/mmu/mux24_b44  (
    .i0(\biu/paddress [44]),
    .i1(\biu/bus_unit/mmu_hwdata [42]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [44]));
  AL_MUX \biu/bus_unit/mmu/mux24_b45  (
    .i0(\biu/paddress [45]),
    .i1(\biu/bus_unit/mmu_hwdata [43]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [45]));
  AL_MUX \biu/bus_unit/mmu/mux24_b46  (
    .i0(\biu/paddress [46]),
    .i1(\biu/bus_unit/mmu_hwdata [44]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [46]));
  AL_MUX \biu/bus_unit/mmu/mux24_b47  (
    .i0(\biu/paddress [47]),
    .i1(\biu/bus_unit/mmu_hwdata [45]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [47]));
  AL_MUX \biu/bus_unit/mmu/mux24_b48  (
    .i0(\biu/paddress [48]),
    .i1(\biu/bus_unit/mmu_hwdata [46]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [48]));
  AL_MUX \biu/bus_unit/mmu/mux24_b49  (
    .i0(\biu/paddress [49]),
    .i1(\biu/bus_unit/mmu_hwdata [47]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [49]));
  AL_MUX \biu/bus_unit/mmu/mux24_b5  (
    .i0(\biu/paddress [5]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [5]));
  AL_MUX \biu/bus_unit/mmu/mux24_b50  (
    .i0(\biu/paddress [50]),
    .i1(\biu/bus_unit/mmu_hwdata [48]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [50]));
  AL_MUX \biu/bus_unit/mmu/mux24_b51  (
    .i0(\biu/paddress [51]),
    .i1(\biu/bus_unit/mmu_hwdata [49]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [51]));
  AL_MUX \biu/bus_unit/mmu/mux24_b52  (
    .i0(\biu/paddress [52]),
    .i1(\biu/bus_unit/mmu_hwdata [50]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [52]));
  AL_MUX \biu/bus_unit/mmu/mux24_b53  (
    .i0(\biu/paddress [53]),
    .i1(\biu/bus_unit/mmu_hwdata [51]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [53]));
  AL_MUX \biu/bus_unit/mmu/mux24_b54  (
    .i0(\biu/paddress [54]),
    .i1(\biu/bus_unit/mmu_hwdata [52]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [54]));
  AL_MUX \biu/bus_unit/mmu/mux24_b55  (
    .i0(\biu/paddress [55]),
    .i1(\biu/bus_unit/mmu_hwdata [53]),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [55]));
  AL_MUX \biu/bus_unit/mmu/mux24_b56  (
    .i0(\biu/paddress [56]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [56]));
  AL_MUX \biu/bus_unit/mmu/mux24_b57  (
    .i0(\biu/paddress [57]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [57]));
  AL_MUX \biu/bus_unit/mmu/mux24_b58  (
    .i0(\biu/paddress [58]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [58]));
  AL_MUX \biu/bus_unit/mmu/mux24_b59  (
    .i0(\biu/paddress [59]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [59]));
  AL_MUX \biu/bus_unit/mmu/mux24_b6  (
    .i0(\biu/paddress [6]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [6]));
  AL_MUX \biu/bus_unit/mmu/mux24_b60  (
    .i0(\biu/paddress [60]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [60]));
  AL_MUX \biu/bus_unit/mmu/mux24_b61  (
    .i0(\biu/paddress [61]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [61]));
  AL_MUX \biu/bus_unit/mmu/mux24_b62  (
    .i0(\biu/paddress [62]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [62]));
  AL_MUX \biu/bus_unit/mmu/mux24_b63  (
    .i0(\biu/paddress [63]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [63]));
  AL_MUX \biu/bus_unit/mmu/mux24_b7  (
    .i0(\biu/paddress [7]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [7]));
  AL_MUX \biu/bus_unit/mmu/mux24_b8  (
    .i0(\biu/paddress [8]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [8]));
  AL_MUX \biu/bus_unit/mmu/mux24_b9  (
    .i0(\biu/paddress [9]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux24_b0_sel_is_1_o ),
    .o(\biu/bus_unit/mmu/n65 [9]));
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b0  (
    .i0(\biu/bus_unit/mmu/n65 [0]),
    .i1(\biu/bus_unit/mmu/n63 [0]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [0]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b1  (
    .i0(\biu/bus_unit/mmu/n65 [1]),
    .i1(\biu/bus_unit/mmu/n63 [1]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [1]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b10  (
    .i0(\biu/bus_unit/mmu/n65 [10]),
    .i1(\biu/bus_unit/mmu/n63 [10]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [10]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b11  (
    .i0(\biu/bus_unit/mmu/n65 [11]),
    .i1(\biu/bus_unit/mmu/n63 [11]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [11]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b12  (
    .i0(\biu/bus_unit/mmu/n65 [12]),
    .i1(\biu/bus_unit/mmu/n63 [12]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [12]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b13  (
    .i0(\biu/bus_unit/mmu/n65 [13]),
    .i1(\biu/bus_unit/mmu/n63 [13]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [13]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b14  (
    .i0(\biu/bus_unit/mmu/n65 [14]),
    .i1(\biu/bus_unit/mmu/n63 [14]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [14]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b15  (
    .i0(\biu/bus_unit/mmu/n65 [15]),
    .i1(\biu/bus_unit/mmu/n63 [15]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [15]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b16  (
    .i0(\biu/bus_unit/mmu/n65 [16]),
    .i1(\biu/bus_unit/mmu/n63 [16]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [16]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b17  (
    .i0(\biu/bus_unit/mmu/n65 [17]),
    .i1(\biu/bus_unit/mmu/n63 [17]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [17]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b18  (
    .i0(\biu/bus_unit/mmu/n65 [18]),
    .i1(\biu/bus_unit/mmu/n63 [18]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [18]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b19  (
    .i0(\biu/bus_unit/mmu/n65 [19]),
    .i1(\biu/bus_unit/mmu/n63 [19]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [19]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b2  (
    .i0(\biu/bus_unit/mmu/n65 [2]),
    .i1(\biu/bus_unit/mmu/n63 [2]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [2]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b20  (
    .i0(\biu/bus_unit/mmu/n65 [20]),
    .i1(\biu/bus_unit/mmu/n63 [20]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [20]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b21  (
    .i0(\biu/bus_unit/mmu/n65 [21]),
    .i1(\biu/bus_unit/mmu/n63 [21]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [21]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b22  (
    .i0(\biu/bus_unit/mmu/n65 [22]),
    .i1(\biu/bus_unit/mmu/n63 [22]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [22]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b23  (
    .i0(\biu/bus_unit/mmu/n65 [23]),
    .i1(\biu/bus_unit/mmu/n63 [23]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [23]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b24  (
    .i0(\biu/bus_unit/mmu/n65 [24]),
    .i1(\biu/bus_unit/mmu/n63 [24]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [24]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b25  (
    .i0(\biu/bus_unit/mmu/n65 [25]),
    .i1(\biu/bus_unit/mmu/n63 [25]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [25]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b26  (
    .i0(\biu/bus_unit/mmu/n65 [26]),
    .i1(\biu/bus_unit/mmu/n63 [26]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [26]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b27  (
    .i0(\biu/bus_unit/mmu/n65 [27]),
    .i1(\biu/bus_unit/mmu/n63 [27]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [27]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b28  (
    .i0(\biu/bus_unit/mmu/n65 [28]),
    .i1(\biu/bus_unit/mmu/n63 [28]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [28]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b29  (
    .i0(\biu/bus_unit/mmu/n65 [29]),
    .i1(\biu/bus_unit/mmu/n63 [29]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [29]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b3  (
    .i0(\biu/bus_unit/mmu/n65 [3]),
    .i1(\biu/bus_unit/mmu/n63 [3]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [3]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b30  (
    .i0(\biu/bus_unit/mmu/n65 [30]),
    .i1(\biu/bus_unit/mmu/n63 [30]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [30]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b31  (
    .i0(\biu/bus_unit/mmu/n65 [31]),
    .i1(\biu/bus_unit/mmu/n63 [31]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [31]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b32  (
    .i0(\biu/bus_unit/mmu/n65 [32]),
    .i1(\biu/bus_unit/mmu/n63 [32]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [32]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b33  (
    .i0(\biu/bus_unit/mmu/n65 [33]),
    .i1(\biu/bus_unit/mmu/n63 [33]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [33]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b34  (
    .i0(\biu/bus_unit/mmu/n65 [34]),
    .i1(\biu/bus_unit/mmu/n63 [34]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [34]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b35  (
    .i0(\biu/bus_unit/mmu/n65 [35]),
    .i1(\biu/bus_unit/mmu/n63 [35]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [35]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b36  (
    .i0(\biu/bus_unit/mmu/n65 [36]),
    .i1(\biu/bus_unit/mmu/n63 [36]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [36]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b37  (
    .i0(\biu/bus_unit/mmu/n65 [37]),
    .i1(\biu/bus_unit/mmu/n63 [37]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [37]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b38  (
    .i0(\biu/bus_unit/mmu/n65 [38]),
    .i1(\biu/bus_unit/mmu/n63 [38]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [38]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b39  (
    .i0(\biu/bus_unit/mmu/n65 [39]),
    .i1(\biu/bus_unit/mmu/n63 [39]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [39]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b4  (
    .i0(\biu/bus_unit/mmu/n65 [4]),
    .i1(\biu/bus_unit/mmu/n63 [4]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [4]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b40  (
    .i0(\biu/bus_unit/mmu/n65 [40]),
    .i1(\biu/bus_unit/mmu/n63 [40]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [40]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b41  (
    .i0(\biu/bus_unit/mmu/n65 [41]),
    .i1(\biu/bus_unit/mmu/n63 [41]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [41]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b42  (
    .i0(\biu/bus_unit/mmu/n65 [42]),
    .i1(\biu/bus_unit/mmu/n63 [42]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [42]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b43  (
    .i0(\biu/bus_unit/mmu/n65 [43]),
    .i1(\biu/bus_unit/mmu/n63 [43]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [43]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b44  (
    .i0(\biu/bus_unit/mmu/n65 [44]),
    .i1(\biu/bus_unit/mmu/n63 [44]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [44]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b45  (
    .i0(\biu/bus_unit/mmu/n65 [45]),
    .i1(\biu/bus_unit/mmu/n63 [45]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [45]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b46  (
    .i0(\biu/bus_unit/mmu/n65 [46]),
    .i1(\biu/bus_unit/mmu/n63 [46]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [46]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b47  (
    .i0(\biu/bus_unit/mmu/n65 [47]),
    .i1(\biu/bus_unit/mmu/n63 [47]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [47]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b48  (
    .i0(\biu/bus_unit/mmu/n65 [48]),
    .i1(\biu/bus_unit/mmu/n63 [48]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [48]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b49  (
    .i0(\biu/bus_unit/mmu/n65 [49]),
    .i1(\biu/bus_unit/mmu/n63 [49]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [49]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b5  (
    .i0(\biu/bus_unit/mmu/n65 [5]),
    .i1(\biu/bus_unit/mmu/n63 [5]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [5]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b50  (
    .i0(\biu/bus_unit/mmu/n65 [50]),
    .i1(\biu/bus_unit/mmu/n63 [50]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [50]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b51  (
    .i0(\biu/bus_unit/mmu/n65 [51]),
    .i1(\biu/bus_unit/mmu/n63 [51]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [51]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b52  (
    .i0(\biu/bus_unit/mmu/n65 [52]),
    .i1(\biu/bus_unit/mmu/n63 [52]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [52]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b53  (
    .i0(\biu/bus_unit/mmu/n65 [53]),
    .i1(\biu/bus_unit/mmu/n63 [53]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [53]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b54  (
    .i0(\biu/bus_unit/mmu/n65 [54]),
    .i1(\biu/bus_unit/mmu/n63 [54]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [54]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b55  (
    .i0(\biu/bus_unit/mmu/n65 [55]),
    .i1(\biu/bus_unit/mmu/n63 [55]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [55]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b56  (
    .i0(\biu/bus_unit/mmu/n65 [56]),
    .i1(\biu/bus_unit/mmu/n63 [56]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [56]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b57  (
    .i0(\biu/bus_unit/mmu/n65 [57]),
    .i1(\biu/bus_unit/mmu/n63 [57]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [57]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b58  (
    .i0(\biu/bus_unit/mmu/n65 [58]),
    .i1(\biu/bus_unit/mmu/n63 [58]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [58]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b59  (
    .i0(\biu/bus_unit/mmu/n65 [59]),
    .i1(\biu/bus_unit/mmu/n63 [59]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [59]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b6  (
    .i0(\biu/bus_unit/mmu/n65 [6]),
    .i1(\biu/bus_unit/mmu/n63 [6]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [6]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b60  (
    .i0(\biu/bus_unit/mmu/n65 [60]),
    .i1(\biu/bus_unit/mmu/n63 [60]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [60]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b61  (
    .i0(\biu/bus_unit/mmu/n65 [61]),
    .i1(\biu/bus_unit/mmu/n63 [61]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [61]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b62  (
    .i0(\biu/bus_unit/mmu/n65 [62]),
    .i1(\biu/bus_unit/mmu/n63 [62]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [62]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b63  (
    .i0(\biu/bus_unit/mmu/n65 [63]),
    .i1(\biu/bus_unit/mmu/n63 [63]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [63]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b7  (
    .i0(\biu/bus_unit/mmu/n65 [7]),
    .i1(\biu/bus_unit/mmu/n63 [7]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [7]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b8  (
    .i0(\biu/bus_unit/mmu/n65 [8]),
    .i1(\biu/bus_unit/mmu/n63 [8]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [8]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux25_b9  (
    .i0(\biu/bus_unit/mmu/n65 [9]),
    .i1(\biu/bus_unit/mmu/n63 [9]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n66 [9]));  // ../../RTL/CPU/BIU/mmu.v(182)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b0  (
    .i0(\biu/paddress [64]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [0]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b1  (
    .i0(\biu/paddress [65]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [1]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b10  (
    .i0(\biu/paddress [74]),
    .i1(\biu/bus_unit/mmu/va_vpn [7]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [10]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b11  (
    .i0(\biu/paddress [75]),
    .i1(\biu/bus_unit/mmu/va_vpn [8]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [11]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b12  (
    .i0(\biu/paddress [76]),
    .i1(satp[0]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [12]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b13  (
    .i0(\biu/paddress [77]),
    .i1(satp[1]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [13]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b14  (
    .i0(\biu/paddress [78]),
    .i1(satp[2]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [14]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b15  (
    .i0(\biu/paddress [79]),
    .i1(satp[3]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [15]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b16  (
    .i0(\biu/paddress [80]),
    .i1(satp[4]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [16]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b17  (
    .i0(\biu/paddress [81]),
    .i1(satp[5]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [17]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b18  (
    .i0(\biu/paddress [82]),
    .i1(satp[6]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [18]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b19  (
    .i0(\biu/paddress [83]),
    .i1(satp[7]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [19]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b2  (
    .i0(\biu/paddress [66]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [2]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b20  (
    .i0(\biu/paddress [84]),
    .i1(satp[8]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [20]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b21  (
    .i0(\biu/paddress [85]),
    .i1(satp[9]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [21]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b22  (
    .i0(\biu/paddress [86]),
    .i1(satp[10]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [22]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b23  (
    .i0(\biu/paddress [87]),
    .i1(satp[11]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [23]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b24  (
    .i0(\biu/paddress [88]),
    .i1(satp[12]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [24]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b25  (
    .i0(\biu/paddress [89]),
    .i1(satp[13]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [25]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b26  (
    .i0(\biu/paddress [90]),
    .i1(satp[14]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [26]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b27  (
    .i0(\biu/paddress [91]),
    .i1(satp[15]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [27]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b28  (
    .i0(\biu/paddress [92]),
    .i1(satp[16]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [28]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b29  (
    .i0(\biu/paddress [93]),
    .i1(satp[17]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [29]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b3  (
    .i0(\biu/paddress [67]),
    .i1(\biu/bus_unit/mmu/va_vpn [0]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [3]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b30  (
    .i0(\biu/paddress [94]),
    .i1(satp[18]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [30]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b31  (
    .i0(\biu/paddress [95]),
    .i1(satp[19]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [31]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b32  (
    .i0(\biu/paddress [96]),
    .i1(satp[20]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [32]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b33  (
    .i0(\biu/paddress [97]),
    .i1(satp[21]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [33]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b34  (
    .i0(\biu/paddress [98]),
    .i1(satp[22]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [34]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b35  (
    .i0(\biu/paddress [99]),
    .i1(satp[23]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [35]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b36  (
    .i0(\biu/paddress [100]),
    .i1(satp[24]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [36]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b37  (
    .i0(\biu/paddress [101]),
    .i1(satp[25]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [37]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b38  (
    .i0(\biu/paddress [102]),
    .i1(satp[26]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [38]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b39  (
    .i0(\biu/paddress [103]),
    .i1(satp[27]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [39]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b4  (
    .i0(\biu/paddress [68]),
    .i1(\biu/bus_unit/mmu/va_vpn [1]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [4]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b40  (
    .i0(\biu/paddress [104]),
    .i1(satp[28]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [40]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b41  (
    .i0(\biu/paddress [105]),
    .i1(satp[29]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [41]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b42  (
    .i0(\biu/paddress [106]),
    .i1(satp[30]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [42]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b43  (
    .i0(\biu/paddress [107]),
    .i1(satp[31]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [43]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b44  (
    .i0(\biu/paddress [108]),
    .i1(satp[32]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [44]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b45  (
    .i0(\biu/paddress [109]),
    .i1(satp[33]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [45]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b46  (
    .i0(\biu/paddress [110]),
    .i1(satp[34]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [46]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b47  (
    .i0(\biu/paddress [111]),
    .i1(satp[35]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [47]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b48  (
    .i0(\biu/paddress [112]),
    .i1(satp[36]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [48]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b49  (
    .i0(\biu/paddress [113]),
    .i1(satp[37]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [49]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b5  (
    .i0(\biu/paddress [69]),
    .i1(\biu/bus_unit/mmu/va_vpn [2]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [5]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b50  (
    .i0(\biu/paddress [114]),
    .i1(satp[38]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [50]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b51  (
    .i0(\biu/paddress [115]),
    .i1(satp[39]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [51]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b52  (
    .i0(\biu/paddress [116]),
    .i1(satp[40]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [52]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b53  (
    .i0(\biu/paddress [117]),
    .i1(satp[41]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [53]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b54  (
    .i0(\biu/paddress [118]),
    .i1(satp[42]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [54]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b55  (
    .i0(\biu/paddress [119]),
    .i1(satp[43]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [55]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b56  (
    .i0(\biu/paddress [120]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [56]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b57  (
    .i0(\biu/paddress [121]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [57]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b58  (
    .i0(\biu/paddress [122]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [58]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b59  (
    .i0(\biu/paddress [123]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [59]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b6  (
    .i0(\biu/paddress [70]),
    .i1(\biu/bus_unit/mmu/va_vpn [3]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [6]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b60  (
    .i0(\biu/paddress [124]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [60]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b61  (
    .i0(\biu/paddress [125]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [61]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b62  (
    .i0(\biu/paddress [126]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [62]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b63  (
    .i0(\biu/paddress [127]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [63]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b7  (
    .i0(\biu/paddress [71]),
    .i1(\biu/bus_unit/mmu/va_vpn [4]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [7]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b8  (
    .i0(\biu/paddress [72]),
    .i1(\biu/bus_unit/mmu/va_vpn [5]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [8]));  // ../../RTL/CPU/BIU/mmu.v(193)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux27_b9  (
    .i0(\biu/paddress [73]),
    .i1(\biu/bus_unit/mmu/va_vpn [6]),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n68 [9]));  // ../../RTL/CPU/BIU/mmu.v(193)
  AL_MUX \biu/bus_unit/mmu/mux29_b0  (
    .i0(\biu/paddress [64]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [0]));
  AL_MUX \biu/bus_unit/mmu/mux29_b1  (
    .i0(\biu/paddress [65]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [1]));
  AL_MUX \biu/bus_unit/mmu/mux29_b10  (
    .i0(\biu/paddress [74]),
    .i1(\biu/bus_unit/mmu/va_vpn [7]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [10]));
  AL_MUX \biu/bus_unit/mmu/mux29_b11  (
    .i0(\biu/paddress [75]),
    .i1(\biu/bus_unit/mmu/va_vpn [8]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [11]));
  AL_MUX \biu/bus_unit/mmu/mux29_b12  (
    .i0(\biu/paddress [76]),
    .i1(\biu/bus_unit/mmu_hwdata [10]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [12]));
  AL_MUX \biu/bus_unit/mmu/mux29_b13  (
    .i0(\biu/paddress [77]),
    .i1(\biu/bus_unit/mmu_hwdata [11]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [13]));
  AL_MUX \biu/bus_unit/mmu/mux29_b14  (
    .i0(\biu/paddress [78]),
    .i1(\biu/bus_unit/mmu_hwdata [12]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [14]));
  AL_MUX \biu/bus_unit/mmu/mux29_b15  (
    .i0(\biu/paddress [79]),
    .i1(\biu/bus_unit/mmu_hwdata [13]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [15]));
  AL_MUX \biu/bus_unit/mmu/mux29_b16  (
    .i0(\biu/paddress [80]),
    .i1(\biu/bus_unit/mmu_hwdata [14]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [16]));
  AL_MUX \biu/bus_unit/mmu/mux29_b17  (
    .i0(\biu/paddress [81]),
    .i1(\biu/bus_unit/mmu_hwdata [15]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [17]));
  AL_MUX \biu/bus_unit/mmu/mux29_b18  (
    .i0(\biu/paddress [82]),
    .i1(\biu/bus_unit/mmu_hwdata [16]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [18]));
  AL_MUX \biu/bus_unit/mmu/mux29_b19  (
    .i0(\biu/paddress [83]),
    .i1(\biu/bus_unit/mmu_hwdata [17]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [19]));
  AL_MUX \biu/bus_unit/mmu/mux29_b2  (
    .i0(\biu/paddress [66]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [2]));
  AL_MUX \biu/bus_unit/mmu/mux29_b20  (
    .i0(\biu/paddress [84]),
    .i1(\biu/bus_unit/mmu_hwdata [18]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [20]));
  AL_MUX \biu/bus_unit/mmu/mux29_b21  (
    .i0(\biu/paddress [85]),
    .i1(\biu/bus_unit/mmu_hwdata [19]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [21]));
  AL_MUX \biu/bus_unit/mmu/mux29_b22  (
    .i0(\biu/paddress [86]),
    .i1(\biu/bus_unit/mmu_hwdata [20]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [22]));
  AL_MUX \biu/bus_unit/mmu/mux29_b23  (
    .i0(\biu/paddress [87]),
    .i1(\biu/bus_unit/mmu_hwdata [21]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [23]));
  AL_MUX \biu/bus_unit/mmu/mux29_b24  (
    .i0(\biu/paddress [88]),
    .i1(\biu/bus_unit/mmu_hwdata [22]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [24]));
  AL_MUX \biu/bus_unit/mmu/mux29_b25  (
    .i0(\biu/paddress [89]),
    .i1(\biu/bus_unit/mmu_hwdata [23]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [25]));
  AL_MUX \biu/bus_unit/mmu/mux29_b26  (
    .i0(\biu/paddress [90]),
    .i1(\biu/bus_unit/mmu_hwdata [24]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [26]));
  AL_MUX \biu/bus_unit/mmu/mux29_b27  (
    .i0(\biu/paddress [91]),
    .i1(\biu/bus_unit/mmu_hwdata [25]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [27]));
  AL_MUX \biu/bus_unit/mmu/mux29_b28  (
    .i0(\biu/paddress [92]),
    .i1(\biu/bus_unit/mmu_hwdata [26]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [28]));
  AL_MUX \biu/bus_unit/mmu/mux29_b29  (
    .i0(\biu/paddress [93]),
    .i1(\biu/bus_unit/mmu_hwdata [27]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [29]));
  AL_MUX \biu/bus_unit/mmu/mux29_b3  (
    .i0(\biu/paddress [67]),
    .i1(\biu/bus_unit/mmu/va_vpn [0]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [3]));
  AL_MUX \biu/bus_unit/mmu/mux29_b30  (
    .i0(\biu/paddress [94]),
    .i1(\biu/bus_unit/mmu_hwdata [28]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [30]));
  AL_MUX \biu/bus_unit/mmu/mux29_b31  (
    .i0(\biu/paddress [95]),
    .i1(\biu/bus_unit/mmu_hwdata [29]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [31]));
  AL_MUX \biu/bus_unit/mmu/mux29_b32  (
    .i0(\biu/paddress [96]),
    .i1(\biu/bus_unit/mmu_hwdata [30]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [32]));
  AL_MUX \biu/bus_unit/mmu/mux29_b33  (
    .i0(\biu/paddress [97]),
    .i1(\biu/bus_unit/mmu_hwdata [31]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [33]));
  AL_MUX \biu/bus_unit/mmu/mux29_b34  (
    .i0(\biu/paddress [98]),
    .i1(\biu/bus_unit/mmu_hwdata [32]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [34]));
  AL_MUX \biu/bus_unit/mmu/mux29_b35  (
    .i0(\biu/paddress [99]),
    .i1(\biu/bus_unit/mmu_hwdata [33]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [35]));
  AL_MUX \biu/bus_unit/mmu/mux29_b36  (
    .i0(\biu/paddress [100]),
    .i1(\biu/bus_unit/mmu_hwdata [34]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [36]));
  AL_MUX \biu/bus_unit/mmu/mux29_b37  (
    .i0(\biu/paddress [101]),
    .i1(\biu/bus_unit/mmu_hwdata [35]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [37]));
  AL_MUX \biu/bus_unit/mmu/mux29_b38  (
    .i0(\biu/paddress [102]),
    .i1(\biu/bus_unit/mmu_hwdata [36]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [38]));
  AL_MUX \biu/bus_unit/mmu/mux29_b39  (
    .i0(\biu/paddress [103]),
    .i1(\biu/bus_unit/mmu_hwdata [37]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [39]));
  AL_MUX \biu/bus_unit/mmu/mux29_b4  (
    .i0(\biu/paddress [68]),
    .i1(\biu/bus_unit/mmu/va_vpn [1]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [4]));
  AL_MUX \biu/bus_unit/mmu/mux29_b40  (
    .i0(\biu/paddress [104]),
    .i1(\biu/bus_unit/mmu_hwdata [38]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [40]));
  AL_MUX \biu/bus_unit/mmu/mux29_b41  (
    .i0(\biu/paddress [105]),
    .i1(\biu/bus_unit/mmu_hwdata [39]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [41]));
  AL_MUX \biu/bus_unit/mmu/mux29_b42  (
    .i0(\biu/paddress [106]),
    .i1(\biu/bus_unit/mmu_hwdata [40]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [42]));
  AL_MUX \biu/bus_unit/mmu/mux29_b43  (
    .i0(\biu/paddress [107]),
    .i1(\biu/bus_unit/mmu_hwdata [41]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [43]));
  AL_MUX \biu/bus_unit/mmu/mux29_b44  (
    .i0(\biu/paddress [108]),
    .i1(\biu/bus_unit/mmu_hwdata [42]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [44]));
  AL_MUX \biu/bus_unit/mmu/mux29_b45  (
    .i0(\biu/paddress [109]),
    .i1(\biu/bus_unit/mmu_hwdata [43]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [45]));
  AL_MUX \biu/bus_unit/mmu/mux29_b46  (
    .i0(\biu/paddress [110]),
    .i1(\biu/bus_unit/mmu_hwdata [44]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [46]));
  AL_MUX \biu/bus_unit/mmu/mux29_b47  (
    .i0(\biu/paddress [111]),
    .i1(\biu/bus_unit/mmu_hwdata [45]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [47]));
  AL_MUX \biu/bus_unit/mmu/mux29_b48  (
    .i0(\biu/paddress [112]),
    .i1(\biu/bus_unit/mmu_hwdata [46]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [48]));
  AL_MUX \biu/bus_unit/mmu/mux29_b49  (
    .i0(\biu/paddress [113]),
    .i1(\biu/bus_unit/mmu_hwdata [47]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [49]));
  AL_MUX \biu/bus_unit/mmu/mux29_b5  (
    .i0(\biu/paddress [69]),
    .i1(\biu/bus_unit/mmu/va_vpn [2]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [5]));
  AL_MUX \biu/bus_unit/mmu/mux29_b50  (
    .i0(\biu/paddress [114]),
    .i1(\biu/bus_unit/mmu_hwdata [48]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [50]));
  AL_MUX \biu/bus_unit/mmu/mux29_b51  (
    .i0(\biu/paddress [115]),
    .i1(\biu/bus_unit/mmu_hwdata [49]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [51]));
  AL_MUX \biu/bus_unit/mmu/mux29_b52  (
    .i0(\biu/paddress [116]),
    .i1(\biu/bus_unit/mmu_hwdata [50]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [52]));
  AL_MUX \biu/bus_unit/mmu/mux29_b53  (
    .i0(\biu/paddress [117]),
    .i1(\biu/bus_unit/mmu_hwdata [51]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [53]));
  AL_MUX \biu/bus_unit/mmu/mux29_b54  (
    .i0(\biu/paddress [118]),
    .i1(\biu/bus_unit/mmu_hwdata [52]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [54]));
  AL_MUX \biu/bus_unit/mmu/mux29_b55  (
    .i0(\biu/paddress [119]),
    .i1(\biu/bus_unit/mmu_hwdata [53]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [55]));
  AL_MUX \biu/bus_unit/mmu/mux29_b56  (
    .i0(\biu/paddress [120]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [56]));
  AL_MUX \biu/bus_unit/mmu/mux29_b57  (
    .i0(\biu/paddress [121]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [57]));
  AL_MUX \biu/bus_unit/mmu/mux29_b58  (
    .i0(\biu/paddress [122]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [58]));
  AL_MUX \biu/bus_unit/mmu/mux29_b59  (
    .i0(\biu/paddress [123]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [59]));
  AL_MUX \biu/bus_unit/mmu/mux29_b6  (
    .i0(\biu/paddress [70]),
    .i1(\biu/bus_unit/mmu/va_vpn [3]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [6]));
  AL_MUX \biu/bus_unit/mmu/mux29_b60  (
    .i0(\biu/paddress [124]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [60]));
  AL_MUX \biu/bus_unit/mmu/mux29_b61  (
    .i0(\biu/paddress [125]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [61]));
  AL_MUX \biu/bus_unit/mmu/mux29_b62  (
    .i0(\biu/paddress [126]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [62]));
  AL_MUX \biu/bus_unit/mmu/mux29_b63  (
    .i0(\biu/paddress [127]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [63]));
  AL_MUX \biu/bus_unit/mmu/mux29_b7  (
    .i0(\biu/paddress [71]),
    .i1(\biu/bus_unit/mmu/va_vpn [4]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [7]));
  AL_MUX \biu/bus_unit/mmu/mux29_b8  (
    .i0(\biu/paddress [72]),
    .i1(\biu/bus_unit/mmu/va_vpn [5]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [8]));
  AL_MUX \biu/bus_unit/mmu/mux29_b9  (
    .i0(\biu/paddress [73]),
    .i1(\biu/bus_unit/mmu/va_vpn [6]),
    .sel(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n70 [9]));
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux2_b0  (
    .i0(\biu/bus_unit/mmu/n29 [0]),
    .i1(\biu/maddress [12]),
    .sel(\biu/bus_unit/mmu/n26 ),
    .o(\biu/bus_unit/mmu/va_vpn [0]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux2_b1  (
    .i0(\biu/bus_unit/mmu/n29 [1]),
    .i1(\biu/maddress [13]),
    .sel(\biu/bus_unit/mmu/n26 ),
    .o(\biu/bus_unit/mmu/va_vpn [1]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux2_b2  (
    .i0(\biu/bus_unit/mmu/n29 [2]),
    .i1(\biu/maddress [14]),
    .sel(\biu/bus_unit/mmu/n26 ),
    .o(\biu/bus_unit/mmu/va_vpn [2]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux2_b3  (
    .i0(\biu/bus_unit/mmu/n29 [3]),
    .i1(\biu/maddress [15]),
    .sel(\biu/bus_unit/mmu/n26 ),
    .o(\biu/bus_unit/mmu/va_vpn [3]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux2_b4  (
    .i0(\biu/bus_unit/mmu/n29 [4]),
    .i1(\biu/maddress [16]),
    .sel(\biu/bus_unit/mmu/n26 ),
    .o(\biu/bus_unit/mmu/va_vpn [4]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux2_b5  (
    .i0(\biu/bus_unit/mmu/n29 [5]),
    .i1(\biu/maddress [17]),
    .sel(\biu/bus_unit/mmu/n26 ),
    .o(\biu/bus_unit/mmu/va_vpn [5]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux2_b6  (
    .i0(\biu/bus_unit/mmu/n29 [6]),
    .i1(\biu/maddress [18]),
    .sel(\biu/bus_unit/mmu/n26 ),
    .o(\biu/bus_unit/mmu/va_vpn [6]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux2_b7  (
    .i0(\biu/bus_unit/mmu/n29 [7]),
    .i1(\biu/maddress [19]),
    .sel(\biu/bus_unit/mmu/n26 ),
    .o(\biu/bus_unit/mmu/va_vpn [7]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux2_b8  (
    .i0(\biu/bus_unit/mmu/n29 [8]),
    .i1(\biu/maddress [20]),
    .sel(\biu/bus_unit/mmu/n26 ),
    .o(\biu/bus_unit/mmu/va_vpn [8]));  // ../../RTL/CPU/BIU/mmu.v(115)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b0  (
    .i0(\biu/bus_unit/mmu/n70 [0]),
    .i1(\biu/bus_unit/mmu/n68 [0]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [0]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b1  (
    .i0(\biu/bus_unit/mmu/n70 [1]),
    .i1(\biu/bus_unit/mmu/n68 [1]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [1]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b10  (
    .i0(\biu/bus_unit/mmu/n70 [10]),
    .i1(\biu/bus_unit/mmu/n68 [10]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [10]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b11  (
    .i0(\biu/bus_unit/mmu/n70 [11]),
    .i1(\biu/bus_unit/mmu/n68 [11]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [11]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b12  (
    .i0(\biu/bus_unit/mmu/n70 [12]),
    .i1(\biu/bus_unit/mmu/n68 [12]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [12]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b13  (
    .i0(\biu/bus_unit/mmu/n70 [13]),
    .i1(\biu/bus_unit/mmu/n68 [13]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [13]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b14  (
    .i0(\biu/bus_unit/mmu/n70 [14]),
    .i1(\biu/bus_unit/mmu/n68 [14]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [14]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b15  (
    .i0(\biu/bus_unit/mmu/n70 [15]),
    .i1(\biu/bus_unit/mmu/n68 [15]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [15]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b16  (
    .i0(\biu/bus_unit/mmu/n70 [16]),
    .i1(\biu/bus_unit/mmu/n68 [16]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [16]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b17  (
    .i0(\biu/bus_unit/mmu/n70 [17]),
    .i1(\biu/bus_unit/mmu/n68 [17]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [17]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b18  (
    .i0(\biu/bus_unit/mmu/n70 [18]),
    .i1(\biu/bus_unit/mmu/n68 [18]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [18]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b19  (
    .i0(\biu/bus_unit/mmu/n70 [19]),
    .i1(\biu/bus_unit/mmu/n68 [19]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [19]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b2  (
    .i0(\biu/bus_unit/mmu/n70 [2]),
    .i1(\biu/bus_unit/mmu/n68 [2]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [2]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b20  (
    .i0(\biu/bus_unit/mmu/n70 [20]),
    .i1(\biu/bus_unit/mmu/n68 [20]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [20]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b21  (
    .i0(\biu/bus_unit/mmu/n70 [21]),
    .i1(\biu/bus_unit/mmu/n68 [21]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [21]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b22  (
    .i0(\biu/bus_unit/mmu/n70 [22]),
    .i1(\biu/bus_unit/mmu/n68 [22]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [22]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b23  (
    .i0(\biu/bus_unit/mmu/n70 [23]),
    .i1(\biu/bus_unit/mmu/n68 [23]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [23]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b24  (
    .i0(\biu/bus_unit/mmu/n70 [24]),
    .i1(\biu/bus_unit/mmu/n68 [24]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [24]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b25  (
    .i0(\biu/bus_unit/mmu/n70 [25]),
    .i1(\biu/bus_unit/mmu/n68 [25]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [25]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b26  (
    .i0(\biu/bus_unit/mmu/n70 [26]),
    .i1(\biu/bus_unit/mmu/n68 [26]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [26]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b27  (
    .i0(\biu/bus_unit/mmu/n70 [27]),
    .i1(\biu/bus_unit/mmu/n68 [27]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [27]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b28  (
    .i0(\biu/bus_unit/mmu/n70 [28]),
    .i1(\biu/bus_unit/mmu/n68 [28]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [28]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b29  (
    .i0(\biu/bus_unit/mmu/n70 [29]),
    .i1(\biu/bus_unit/mmu/n68 [29]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [29]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b3  (
    .i0(\biu/bus_unit/mmu/n70 [3]),
    .i1(\biu/bus_unit/mmu/n68 [3]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [3]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b30  (
    .i0(\biu/bus_unit/mmu/n70 [30]),
    .i1(\biu/bus_unit/mmu/n68 [30]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [30]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b31  (
    .i0(\biu/bus_unit/mmu/n70 [31]),
    .i1(\biu/bus_unit/mmu/n68 [31]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [31]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b32  (
    .i0(\biu/bus_unit/mmu/n70 [32]),
    .i1(\biu/bus_unit/mmu/n68 [32]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [32]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b33  (
    .i0(\biu/bus_unit/mmu/n70 [33]),
    .i1(\biu/bus_unit/mmu/n68 [33]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [33]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b34  (
    .i0(\biu/bus_unit/mmu/n70 [34]),
    .i1(\biu/bus_unit/mmu/n68 [34]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [34]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b35  (
    .i0(\biu/bus_unit/mmu/n70 [35]),
    .i1(\biu/bus_unit/mmu/n68 [35]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [35]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b36  (
    .i0(\biu/bus_unit/mmu/n70 [36]),
    .i1(\biu/bus_unit/mmu/n68 [36]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [36]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b37  (
    .i0(\biu/bus_unit/mmu/n70 [37]),
    .i1(\biu/bus_unit/mmu/n68 [37]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [37]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b38  (
    .i0(\biu/bus_unit/mmu/n70 [38]),
    .i1(\biu/bus_unit/mmu/n68 [38]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [38]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b39  (
    .i0(\biu/bus_unit/mmu/n70 [39]),
    .i1(\biu/bus_unit/mmu/n68 [39]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [39]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b4  (
    .i0(\biu/bus_unit/mmu/n70 [4]),
    .i1(\biu/bus_unit/mmu/n68 [4]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [4]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b40  (
    .i0(\biu/bus_unit/mmu/n70 [40]),
    .i1(\biu/bus_unit/mmu/n68 [40]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [40]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b41  (
    .i0(\biu/bus_unit/mmu/n70 [41]),
    .i1(\biu/bus_unit/mmu/n68 [41]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [41]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b42  (
    .i0(\biu/bus_unit/mmu/n70 [42]),
    .i1(\biu/bus_unit/mmu/n68 [42]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [42]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b43  (
    .i0(\biu/bus_unit/mmu/n70 [43]),
    .i1(\biu/bus_unit/mmu/n68 [43]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [43]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b44  (
    .i0(\biu/bus_unit/mmu/n70 [44]),
    .i1(\biu/bus_unit/mmu/n68 [44]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [44]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b45  (
    .i0(\biu/bus_unit/mmu/n70 [45]),
    .i1(\biu/bus_unit/mmu/n68 [45]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [45]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b46  (
    .i0(\biu/bus_unit/mmu/n70 [46]),
    .i1(\biu/bus_unit/mmu/n68 [46]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [46]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b47  (
    .i0(\biu/bus_unit/mmu/n70 [47]),
    .i1(\biu/bus_unit/mmu/n68 [47]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [47]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b48  (
    .i0(\biu/bus_unit/mmu/n70 [48]),
    .i1(\biu/bus_unit/mmu/n68 [48]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [48]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b49  (
    .i0(\biu/bus_unit/mmu/n70 [49]),
    .i1(\biu/bus_unit/mmu/n68 [49]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [49]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b5  (
    .i0(\biu/bus_unit/mmu/n70 [5]),
    .i1(\biu/bus_unit/mmu/n68 [5]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [5]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b50  (
    .i0(\biu/bus_unit/mmu/n70 [50]),
    .i1(\biu/bus_unit/mmu/n68 [50]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [50]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b51  (
    .i0(\biu/bus_unit/mmu/n70 [51]),
    .i1(\biu/bus_unit/mmu/n68 [51]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [51]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b52  (
    .i0(\biu/bus_unit/mmu/n70 [52]),
    .i1(\biu/bus_unit/mmu/n68 [52]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [52]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b53  (
    .i0(\biu/bus_unit/mmu/n70 [53]),
    .i1(\biu/bus_unit/mmu/n68 [53]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [53]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b54  (
    .i0(\biu/bus_unit/mmu/n70 [54]),
    .i1(\biu/bus_unit/mmu/n68 [54]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [54]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b55  (
    .i0(\biu/bus_unit/mmu/n70 [55]),
    .i1(\biu/bus_unit/mmu/n68 [55]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [55]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b56  (
    .i0(\biu/bus_unit/mmu/n70 [56]),
    .i1(\biu/bus_unit/mmu/n68 [56]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [56]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b57  (
    .i0(\biu/bus_unit/mmu/n70 [57]),
    .i1(\biu/bus_unit/mmu/n68 [57]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [57]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b58  (
    .i0(\biu/bus_unit/mmu/n70 [58]),
    .i1(\biu/bus_unit/mmu/n68 [58]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [58]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b59  (
    .i0(\biu/bus_unit/mmu/n70 [59]),
    .i1(\biu/bus_unit/mmu/n68 [59]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [59]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b6  (
    .i0(\biu/bus_unit/mmu/n70 [6]),
    .i1(\biu/bus_unit/mmu/n68 [6]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [6]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b60  (
    .i0(\biu/bus_unit/mmu/n70 [60]),
    .i1(\biu/bus_unit/mmu/n68 [60]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [60]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b61  (
    .i0(\biu/bus_unit/mmu/n70 [61]),
    .i1(\biu/bus_unit/mmu/n68 [61]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [61]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b62  (
    .i0(\biu/bus_unit/mmu/n70 [62]),
    .i1(\biu/bus_unit/mmu/n68 [62]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [62]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b63  (
    .i0(\biu/bus_unit/mmu/n70 [63]),
    .i1(\biu/bus_unit/mmu/n68 [63]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [63]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b7  (
    .i0(\biu/bus_unit/mmu/n70 [7]),
    .i1(\biu/bus_unit/mmu/n68 [7]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [7]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b8  (
    .i0(\biu/bus_unit/mmu/n70 [8]),
    .i1(\biu/bus_unit/mmu/n68 [8]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [8]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux30_b9  (
    .i0(\biu/bus_unit/mmu/n70 [9]),
    .i1(\biu/bus_unit/mmu/n68 [9]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n71 [9]));  // ../../RTL/CPU/BIU/mmu.v(198)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b0  (
    .i0(\biu/bus_unit/mmu_hwdata [0]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [0]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b1  (
    .i0(\biu/bus_unit/mmu_hwdata [1]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [1]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b10  (
    .i0(\biu/bus_unit/mmu_hwdata [10]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [10]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b11  (
    .i0(\biu/bus_unit/mmu_hwdata [11]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [11]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b12  (
    .i0(\biu/bus_unit/mmu_hwdata [12]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [12]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b13  (
    .i0(\biu/bus_unit/mmu_hwdata [13]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [13]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b14  (
    .i0(\biu/bus_unit/mmu_hwdata [14]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [14]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b15  (
    .i0(\biu/bus_unit/mmu_hwdata [15]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [15]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b16  (
    .i0(\biu/bus_unit/mmu_hwdata [16]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [16]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b17  (
    .i0(\biu/bus_unit/mmu_hwdata [17]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [17]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b18  (
    .i0(\biu/bus_unit/mmu_hwdata [18]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [18]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b19  (
    .i0(\biu/bus_unit/mmu_hwdata [19]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [19]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b2  (
    .i0(\biu/bus_unit/mmu_hwdata [2]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [2]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b20  (
    .i0(\biu/bus_unit/mmu_hwdata [20]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [20]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b21  (
    .i0(\biu/bus_unit/mmu_hwdata [21]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [21]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b22  (
    .i0(\biu/bus_unit/mmu_hwdata [22]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [22]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b23  (
    .i0(\biu/bus_unit/mmu_hwdata [23]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [23]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b24  (
    .i0(\biu/bus_unit/mmu_hwdata [24]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [24]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b25  (
    .i0(\biu/bus_unit/mmu_hwdata [25]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [25]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b26  (
    .i0(\biu/bus_unit/mmu_hwdata [26]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [26]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b27  (
    .i0(\biu/bus_unit/mmu_hwdata [27]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [27]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b28  (
    .i0(\biu/bus_unit/mmu_hwdata [28]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [28]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b29  (
    .i0(\biu/bus_unit/mmu_hwdata [29]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [29]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b3  (
    .i0(\biu/bus_unit/mmu_hwdata [3]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [3]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b30  (
    .i0(\biu/bus_unit/mmu_hwdata [30]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [30]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b31  (
    .i0(\biu/bus_unit/mmu_hwdata [31]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [31]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b32  (
    .i0(\biu/bus_unit/mmu_hwdata [32]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [32]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b33  (
    .i0(\biu/bus_unit/mmu_hwdata [33]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [33]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b34  (
    .i0(\biu/bus_unit/mmu_hwdata [34]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [34]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b35  (
    .i0(\biu/bus_unit/mmu_hwdata [35]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [35]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b36  (
    .i0(\biu/bus_unit/mmu_hwdata [36]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [36]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b37  (
    .i0(\biu/bus_unit/mmu_hwdata [37]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [37]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b38  (
    .i0(\biu/bus_unit/mmu_hwdata [38]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [38]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b39  (
    .i0(\biu/bus_unit/mmu_hwdata [39]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [39]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b4  (
    .i0(\biu/bus_unit/mmu_hwdata [4]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [4]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b40  (
    .i0(\biu/bus_unit/mmu_hwdata [40]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [40]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b41  (
    .i0(\biu/bus_unit/mmu_hwdata [41]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [41]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b42  (
    .i0(\biu/bus_unit/mmu_hwdata [42]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [42]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b43  (
    .i0(\biu/bus_unit/mmu_hwdata [43]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [43]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b44  (
    .i0(\biu/bus_unit/mmu_hwdata [44]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [44]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b45  (
    .i0(\biu/bus_unit/mmu_hwdata [45]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [45]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b46  (
    .i0(\biu/bus_unit/mmu_hwdata [46]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [46]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b47  (
    .i0(\biu/bus_unit/mmu_hwdata [47]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [47]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b48  (
    .i0(\biu/bus_unit/mmu_hwdata [48]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [48]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b49  (
    .i0(\biu/bus_unit/mmu_hwdata [49]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [49]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b5  (
    .i0(\biu/bus_unit/mmu_hwdata [5]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [5]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b50  (
    .i0(\biu/bus_unit/mmu_hwdata [50]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [50]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b51  (
    .i0(\biu/bus_unit/mmu_hwdata [51]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [51]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b52  (
    .i0(\biu/bus_unit/mmu_hwdata [52]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [52]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b53  (
    .i0(\biu/bus_unit/mmu_hwdata [53]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [53]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b54  (
    .i0(\biu/bus_unit/mmu_hwdata [54]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [54]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b55  (
    .i0(\biu/bus_unit/mmu_hwdata [55]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [55]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b56  (
    .i0(\biu/bus_unit/mmu_hwdata [56]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [56]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b57  (
    .i0(\biu/bus_unit/mmu_hwdata [57]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [57]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b58  (
    .i0(\biu/bus_unit/mmu_hwdata [58]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [58]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b59  (
    .i0(\biu/bus_unit/mmu_hwdata [59]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [59]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b6  (
    .i0(\biu/bus_unit/mmu_hwdata [6]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [6]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b60  (
    .i0(\biu/bus_unit/mmu_hwdata [60]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [60]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b61  (
    .i0(\biu/bus_unit/mmu_hwdata [61]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [61]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b62  (
    .i0(\biu/bus_unit/mmu_hwdata [62]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [62]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b63  (
    .i0(\biu/bus_unit/mmu_hwdata [63]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [63]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b7  (
    .i0(\biu/bus_unit/mmu_hwdata [7]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [7]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b8  (
    .i0(\biu/bus_unit/mmu_hwdata [8]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [8]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux32_b9  (
    .i0(\biu/bus_unit/mmu_hwdata [9]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n74 ),
    .o(\biu/bus_unit/mmu/n75 [9]));  // ../../RTL/CPU/BIU/mmu.v(209)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux33_b6  (
    .i0(\biu/bus_unit/mmu_hwdata [6]),
    .i1(hrdata[6]),
    .sel(hready),
    .o(\biu/bus_unit/mmu/n76 [6]));  // ../../RTL/CPU/BIU/mmu.v(212)
  AL_MUX \biu/bus_unit/mmu/mux34_b0  (
    .i0(\biu/bus_unit/mmu_hwdata [0]),
    .i1(hrdata[0]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [0]));
  and \biu/bus_unit/mmu/mux34_b0_sel_is_3  (\biu/bus_unit/mmu/mux34_b0_sel_is_3_o , \biu/bus_unit/mmu/n35 , hready);
  AL_MUX \biu/bus_unit/mmu/mux34_b1  (
    .i0(\biu/bus_unit/mmu_hwdata [1]),
    .i1(hrdata[1]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [1]));
  AL_MUX \biu/bus_unit/mmu/mux34_b10  (
    .i0(\biu/bus_unit/mmu_hwdata [10]),
    .i1(hrdata[10]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [10]));
  AL_MUX \biu/bus_unit/mmu/mux34_b11  (
    .i0(\biu/bus_unit/mmu_hwdata [11]),
    .i1(hrdata[11]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [11]));
  AL_MUX \biu/bus_unit/mmu/mux34_b12  (
    .i0(\biu/bus_unit/mmu_hwdata [12]),
    .i1(hrdata[12]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [12]));
  AL_MUX \biu/bus_unit/mmu/mux34_b13  (
    .i0(\biu/bus_unit/mmu_hwdata [13]),
    .i1(hrdata[13]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [13]));
  AL_MUX \biu/bus_unit/mmu/mux34_b14  (
    .i0(\biu/bus_unit/mmu_hwdata [14]),
    .i1(hrdata[14]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [14]));
  AL_MUX \biu/bus_unit/mmu/mux34_b15  (
    .i0(\biu/bus_unit/mmu_hwdata [15]),
    .i1(hrdata[15]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [15]));
  AL_MUX \biu/bus_unit/mmu/mux34_b16  (
    .i0(\biu/bus_unit/mmu_hwdata [16]),
    .i1(hrdata[16]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [16]));
  AL_MUX \biu/bus_unit/mmu/mux34_b17  (
    .i0(\biu/bus_unit/mmu_hwdata [17]),
    .i1(hrdata[17]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [17]));
  AL_MUX \biu/bus_unit/mmu/mux34_b18  (
    .i0(\biu/bus_unit/mmu_hwdata [18]),
    .i1(hrdata[18]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [18]));
  AL_MUX \biu/bus_unit/mmu/mux34_b19  (
    .i0(\biu/bus_unit/mmu_hwdata [19]),
    .i1(hrdata[19]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [19]));
  AL_MUX \biu/bus_unit/mmu/mux34_b2  (
    .i0(\biu/bus_unit/mmu_hwdata [2]),
    .i1(hrdata[2]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [2]));
  AL_MUX \biu/bus_unit/mmu/mux34_b20  (
    .i0(\biu/bus_unit/mmu_hwdata [20]),
    .i1(hrdata[20]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [20]));
  AL_MUX \biu/bus_unit/mmu/mux34_b21  (
    .i0(\biu/bus_unit/mmu_hwdata [21]),
    .i1(hrdata[21]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [21]));
  AL_MUX \biu/bus_unit/mmu/mux34_b22  (
    .i0(\biu/bus_unit/mmu_hwdata [22]),
    .i1(hrdata[22]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [22]));
  AL_MUX \biu/bus_unit/mmu/mux34_b23  (
    .i0(\biu/bus_unit/mmu_hwdata [23]),
    .i1(hrdata[23]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [23]));
  AL_MUX \biu/bus_unit/mmu/mux34_b24  (
    .i0(\biu/bus_unit/mmu_hwdata [24]),
    .i1(hrdata[24]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [24]));
  AL_MUX \biu/bus_unit/mmu/mux34_b25  (
    .i0(\biu/bus_unit/mmu_hwdata [25]),
    .i1(hrdata[25]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [25]));
  AL_MUX \biu/bus_unit/mmu/mux34_b26  (
    .i0(\biu/bus_unit/mmu_hwdata [26]),
    .i1(hrdata[26]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [26]));
  AL_MUX \biu/bus_unit/mmu/mux34_b27  (
    .i0(\biu/bus_unit/mmu_hwdata [27]),
    .i1(hrdata[27]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [27]));
  AL_MUX \biu/bus_unit/mmu/mux34_b28  (
    .i0(\biu/bus_unit/mmu_hwdata [28]),
    .i1(hrdata[28]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [28]));
  AL_MUX \biu/bus_unit/mmu/mux34_b29  (
    .i0(\biu/bus_unit/mmu_hwdata [29]),
    .i1(hrdata[29]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [29]));
  AL_MUX \biu/bus_unit/mmu/mux34_b3  (
    .i0(\biu/bus_unit/mmu_hwdata [3]),
    .i1(hrdata[3]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [3]));
  AL_MUX \biu/bus_unit/mmu/mux34_b30  (
    .i0(\biu/bus_unit/mmu_hwdata [30]),
    .i1(hrdata[30]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [30]));
  AL_MUX \biu/bus_unit/mmu/mux34_b31  (
    .i0(\biu/bus_unit/mmu_hwdata [31]),
    .i1(hrdata[31]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [31]));
  AL_MUX \biu/bus_unit/mmu/mux34_b32  (
    .i0(\biu/bus_unit/mmu_hwdata [32]),
    .i1(hrdata[32]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [32]));
  AL_MUX \biu/bus_unit/mmu/mux34_b33  (
    .i0(\biu/bus_unit/mmu_hwdata [33]),
    .i1(hrdata[33]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [33]));
  AL_MUX \biu/bus_unit/mmu/mux34_b34  (
    .i0(\biu/bus_unit/mmu_hwdata [34]),
    .i1(hrdata[34]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [34]));
  AL_MUX \biu/bus_unit/mmu/mux34_b35  (
    .i0(\biu/bus_unit/mmu_hwdata [35]),
    .i1(hrdata[35]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [35]));
  AL_MUX \biu/bus_unit/mmu/mux34_b36  (
    .i0(\biu/bus_unit/mmu_hwdata [36]),
    .i1(hrdata[36]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [36]));
  AL_MUX \biu/bus_unit/mmu/mux34_b37  (
    .i0(\biu/bus_unit/mmu_hwdata [37]),
    .i1(hrdata[37]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [37]));
  AL_MUX \biu/bus_unit/mmu/mux34_b38  (
    .i0(\biu/bus_unit/mmu_hwdata [38]),
    .i1(hrdata[38]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [38]));
  AL_MUX \biu/bus_unit/mmu/mux34_b39  (
    .i0(\biu/bus_unit/mmu_hwdata [39]),
    .i1(hrdata[39]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [39]));
  AL_MUX \biu/bus_unit/mmu/mux34_b4  (
    .i0(\biu/bus_unit/mmu_hwdata [4]),
    .i1(hrdata[4]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [4]));
  AL_MUX \biu/bus_unit/mmu/mux34_b40  (
    .i0(\biu/bus_unit/mmu_hwdata [40]),
    .i1(hrdata[40]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [40]));
  AL_MUX \biu/bus_unit/mmu/mux34_b41  (
    .i0(\biu/bus_unit/mmu_hwdata [41]),
    .i1(hrdata[41]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [41]));
  AL_MUX \biu/bus_unit/mmu/mux34_b42  (
    .i0(\biu/bus_unit/mmu_hwdata [42]),
    .i1(hrdata[42]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [42]));
  AL_MUX \biu/bus_unit/mmu/mux34_b43  (
    .i0(\biu/bus_unit/mmu_hwdata [43]),
    .i1(hrdata[43]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [43]));
  AL_MUX \biu/bus_unit/mmu/mux34_b44  (
    .i0(\biu/bus_unit/mmu_hwdata [44]),
    .i1(hrdata[44]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [44]));
  AL_MUX \biu/bus_unit/mmu/mux34_b45  (
    .i0(\biu/bus_unit/mmu_hwdata [45]),
    .i1(hrdata[45]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [45]));
  AL_MUX \biu/bus_unit/mmu/mux34_b46  (
    .i0(\biu/bus_unit/mmu_hwdata [46]),
    .i1(hrdata[46]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [46]));
  AL_MUX \biu/bus_unit/mmu/mux34_b47  (
    .i0(\biu/bus_unit/mmu_hwdata [47]),
    .i1(hrdata[47]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [47]));
  AL_MUX \biu/bus_unit/mmu/mux34_b48  (
    .i0(\biu/bus_unit/mmu_hwdata [48]),
    .i1(hrdata[48]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [48]));
  AL_MUX \biu/bus_unit/mmu/mux34_b49  (
    .i0(\biu/bus_unit/mmu_hwdata [49]),
    .i1(hrdata[49]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [49]));
  AL_MUX \biu/bus_unit/mmu/mux34_b5  (
    .i0(\biu/bus_unit/mmu_hwdata [5]),
    .i1(hrdata[5]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [5]));
  AL_MUX \biu/bus_unit/mmu/mux34_b50  (
    .i0(\biu/bus_unit/mmu_hwdata [50]),
    .i1(hrdata[50]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [50]));
  AL_MUX \biu/bus_unit/mmu/mux34_b51  (
    .i0(\biu/bus_unit/mmu_hwdata [51]),
    .i1(hrdata[51]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [51]));
  AL_MUX \biu/bus_unit/mmu/mux34_b52  (
    .i0(\biu/bus_unit/mmu_hwdata [52]),
    .i1(hrdata[52]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [52]));
  AL_MUX \biu/bus_unit/mmu/mux34_b53  (
    .i0(\biu/bus_unit/mmu_hwdata [53]),
    .i1(hrdata[53]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [53]));
  AL_MUX \biu/bus_unit/mmu/mux34_b54  (
    .i0(\biu/bus_unit/mmu_hwdata [54]),
    .i1(hrdata[54]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [54]));
  AL_MUX \biu/bus_unit/mmu/mux34_b55  (
    .i0(\biu/bus_unit/mmu_hwdata [55]),
    .i1(hrdata[55]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [55]));
  AL_MUX \biu/bus_unit/mmu/mux34_b56  (
    .i0(\biu/bus_unit/mmu_hwdata [56]),
    .i1(hrdata[56]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [56]));
  AL_MUX \biu/bus_unit/mmu/mux34_b57  (
    .i0(\biu/bus_unit/mmu_hwdata [57]),
    .i1(hrdata[57]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [57]));
  AL_MUX \biu/bus_unit/mmu/mux34_b58  (
    .i0(\biu/bus_unit/mmu_hwdata [58]),
    .i1(hrdata[58]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [58]));
  AL_MUX \biu/bus_unit/mmu/mux34_b59  (
    .i0(\biu/bus_unit/mmu_hwdata [59]),
    .i1(hrdata[59]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [59]));
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux34_b6  (
    .i0(\biu/bus_unit/mmu/n77 ),
    .i1(\biu/bus_unit/mmu/n76 [6]),
    .sel(\biu/bus_unit/mmu/n35 ),
    .o(\biu/bus_unit/mmu/n78 [6]));  // ../../RTL/CPU/BIU/mmu.v(217)
  AL_MUX \biu/bus_unit/mmu/mux34_b60  (
    .i0(\biu/bus_unit/mmu_hwdata [60]),
    .i1(hrdata[60]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [60]));
  AL_MUX \biu/bus_unit/mmu/mux34_b61  (
    .i0(\biu/bus_unit/mmu_hwdata [61]),
    .i1(hrdata[61]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [61]));
  AL_MUX \biu/bus_unit/mmu/mux34_b62  (
    .i0(\biu/bus_unit/mmu_hwdata [62]),
    .i1(hrdata[62]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [62]));
  AL_MUX \biu/bus_unit/mmu/mux34_b63  (
    .i0(\biu/bus_unit/mmu_hwdata [63]),
    .i1(hrdata[63]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [63]));
  AL_MUX \biu/bus_unit/mmu/mux34_b7  (
    .i0(\biu/bus_unit/mmu_hwdata [7]),
    .i1(hrdata[7]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [7]));
  AL_MUX \biu/bus_unit/mmu/mux34_b8  (
    .i0(\biu/bus_unit/mmu_hwdata [8]),
    .i1(hrdata[8]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [8]));
  AL_MUX \biu/bus_unit/mmu/mux34_b9  (
    .i0(\biu/bus_unit/mmu_hwdata [9]),
    .i1(hrdata[9]),
    .sel(\biu/bus_unit/mmu/mux34_b0_sel_is_3_o ),
    .o(\biu/bus_unit/mmu/n78 [9]));
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b0  (
    .i0(\biu/bus_unit/mmu/n78 [0]),
    .i1(\biu/bus_unit/mmu/n75 [0]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [0]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b1  (
    .i0(\biu/bus_unit/mmu/n78 [1]),
    .i1(\biu/bus_unit/mmu/n75 [1]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [1]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b10  (
    .i0(\biu/bus_unit/mmu/n78 [10]),
    .i1(\biu/bus_unit/mmu/n75 [10]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [10]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b11  (
    .i0(\biu/bus_unit/mmu/n78 [11]),
    .i1(\biu/bus_unit/mmu/n75 [11]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [11]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b12  (
    .i0(\biu/bus_unit/mmu/n78 [12]),
    .i1(\biu/bus_unit/mmu/n75 [12]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [12]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b13  (
    .i0(\biu/bus_unit/mmu/n78 [13]),
    .i1(\biu/bus_unit/mmu/n75 [13]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [13]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b14  (
    .i0(\biu/bus_unit/mmu/n78 [14]),
    .i1(\biu/bus_unit/mmu/n75 [14]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [14]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b15  (
    .i0(\biu/bus_unit/mmu/n78 [15]),
    .i1(\biu/bus_unit/mmu/n75 [15]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [15]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b16  (
    .i0(\biu/bus_unit/mmu/n78 [16]),
    .i1(\biu/bus_unit/mmu/n75 [16]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [16]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b17  (
    .i0(\biu/bus_unit/mmu/n78 [17]),
    .i1(\biu/bus_unit/mmu/n75 [17]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [17]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b18  (
    .i0(\biu/bus_unit/mmu/n78 [18]),
    .i1(\biu/bus_unit/mmu/n75 [18]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [18]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b19  (
    .i0(\biu/bus_unit/mmu/n78 [19]),
    .i1(\biu/bus_unit/mmu/n75 [19]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [19]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b2  (
    .i0(\biu/bus_unit/mmu/n78 [2]),
    .i1(\biu/bus_unit/mmu/n75 [2]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [2]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b20  (
    .i0(\biu/bus_unit/mmu/n78 [20]),
    .i1(\biu/bus_unit/mmu/n75 [20]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [20]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b21  (
    .i0(\biu/bus_unit/mmu/n78 [21]),
    .i1(\biu/bus_unit/mmu/n75 [21]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [21]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b22  (
    .i0(\biu/bus_unit/mmu/n78 [22]),
    .i1(\biu/bus_unit/mmu/n75 [22]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [22]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b23  (
    .i0(\biu/bus_unit/mmu/n78 [23]),
    .i1(\biu/bus_unit/mmu/n75 [23]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [23]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b24  (
    .i0(\biu/bus_unit/mmu/n78 [24]),
    .i1(\biu/bus_unit/mmu/n75 [24]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [24]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b25  (
    .i0(\biu/bus_unit/mmu/n78 [25]),
    .i1(\biu/bus_unit/mmu/n75 [25]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [25]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b26  (
    .i0(\biu/bus_unit/mmu/n78 [26]),
    .i1(\biu/bus_unit/mmu/n75 [26]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [26]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b27  (
    .i0(\biu/bus_unit/mmu/n78 [27]),
    .i1(\biu/bus_unit/mmu/n75 [27]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [27]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b28  (
    .i0(\biu/bus_unit/mmu/n78 [28]),
    .i1(\biu/bus_unit/mmu/n75 [28]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [28]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b29  (
    .i0(\biu/bus_unit/mmu/n78 [29]),
    .i1(\biu/bus_unit/mmu/n75 [29]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [29]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b3  (
    .i0(\biu/bus_unit/mmu/n78 [3]),
    .i1(\biu/bus_unit/mmu/n75 [3]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [3]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b30  (
    .i0(\biu/bus_unit/mmu/n78 [30]),
    .i1(\biu/bus_unit/mmu/n75 [30]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [30]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b31  (
    .i0(\biu/bus_unit/mmu/n78 [31]),
    .i1(\biu/bus_unit/mmu/n75 [31]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [31]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b32  (
    .i0(\biu/bus_unit/mmu/n78 [32]),
    .i1(\biu/bus_unit/mmu/n75 [32]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [32]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b33  (
    .i0(\biu/bus_unit/mmu/n78 [33]),
    .i1(\biu/bus_unit/mmu/n75 [33]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [33]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b34  (
    .i0(\biu/bus_unit/mmu/n78 [34]),
    .i1(\biu/bus_unit/mmu/n75 [34]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [34]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b35  (
    .i0(\biu/bus_unit/mmu/n78 [35]),
    .i1(\biu/bus_unit/mmu/n75 [35]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [35]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b36  (
    .i0(\biu/bus_unit/mmu/n78 [36]),
    .i1(\biu/bus_unit/mmu/n75 [36]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [36]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b37  (
    .i0(\biu/bus_unit/mmu/n78 [37]),
    .i1(\biu/bus_unit/mmu/n75 [37]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [37]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b38  (
    .i0(\biu/bus_unit/mmu/n78 [38]),
    .i1(\biu/bus_unit/mmu/n75 [38]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [38]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b39  (
    .i0(\biu/bus_unit/mmu/n78 [39]),
    .i1(\biu/bus_unit/mmu/n75 [39]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [39]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b4  (
    .i0(\biu/bus_unit/mmu/n78 [4]),
    .i1(\biu/bus_unit/mmu/n75 [4]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [4]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b40  (
    .i0(\biu/bus_unit/mmu/n78 [40]),
    .i1(\biu/bus_unit/mmu/n75 [40]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [40]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b41  (
    .i0(\biu/bus_unit/mmu/n78 [41]),
    .i1(\biu/bus_unit/mmu/n75 [41]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [41]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b42  (
    .i0(\biu/bus_unit/mmu/n78 [42]),
    .i1(\biu/bus_unit/mmu/n75 [42]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [42]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b43  (
    .i0(\biu/bus_unit/mmu/n78 [43]),
    .i1(\biu/bus_unit/mmu/n75 [43]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [43]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b44  (
    .i0(\biu/bus_unit/mmu/n78 [44]),
    .i1(\biu/bus_unit/mmu/n75 [44]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [44]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b45  (
    .i0(\biu/bus_unit/mmu/n78 [45]),
    .i1(\biu/bus_unit/mmu/n75 [45]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [45]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b46  (
    .i0(\biu/bus_unit/mmu/n78 [46]),
    .i1(\biu/bus_unit/mmu/n75 [46]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [46]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b47  (
    .i0(\biu/bus_unit/mmu/n78 [47]),
    .i1(\biu/bus_unit/mmu/n75 [47]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [47]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b48  (
    .i0(\biu/bus_unit/mmu/n78 [48]),
    .i1(\biu/bus_unit/mmu/n75 [48]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [48]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b49  (
    .i0(\biu/bus_unit/mmu/n78 [49]),
    .i1(\biu/bus_unit/mmu/n75 [49]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [49]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b5  (
    .i0(\biu/bus_unit/mmu/n78 [5]),
    .i1(\biu/bus_unit/mmu/n75 [5]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [5]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b50  (
    .i0(\biu/bus_unit/mmu/n78 [50]),
    .i1(\biu/bus_unit/mmu/n75 [50]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [50]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b51  (
    .i0(\biu/bus_unit/mmu/n78 [51]),
    .i1(\biu/bus_unit/mmu/n75 [51]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [51]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b52  (
    .i0(\biu/bus_unit/mmu/n78 [52]),
    .i1(\biu/bus_unit/mmu/n75 [52]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [52]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b53  (
    .i0(\biu/bus_unit/mmu/n78 [53]),
    .i1(\biu/bus_unit/mmu/n75 [53]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [53]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b54  (
    .i0(\biu/bus_unit/mmu/n78 [54]),
    .i1(\biu/bus_unit/mmu/n75 [54]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [54]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b55  (
    .i0(\biu/bus_unit/mmu/n78 [55]),
    .i1(\biu/bus_unit/mmu/n75 [55]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [55]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b56  (
    .i0(\biu/bus_unit/mmu/n78 [56]),
    .i1(\biu/bus_unit/mmu/n75 [56]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [56]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b57  (
    .i0(\biu/bus_unit/mmu/n78 [57]),
    .i1(\biu/bus_unit/mmu/n75 [57]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [57]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b58  (
    .i0(\biu/bus_unit/mmu/n78 [58]),
    .i1(\biu/bus_unit/mmu/n75 [58]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [58]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b59  (
    .i0(\biu/bus_unit/mmu/n78 [59]),
    .i1(\biu/bus_unit/mmu/n75 [59]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [59]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b6  (
    .i0(\biu/bus_unit/mmu/n78 [6]),
    .i1(\biu/bus_unit/mmu/n75 [6]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [6]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b60  (
    .i0(\biu/bus_unit/mmu/n78 [60]),
    .i1(\biu/bus_unit/mmu/n75 [60]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [60]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b61  (
    .i0(\biu/bus_unit/mmu/n78 [61]),
    .i1(\biu/bus_unit/mmu/n75 [61]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [61]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b62  (
    .i0(\biu/bus_unit/mmu/n78 [62]),
    .i1(\biu/bus_unit/mmu/n75 [62]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [62]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b63  (
    .i0(\biu/bus_unit/mmu/n78 [63]),
    .i1(\biu/bus_unit/mmu/n75 [63]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [63]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b7  (
    .i0(\biu/bus_unit/mmu/n78 [7]),
    .i1(\biu/bus_unit/mmu/n75 [7]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [7]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b8  (
    .i0(\biu/bus_unit/mmu/n78 [8]),
    .i1(\biu/bus_unit/mmu/n75 [8]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [8]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux35_b9  (
    .i0(\biu/bus_unit/mmu/n78 [9]),
    .i1(\biu/bus_unit/mmu/n75 [9]),
    .sel(\biu/bus_unit/mmu/n30 ),
    .o(\biu/bus_unit/mmu/n79 [9]));  // ../../RTL/CPU/BIU/mmu.v(217)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux3_b0  (
    .i0(\biu/pa_cov ),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n33 [0]));  // ../../RTL/CPU/BIU/mmu.v(125)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux3_b1  (
    .i0(\biu/pa_cov ),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n32 ),
    .o(\biu/bus_unit/mmu/n33 [1]));  // ../../RTL/CPU/BIU/mmu.v(125)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux4_b0  (
    .i0(hready),
    .i1(1'b1),
    .sel(hresp),
    .o(\biu/bus_unit/mmu/n36 [0]));  // ../../RTL/CPU/BIU/mmu.v(131)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux4_b1  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(hresp),
    .o(\biu/bus_unit/mmu/n36 [1]));  // ../../RTL/CPU/BIU/mmu.v(131)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux4_b3  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(hresp),
    .o(\biu/bus_unit/mmu/n36 [3]));  // ../../RTL/CPU/BIU/mmu.v(131)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux5_b0  (
    .i0(\biu/bus_unit/mmu/n38 [0]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/pointer_page ),
    .o(\biu/bus_unit/mmu/n39 [0]));  // ../../RTL/CPU/BIU/mmu.v(134)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux6_b0  (
    .i0(\biu/bus_unit/mmu/n39 [0]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/page_unvalid ),
    .o(\biu/bus_unit/mmu/n40 [0]));  // ../../RTL/CPU/BIU/mmu.v(134)
  AL_MUX \biu/bus_unit/mmu/mux6_b1  (
    .i0(1'b0),
    .i1(\biu/bus_unit/mmu/n38 [0]),
    .sel(\biu/bus_unit/mmu/mux6_b1_sel_is_0_o ),
    .o(\biu/bus_unit/mmu/n40 [1]));
  and \biu/bus_unit/mmu/mux6_b1_sel_is_0  (\biu/bus_unit/mmu/mux6_b1_sel_is_0_o , \biu/bus_unit/mmu/page_unvalid_neg , \biu/bus_unit/mmu/pointer_page_neg );
  AL_MUX \biu/bus_unit/mmu/mux6_b2  (
    .i0(1'b0),
    .i1(\biu/bus_unit/mmu/leaf_page ),
    .sel(\biu/bus_unit/mmu/mux6_b1_sel_is_0_o ),
    .o(\biu/bus_unit/mmu/n40 [2]));
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux6_b3  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/page_unvalid ),
    .o(\biu/bus_unit/mmu/n40 [3]));  // ../../RTL/CPU/BIU/mmu.v(134)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux7_b0  (
    .i0(\biu/bus_unit/mmu/page_chk_ok ),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n42 ),
    .o(\biu/bus_unit/mmu/n44 [0]));  // ../../RTL/CPU/BIU/mmu.v(137)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux7_b1  (
    .i0(\biu/bus_unit/mmu/page_chk_ok ),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n42 ),
    .o(\biu/bus_unit/mmu/n44 [1]));  // ../../RTL/CPU/BIU/mmu.v(137)
  binary_mux_s1_w1 \biu/bus_unit/mmu/mux7_b3  (
    .i0(\biu/bus_unit/mmu/n43 [3]),
    .i1(1'b0),
    .sel(\biu/bus_unit/mmu/n42 ),
    .o(\biu/bus_unit/mmu/n44 [3]));  // ../../RTL/CPU/BIU/mmu.v(137)
  and \biu/bus_unit/mmu/mux9_b0_sel_is_0  (\biu/bus_unit/mmu/mux9_b0_sel_is_0_o , \biu/bus_unit/mmu_page_fault_neg , \biu/bus_unit/mmu_acc_fault_neg );
  not \biu/bus_unit/mmu/n30_inv  (\biu/bus_unit/mmu/n30_neg , \biu/bus_unit/mmu/n30 );
  not \biu/bus_unit/mmu/n34_inv  (\biu/bus_unit/mmu/n34_neg , \biu/bus_unit/mmu/n34 );
  not \biu/bus_unit/mmu/n35_inv  (\biu/bus_unit/mmu/n35_neg , \biu/bus_unit/mmu/n35 );
  ne_w4 \biu/bus_unit/mmu/neq0  (
    .i0(satp[63:60]),
    .i1(4'b1000),
    .o(\biu/bus_unit/mmu/n73 ));  // ../../RTL/CPU/BIU/mmu.v(209)
  not \biu/bus_unit/mmu/page_unvalid_inv  (\biu/bus_unit/mmu/page_unvalid_neg , \biu/bus_unit/mmu/page_unvalid );
  not \biu/bus_unit/mmu/pointer_page_inv  (\biu/bus_unit/mmu/pointer_page_neg , \biu/bus_unit/mmu/pointer_page );
  reg_sr_as_w1 \biu/bus_unit/mmu/reg0_b0  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n59 [0]),
    .en(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/mmu/n58 ),
    .set(1'b0),
    .q(\biu/bus_unit/mmu/i [0]));  // ../../RTL/CPU/BIU/mmu.v(166)
  reg_ar_ss_w1 \biu/bus_unit/mmu/reg0_b1  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n59 [1]),
    .en(\biu/bus_unit/mmu/mux20_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(\biu/bus_unit/mmu/n58 ),
    .q(\biu/bus_unit/mmu/i [1]));  // ../../RTL/CPU/BIU/mmu.v(166)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b0  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [0]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b1  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [1]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b10  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [10]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b11  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [11]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b12  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [12]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b13  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [13]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b14  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [14]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b15  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [15]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b16  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [16]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b17  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [17]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b18  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [18]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b19  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [19]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b2  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [2]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b20  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [20]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b21  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [21]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b22  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [22]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b23  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [23]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b24  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [24]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b25  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [25]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b26  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [26]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b27  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [27]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b28  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [28]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b29  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [29]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b3  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [3]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b30  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [30]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b31  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [31]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b32  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [32]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b33  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [33]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b34  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [34]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b35  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [35]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b36  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [36]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b37  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [37]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b38  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [38]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b39  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [39]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b4  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [4]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b40  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [40]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b41  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [41]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b42  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [42]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b43  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [43]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b44  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [44]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b45  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [45]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b46  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [46]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b47  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [47]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b48  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [48]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b49  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [49]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b5  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [5]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b50  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [50]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b51  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [51]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b52  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [52]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b53  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [53]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b54  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [54]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b55  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [55]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b56  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [56]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b57  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [57]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b58  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [58]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b59  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [59]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b6  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [6]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b60  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [60]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b61  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [61]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b62  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [62]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b63  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [63]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b7  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [7]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b8  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [8]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg1_b9  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n66 [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [9]));  // ../../RTL/CPU/BIU/mmu.v(183)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b0  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [64]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b1  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [65]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b10  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [74]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b11  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [75]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b12  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [76]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b13  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [77]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b14  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [78]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b15  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [79]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b16  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [80]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b17  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [81]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b18  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [82]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b19  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [83]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b2  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [66]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b20  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [84]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b21  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [85]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b22  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [86]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b23  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [87]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b24  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [88]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b25  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [89]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b26  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [90]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b27  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [91]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b28  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [92]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b29  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [93]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b3  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [67]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b30  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [94]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b31  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [95]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b32  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [96]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b33  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [97]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b34  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [98]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b35  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [99]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b36  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [100]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b37  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [101]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b38  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [102]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b39  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [103]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b4  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [68]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b40  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [104]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b41  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [105]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b42  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [106]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b43  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [107]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b44  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [108]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b45  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [109]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b46  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [110]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b47  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [111]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b48  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [112]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b49  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [113]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b5  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [69]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b50  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [114]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b51  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [115]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b52  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [116]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b53  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [117]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b54  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [118]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b55  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [119]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b56  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [120]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b57  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [121]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b58  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [122]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b59  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [123]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b6  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [70]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b60  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [124]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b61  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [125]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b62  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [126]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b63  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [127]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b7  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [71]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b8  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [72]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg2_b9  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n71 [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/paddress [73]));  // ../../RTL/CPU/BIU/mmu.v(200)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b0  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [0]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b1  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [1]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b10  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [10]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b11  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [11]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b12  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [12]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b13  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [13]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b14  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [14]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b15  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [15]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b16  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [16]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b17  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [17]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b18  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [18]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b19  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [19]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b2  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [2]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b20  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [20]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b21  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [21]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b22  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [22]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b23  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [23]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b24  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [24]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b25  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [25]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b26  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [26]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b27  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [27]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b28  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [28]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b29  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [29]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b3  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [3]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b30  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [30]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b31  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [31]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b32  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [32]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b33  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [33]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b34  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [34]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b35  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [35]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b36  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [36]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b37  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [37]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b38  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [38]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b39  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [39]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b4  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [4]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b40  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [40]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b41  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [41]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b42  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [42]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b43  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [43]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b44  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [44]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b45  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [45]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b46  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [46]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b47  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [47]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b48  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [48]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b49  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [49]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b5  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [5]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b50  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [50]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b51  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [51]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b52  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [52]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b53  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [53]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b54  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [54]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b55  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [55]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b56  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [56]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b57  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [57]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b58  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [58]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b59  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [59]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b6  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [6]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b60  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [60]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b61  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [61]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b62  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [62]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b63  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [63]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b7  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [7]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b8  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [8]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg3_b9  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n79 [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu_hwdata [9]));  // ../../RTL/CPU/BIU/mmu.v(218)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg4_b0  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n56 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu/statu [0]));  // ../../RTL/CPU/BIU/mmu.v(154)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg4_b1  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n56 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu/statu [1]));  // ../../RTL/CPU/BIU/mmu.v(154)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg4_b2  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n56 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/mmu/statu [2]));  // ../../RTL/CPU/BIU/mmu.v(154)
  reg_sr_as_w1 \biu/bus_unit/mmu/reg4_b3  (
    .clk(clk),
    .d(\biu/bus_unit/mmu/n54 [3]),
    .en(1'b1),
    .reset(~\biu/bus_unit/mmu/mux18_b3_sel_is_2_o ),
    .set(1'b0),
    .q(\biu/bus_unit/mmu/statu [3]));  // ../../RTL/CPU/BIU/mmu.v(154)
  add_pu2_mu2_o2 \biu/bus_unit/mmu/sub0  (
    .i0(\biu/bus_unit/mmu/i ),
    .i1(2'b01),
    .o(\biu/bus_unit/mmu/n59 ));  // ../../RTL/CPU/BIU/mmu.v(164)
  not \biu/bus_unit/mmu/u10  (\biu/bus_unit/mmu/n6 , \biu/bus_unit/mmu_hwdata [1]);  // ../../RTL/CPU/BIU/mmu.v(106)
  and \biu/bus_unit/mmu/u11  (\biu/bus_unit/mmu/pointer_page , \biu/bus_unit/mmu/n5 , \biu/bus_unit/mmu/n6 );  // ../../RTL/CPU/BIU/mmu.v(106)
  or \biu/bus_unit/mmu/u12  (\biu/bus_unit/mmu/leaf_page , \biu/bus_unit/mmu_hwdata [1], \biu/bus_unit/mmu_hwdata [3]);  // ../../RTL/CPU/BIU/mmu.v(107)
  and \biu/bus_unit/mmu/u13  (\biu/bus_unit/mmu/n9 , \biu/bus_unit/mmu/n8 , sum);  // ../../RTL/CPU/BIU/mmu.v(110)
  or \biu/bus_unit/mmu/u14  (\biu/bus_unit/mmu/n10 , \biu/bus_unit/mmu/n7 , \biu/bus_unit/mmu/n9 );  // ../../RTL/CPU/BIU/mmu.v(110)
  and \biu/bus_unit/mmu/u15  (\biu/bus_unit/mmu/n11 , \biu/bus_unit/mmu_hwdata [4], \biu/bus_unit/mmu/n10 );  // ../../RTL/CPU/BIU/mmu.v(110)
  and \biu/bus_unit/mmu/u16  (\biu/bus_unit/mmu/n13 , \biu/bus_unit/mmu/n12 , \biu/bus_unit/mmu_hwdata [2]);  // ../../RTL/CPU/BIU/mmu.v(111)
  and \biu/bus_unit/mmu/u17  (\biu/bus_unit/mmu/n15 , mxr, \biu/bus_unit/mmu_hwdata [3]);  // ../../RTL/CPU/BIU/mmu.v(111)
  or \biu/bus_unit/mmu/u18  (\biu/bus_unit/mmu/n16 , \biu/bus_unit/mmu_hwdata [1], \biu/bus_unit/mmu/n15 );  // ../../RTL/CPU/BIU/mmu.v(111)
  and \biu/bus_unit/mmu/u19  (\biu/bus_unit/mmu/n17 , \biu/bus_unit/mmu/n14 , \biu/bus_unit/mmu/n16 );  // ../../RTL/CPU/BIU/mmu.v(111)
  not \biu/bus_unit/mmu/u2  (\biu/bus_unit/mmu/n46 [1], hresp);  // ../../RTL/CPU/BIU/mmu.v(143)
  or \biu/bus_unit/mmu/u20  (\biu/bus_unit/mmu/n18 , \biu/bus_unit/mmu/n13 , \biu/bus_unit/mmu/n17 );  // ../../RTL/CPU/BIU/mmu.v(111)
  and \biu/bus_unit/mmu/u21  (\biu/bus_unit/mmu/n20 , \biu/bus_unit/mmu/n19 , \biu/bus_unit/mmu_hwdata [3]);  // ../../RTL/CPU/BIU/mmu.v(111)
  or \biu/bus_unit/mmu/u22  (\biu/bus_unit/mmu/n21 , \biu/bus_unit/mmu/n18 , \biu/bus_unit/mmu/n20 );  // ../../RTL/CPU/BIU/mmu.v(111)
  and \biu/bus_unit/mmu/u23  (\biu/bus_unit/mmu/n22 , \biu/bus_unit/mmu/n11 , \biu/bus_unit/mmu/n21 );  // ../../RTL/CPU/BIU/mmu.v(111)
  not \biu/bus_unit/mmu/u3  (\biu/bus_unit/mmu/n38 [0], \biu/bus_unit/mmu/leaf_page );  // ../../RTL/CPU/BIU/mmu.v(134)
  and \biu/bus_unit/mmu/u35  (\biu/bus_unit/mmu/n23 , \biu/bus_unit/mmu/n8 , \biu/bus_unit/mmu/n21 );  // ../../RTL/CPU/BIU/mmu.v(112)
  or \biu/bus_unit/mmu/u36  (\biu/bus_unit/mmu/n24 , \biu/bus_unit/mmu/n22 , \biu/bus_unit/mmu/n23 );  // ../../RTL/CPU/BIU/mmu.v(112)
  or \biu/bus_unit/mmu/u37  (\biu/bus_unit/mmu/page_chk_ok , \biu/bus_unit/mmu/n24 , \biu/bus_unit/mmu/n25 );  // ../../RTL/CPU/BIU/mmu.v(113)
  and \biu/bus_unit/mmu/u39  (\biu/bus_unit/mmu/n32 , \biu/pa_cov , \biu/bus_unit/mmu/n31 );  // ../../RTL/CPU/BIU/mmu.v(125)
  not \biu/bus_unit/mmu/u4  (\biu/bus_unit/mmu/n0 , \biu/bus_unit/mmu_hwdata [6]);  // ../../RTL/CPU/BIU/mmu.v(105)
  not \biu/bus_unit/mmu/u41  (\biu/bus_unit/mmu/n43 [3], \biu/bus_unit/mmu/page_chk_ok );  // ../../RTL/CPU/BIU/mmu.v(137)
  and \biu/bus_unit/mmu/u43  (\biu/bus_unit/mmu/n42 , \biu/bus_unit/mmu/page_chk_ok , \biu/bus_unit/mmu/n0 );  // ../../RTL/CPU/BIU/mmu.v(137)
  or \biu/bus_unit/mmu/u47  (\biu/bus_unit/mmu/n58 , rst, \biu/bus_unit/mmu/n30 );  // ../../RTL/CPU/BIU/mmu.v(160)
  and \biu/bus_unit/mmu/u5  (\biu/bus_unit/mmu/n2 , \biu/bus_unit/mmu/pointer_page , \biu/bus_unit/mmu/n1 );  // ../../RTL/CPU/BIU/mmu.v(105)
  and \biu/bus_unit/mmu/u56  (\biu/bus_unit/mmu/n74 , \biu/bus_unit/mmu/n73 , \biu/pa_cov );  // ../../RTL/CPU/BIU/mmu.v(209)
  AL_MUX \biu/bus_unit/mmu/u59  (
    .i0(\biu/bus_unit/mmu_hwdata [6]),
    .i1(1'b1),
    .sel(\biu/bus_unit/mmu/n41 ),
    .o(\biu/bus_unit/mmu/n77 ));  // ../../RTL/CPU/BIU/mmu.v(217)
  or \biu/bus_unit/mmu/u6  (\biu/bus_unit/mmu/page_unvalid , \biu/bus_unit/mmu/n0 , \biu/bus_unit/mmu/n2 );  // ../../RTL/CPU/BIU/mmu.v(105)
  and \biu/bus_unit/mmu/u61  (\biu/cacheable , \biu/bus_unit/mmu_trans_rdy , \biu/bus_unit/mmu/n81 );  // ../../RTL/CPU/BIU/mmu.v(221)
  not \biu/bus_unit/mmu/u7  (\biu/bus_unit/mmu/n3 , \biu/bus_unit/mmu_hwdata [3]);  // ../../RTL/CPU/BIU/mmu.v(106)
  or \biu/bus_unit/mmu/u75  (\biu/bus_unit/mmu_htrans [1], \biu/bus_unit/mmu/n34 , \biu/bus_unit/mmu_hwrite );  // ../../RTL/CPU/BIU/mmu.v(238)
  not \biu/bus_unit/mmu/u8  (\biu/bus_unit/mmu/n4 , \biu/bus_unit/mmu_hwdata [2]);  // ../../RTL/CPU/BIU/mmu.v(106)
  and \biu/bus_unit/mmu/u9  (\biu/bus_unit/mmu/n5 , \biu/bus_unit/mmu/n3 , \biu/bus_unit/mmu/n4 );  // ../../RTL/CPU/BIU/mmu.v(106)
  not \biu/bus_unit/mmu_acc_fault_inv  (\biu/bus_unit/mmu_acc_fault_neg , \biu/bus_unit/mmu_acc_fault );
  not \biu/bus_unit/mmu_page_fault_inv  (\biu/bus_unit/mmu_page_fault_neg , \biu/bus_unit/mmu_page_fault );
  not \biu/bus_unit/mmu_trans_rdy_inv  (\biu/bus_unit/mmu_trans_rdy_neg , \biu/bus_unit/mmu_trans_rdy );
  AL_MUX \biu/bus_unit/mux10_b0  (
    .i0(\biu/bus_unit/n19 [0]),
    .i1(\biu/bus_unit/n26 [0]),
    .sel(\biu/bus_unit/mux10_b0_sel_is_2_o ),
    .o(\biu/bus_unit/n29 [0]));
  and \biu/bus_unit/mux10_b0_sel_is_2  (\biu/bus_unit/mux10_b0_sel_is_2_o , \biu/bus_unit/n18_neg , \biu/bus_unit/mux9_b0_sel_is_0_o );
  binary_mux_s1_w1 \biu/bus_unit/mux10_b1  (
    .i0(\biu/bus_unit/n28 [1]),
    .i1(\biu/bus_unit/n19 [0]),
    .sel(\biu/bus_unit/n18 ),
    .o(\biu/bus_unit/n29 [1]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  AL_MUX \biu/bus_unit/mux10_b3  (
    .i0(\biu/bus_unit/mmu/n36 [3]),
    .i1(\biu/bus_unit/n27 [3]),
    .sel(\biu/bus_unit/mux10_b3_sel_is_0_o ),
    .o(\biu/bus_unit/n29 [3]));
  and \biu/bus_unit/mux10_b3_sel_is_0  (\biu/bus_unit/mux10_b3_sel_is_0_o , \biu/bus_unit/n18_neg , \biu/bus_unit/n20_neg );
  binary_mux_s1_w1 \biu/bus_unit/mux11_b0  (
    .i0(\biu/bus_unit/n29 [0]),
    .i1(\biu/bus_unit/n17 [0]),
    .sel(\biu/bus_unit/n14 ),
    .o(\biu/bus_unit/n30 [0]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux11_b1  (
    .i0(\biu/bus_unit/n29 [1]),
    .i1(1'b1),
    .sel(\biu/bus_unit/n14 ),
    .o(\biu/bus_unit/n30 [1]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  AL_MUX \biu/bus_unit/mux11_b2  (
    .i0(\biu/bus_unit/mmu/n36 [3]),
    .i1(\biu/bus_unit/n28 [2]),
    .sel(\biu/bus_unit/mux11_b2_sel_is_0_o ),
    .o(\biu/bus_unit/n30 [2]));
  and \biu/bus_unit/mux11_b2_sel_is_0  (\biu/bus_unit/mux11_b2_sel_is_0_o , \biu/bus_unit/n14_neg , \biu/bus_unit/n18_neg );
  binary_mux_s1_w1 \biu/bus_unit/mux11_b3  (
    .i0(\biu/bus_unit/n29 [3]),
    .i1(1'b1),
    .sel(\biu/bus_unit/n14 ),
    .o(\biu/bus_unit/n30 [3]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  AL_MUX \biu/bus_unit/mux11_b4  (
    .i0(\biu/bus_unit/mmu/n36 [3]),
    .i1(\biu/bus_unit/n26 [4]),
    .sel(\biu/bus_unit/mux11_b4_sel_is_2_o ),
    .o(\biu/bus_unit/n30 [4]));
  and \biu/bus_unit/mux11_b4_sel_is_2  (\biu/bus_unit/mux11_b4_sel_is_2_o , \biu/bus_unit/n14_neg , \biu/bus_unit/mux10_b0_sel_is_2_o );
  binary_mux_s1_w1 \biu/bus_unit/mux12_b1  (
    .i0(\biu/bus_unit/n30 [1]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n13 ),
    .o(\biu/bus_unit/n31 [1]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux12_b2  (
    .i0(\biu/bus_unit/n30 [2]),
    .i1(1'b1),
    .sel(\biu/bus_unit/n13 ),
    .o(\biu/bus_unit/n31 [2]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  AL_MUX \biu/bus_unit/mux13_b0  (
    .i0(1'b1),
    .i1(\biu/bus_unit/n30 [0]),
    .sel(\biu/bus_unit/mux13_b0_sel_is_0_o ),
    .o(\biu/bus_unit/n32 [0]));
  and \biu/bus_unit/mux13_b0_sel_is_0  (\biu/bus_unit/mux13_b0_sel_is_0_o , \biu/bus_unit/n12_neg , \biu/bus_unit/n13_neg );
  AL_MUX \biu/bus_unit/mux13_b3  (
    .i0(1'b0),
    .i1(\biu/bus_unit/n30 [3]),
    .sel(\biu/bus_unit/mux13_b0_sel_is_0_o ),
    .o(\biu/bus_unit/n32 [3]));
  binary_mux_s1_w1 \biu/bus_unit/mux14_b0  (
    .i0(\biu/bus_unit/n32 [0]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n11 ),
    .o(\biu/bus_unit/n33 [0]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  AL_MUX \biu/bus_unit/mux14_b1  (
    .i0(1'b1),
    .i1(\biu/bus_unit/n31 [1]),
    .sel(\biu/bus_unit/mux14_b1_sel_is_0_o ),
    .o(\biu/bus_unit/n33 [1]));
  and \biu/bus_unit/mux14_b1_sel_is_0  (\biu/bus_unit/mux14_b1_sel_is_0_o , \biu/bus_unit/n11_neg , \biu/bus_unit/n12_neg );
  binary_mux_s1_w1 \biu/bus_unit/mux14_b3  (
    .i0(\biu/bus_unit/n32 [3]),
    .i1(1'b1),
    .sel(\biu/bus_unit/n11 ),
    .o(\biu/bus_unit/n33 [3]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  and \biu/bus_unit/mux14_b4_sel_is_2  (\biu/bus_unit/mux14_b4_sel_is_2_o , \biu/bus_unit/n11_neg , \biu/bus_unit/mux13_b0_sel_is_0_o );
  binary_mux_s1_w1 \biu/bus_unit/mux15_b0  (
    .i0(\biu/bus_unit/n33 [0]),
    .i1(\biu/bus_unit/n10 ),
    .sel(\biu/bus_unit/n7 ),
    .o(\biu/bus_unit/n34 [0]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux15_b1  (
    .i0(\biu/bus_unit/n33 [1]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(\biu/bus_unit/n34 [1]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  AL_MUX \biu/bus_unit/mux15_b2  (
    .i0(1'b0),
    .i1(\biu/bus_unit/n31 [2]),
    .sel(\biu/bus_unit/mux15_b2_sel_is_2_o ),
    .o(\biu/bus_unit/n34 [2]));
  and \biu/bus_unit/mux15_b2_sel_is_2  (\biu/bus_unit/mux15_b2_sel_is_2_o , \biu/bus_unit/n7_neg , \biu/bus_unit/mux14_b1_sel_is_0_o );
  binary_mux_s1_w1 \biu/bus_unit/mux15_b3  (
    .i0(\biu/bus_unit/n33 [3]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(\biu/bus_unit/n34 [3]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  and \biu/bus_unit/mux15_b4_sel_is_2  (\biu/bus_unit/mux15_b4_sel_is_2_o , \biu/bus_unit/n7_neg , \biu/bus_unit/mux14_b4_sel_is_2_o );
  binary_mux_s1_w1 \biu/bus_unit/mux16_b0  (
    .i0(\biu/bus_unit/n34 [0]),
    .i1(\biu/bus_unit/n6 [0]),
    .sel(\biu/bus_unit/n0 ),
    .o(\biu/bus_unit/n35 [0]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux16_b1  (
    .i0(\biu/bus_unit/n34 [1]),
    .i1(\biu/bus_unit/n6 [1]),
    .sel(\biu/bus_unit/n0 ),
    .o(\biu/bus_unit/n35 [1]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux16_b2  (
    .i0(\biu/bus_unit/n34 [2]),
    .i1(\biu/bus_unit/n6 [2]),
    .sel(\biu/bus_unit/n0 ),
    .o(\biu/bus_unit/n35 [2]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux16_b3  (
    .i0(\biu/bus_unit/n34 [3]),
    .i1(\biu/bus_unit/n6 [3]),
    .sel(\biu/bus_unit/n0 ),
    .o(\biu/bus_unit/n35 [3]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  and \biu/bus_unit/mux16_b4_sel_is_2  (\biu/bus_unit/mux16_b4_sel_is_2_o , \biu/bus_unit/n0_neg , \biu/bus_unit/mux15_b4_sel_is_2_o );
  and \biu/bus_unit/mux17_b4_sel_is_2  (\biu/bus_unit/mux17_b4_sel_is_2_o , rst_neg, \biu/bus_unit/mux16_b4_sel_is_2_o );
  and \biu/bus_unit/mux19_b0_sel_is_3  (\biu/bus_unit/mux19_b0_sel_is_3_o , \biu/bus_unit/n38 , hready);
  and \biu/bus_unit/mux1_b1_sel_is_0  (\biu/bus_unit/mux1_b1_sel_is_0_o , \biu/bus_unit/n1_neg , \biu/bus_unit/n2_neg );
  and \biu/bus_unit/mux1_b2_sel_is_2  (\biu/bus_unit/mux1_b2_sel_is_2_o , \biu/bus_unit/n1_neg , \biu/bus_unit/n2 );
  binary_mux_s1_w1 \biu/bus_unit/mux22_b0  (
    .i0(\biu/maddress [0]),
    .i1(\biu/paddress [64]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[0]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b1  (
    .i0(\biu/maddress [1]),
    .i1(\biu/paddress [65]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[1]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b10  (
    .i0(\biu/bus_unit/n49 [7]),
    .i1(\biu/paddress [74]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[10]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b11  (
    .i0(\biu/bus_unit/n49 [8]),
    .i1(\biu/paddress [75]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[11]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b12  (
    .i0(\biu/bus_unit/n49 [9]),
    .i1(\biu/paddress [76]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[12]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b13  (
    .i0(\biu/bus_unit/n49 [10]),
    .i1(\biu/paddress [77]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[13]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b14  (
    .i0(\biu/bus_unit/n49 [11]),
    .i1(\biu/paddress [78]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[14]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b15  (
    .i0(\biu/bus_unit/n49 [12]),
    .i1(\biu/paddress [79]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[15]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b16  (
    .i0(\biu/bus_unit/n49 [13]),
    .i1(\biu/paddress [80]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[16]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b17  (
    .i0(\biu/bus_unit/n49 [14]),
    .i1(\biu/paddress [81]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[17]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b18  (
    .i0(\biu/bus_unit/n49 [15]),
    .i1(\biu/paddress [82]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[18]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b19  (
    .i0(\biu/bus_unit/n49 [16]),
    .i1(\biu/paddress [83]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[19]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b2  (
    .i0(\biu/maddress [2]),
    .i1(\biu/paddress [66]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[2]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b20  (
    .i0(\biu/bus_unit/n49 [17]),
    .i1(\biu/paddress [84]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[20]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b21  (
    .i0(\biu/bus_unit/n49 [18]),
    .i1(\biu/paddress [85]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[21]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b22  (
    .i0(\biu/bus_unit/n49 [19]),
    .i1(\biu/paddress [86]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[22]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b23  (
    .i0(\biu/bus_unit/n49 [20]),
    .i1(\biu/paddress [87]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[23]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b24  (
    .i0(\biu/bus_unit/n49 [21]),
    .i1(\biu/paddress [88]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[24]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b25  (
    .i0(\biu/bus_unit/n49 [22]),
    .i1(\biu/paddress [89]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[25]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b26  (
    .i0(\biu/bus_unit/n49 [23]),
    .i1(\biu/paddress [90]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[26]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b27  (
    .i0(\biu/bus_unit/n49 [24]),
    .i1(\biu/paddress [91]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[27]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b28  (
    .i0(\biu/bus_unit/n49 [25]),
    .i1(\biu/paddress [92]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[28]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b29  (
    .i0(\biu/bus_unit/n49 [26]),
    .i1(\biu/paddress [93]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[29]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b3  (
    .i0(\biu/bus_unit/n49 [0]),
    .i1(\biu/paddress [67]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[3]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b30  (
    .i0(\biu/bus_unit/n49 [27]),
    .i1(\biu/paddress [94]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[30]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b31  (
    .i0(\biu/bus_unit/n49 [28]),
    .i1(\biu/paddress [95]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[31]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b32  (
    .i0(\biu/bus_unit/n49 [29]),
    .i1(\biu/paddress [96]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[32]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b33  (
    .i0(\biu/bus_unit/n49 [30]),
    .i1(\biu/paddress [97]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[33]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b34  (
    .i0(\biu/bus_unit/n49 [31]),
    .i1(\biu/paddress [98]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[34]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b35  (
    .i0(\biu/bus_unit/n49 [32]),
    .i1(\biu/paddress [99]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[35]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b36  (
    .i0(\biu/bus_unit/n49 [33]),
    .i1(\biu/paddress [100]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[36]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b37  (
    .i0(\biu/bus_unit/n49 [34]),
    .i1(\biu/paddress [101]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[37]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b38  (
    .i0(\biu/bus_unit/n49 [35]),
    .i1(\biu/paddress [102]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[38]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b39  (
    .i0(\biu/bus_unit/n49 [36]),
    .i1(\biu/paddress [103]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[39]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b4  (
    .i0(\biu/bus_unit/n49 [1]),
    .i1(\biu/paddress [68]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[4]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b40  (
    .i0(\biu/bus_unit/n49 [37]),
    .i1(\biu/paddress [104]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[40]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b41  (
    .i0(\biu/bus_unit/n49 [38]),
    .i1(\biu/paddress [105]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[41]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b42  (
    .i0(\biu/bus_unit/n49 [39]),
    .i1(\biu/paddress [106]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[42]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b43  (
    .i0(\biu/bus_unit/n49 [40]),
    .i1(\biu/paddress [107]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[43]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b44  (
    .i0(\biu/bus_unit/n49 [41]),
    .i1(\biu/paddress [108]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[44]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b45  (
    .i0(\biu/bus_unit/n49 [42]),
    .i1(\biu/paddress [109]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[45]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b46  (
    .i0(\biu/bus_unit/n49 [43]),
    .i1(\biu/paddress [110]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[46]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b47  (
    .i0(\biu/bus_unit/n49 [44]),
    .i1(\biu/paddress [111]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[47]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b48  (
    .i0(\biu/bus_unit/n49 [45]),
    .i1(\biu/paddress [112]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[48]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b49  (
    .i0(\biu/bus_unit/n49 [46]),
    .i1(\biu/paddress [113]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[49]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b5  (
    .i0(\biu/bus_unit/n49 [2]),
    .i1(\biu/paddress [69]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[5]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b50  (
    .i0(\biu/bus_unit/n49 [47]),
    .i1(\biu/paddress [114]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[50]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b51  (
    .i0(\biu/bus_unit/n49 [48]),
    .i1(\biu/paddress [115]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[51]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b52  (
    .i0(\biu/bus_unit/n49 [49]),
    .i1(\biu/paddress [116]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[52]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b53  (
    .i0(\biu/bus_unit/n49 [50]),
    .i1(\biu/paddress [117]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[53]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b54  (
    .i0(\biu/bus_unit/n49 [51]),
    .i1(\biu/paddress [118]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[54]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b55  (
    .i0(\biu/bus_unit/n49 [52]),
    .i1(\biu/paddress [119]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[55]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b56  (
    .i0(\biu/bus_unit/n49 [53]),
    .i1(\biu/paddress [120]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[56]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b57  (
    .i0(\biu/bus_unit/n49 [54]),
    .i1(\biu/paddress [121]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[57]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b58  (
    .i0(\biu/bus_unit/n49 [55]),
    .i1(\biu/paddress [122]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[58]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b59  (
    .i0(\biu/bus_unit/n49 [56]),
    .i1(\biu/paddress [123]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[59]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b6  (
    .i0(\biu/bus_unit/n49 [3]),
    .i1(\biu/paddress [70]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[6]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b60  (
    .i0(\biu/bus_unit/n49 [57]),
    .i1(\biu/paddress [124]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[60]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b61  (
    .i0(\biu/bus_unit/n49 [58]),
    .i1(\biu/paddress [125]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[61]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b62  (
    .i0(\biu/bus_unit/n49 [59]),
    .i1(\biu/paddress [126]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[62]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b63  (
    .i0(\biu/bus_unit/n49 [60]),
    .i1(\biu/paddress [127]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[63]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b7  (
    .i0(\biu/bus_unit/n49 [4]),
    .i1(\biu/paddress [71]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[7]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b8  (
    .i0(\biu/bus_unit/n49 [5]),
    .i1(\biu/paddress [72]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[8]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux22_b9  (
    .i0(\biu/bus_unit/n49 [6]),
    .i1(\biu/paddress [73]),
    .sel(\biu/bus_unit/n7 ),
    .o(haddr[9]));  // ../../RTL/CPU/BIU/bus_unit.v(189)
  binary_mux_s1_w1 \biu/bus_unit/mux23_b0  (
    .i0(\biu/bus_unit/n53 ),
    .i1(1'b1),
    .sel(\biu/bus_unit/n51 ),
    .o(\biu/bus_unit/n54 [0]));  // ../../RTL/CPU/BIU/bus_unit.v(191)
  binary_mux_s1_w1 \biu/bus_unit/mux24_b0  (
    .i0(\biu/bus_unit/n54 [0]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n50 ),
    .o(\biu/bus_unit/n55 [0]));  // ../../RTL/CPU/BIU/bus_unit.v(191)
  and \biu/bus_unit/mux24_b1_sel_is_0  (\biu/bus_unit/mux24_b1_sel_is_0_o , \biu/bus_unit/n50_neg , \biu/bus_unit/n51_neg );
  not \biu/bus_unit/mux24_b1_sel_is_0_o_inv  (\biu/bus_unit/mux24_b1_sel_is_0_o_neg , \biu/bus_unit/mux24_b1_sel_is_0_o );
  binary_mux_s1_w1 \biu/bus_unit/mux25_b0  (
    .i0(\biu/bus_unit/n55 [0]),
    .i1(1'b1),
    .sel(\biu/bus_unit/n7 ),
    .o(hsize[0]));  // ../../RTL/CPU/BIU/bus_unit.v(191)
  AL_MUX \biu/bus_unit/mux25_b1  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\biu/bus_unit/mux25_b1_sel_is_0_o ),
    .o(hsize[1]));
  and \biu/bus_unit/mux25_b1_sel_is_0  (\biu/bus_unit/mux25_b1_sel_is_0_o , \biu/bus_unit/n7_neg , \biu/bus_unit/mux24_b1_sel_is_0_o_neg );
  AL_MUX \biu/bus_unit/mux26_b0  (
    .i0(1'b0),
    .i1(\biu/bus_unit/n38 ),
    .sel(\biu/bus_unit/mux26_b0_sel_is_0_o ),
    .o(hburst[0]));
  and \biu/bus_unit/mux26_b0_sel_is_0  (\biu/bus_unit/mux26_b0_sel_is_0_o , \biu/bus_unit/n7_neg , \biu/bus_unit/n56_neg );
  binary_mux_s1_w1 \biu/bus_unit/mux27_b1  (
    .i0(\biu/bus_unit/n14 ),
    .i1(1'b1),
    .sel(\biu/bus_unit/n58 ),
    .o(\biu/bus_unit/n59 [1]));  // ../../RTL/CPU/BIU/bus_unit.v(195)
  AL_MUX \biu/bus_unit/mux28_b0  (
    .i0(1'b0),
    .i1(\biu/bus_unit/n14 ),
    .sel(\biu/bus_unit/mux28_b0_sel_is_0_o ),
    .o(htrans[0]));
  and \biu/bus_unit/mux28_b0_sel_is_0  (\biu/bus_unit/mux28_b0_sel_is_0_o , \biu/bus_unit/n7_neg , \biu/bus_unit/n58_neg );
  binary_mux_s1_w1 \biu/bus_unit/mux28_b1  (
    .i0(\biu/bus_unit/n59 [1]),
    .i1(\biu/bus_unit/mmu_htrans [1]),
    .sel(\biu/bus_unit/n7 ),
    .o(htrans[1]));  // ../../RTL/CPU/BIU/bus_unit.v(195)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b0  (
    .i0(\biu/write_data [0]),
    .i1(\biu/bus_unit/mmu_hwdata [0]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[0]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b1  (
    .i0(\biu/write_data [1]),
    .i1(\biu/bus_unit/mmu_hwdata [1]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[1]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b10  (
    .i0(\biu/write_data [10]),
    .i1(\biu/bus_unit/mmu_hwdata [10]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[10]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b11  (
    .i0(\biu/write_data [11]),
    .i1(\biu/bus_unit/mmu_hwdata [11]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[11]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b12  (
    .i0(\biu/write_data [12]),
    .i1(\biu/bus_unit/mmu_hwdata [12]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[12]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b13  (
    .i0(\biu/write_data [13]),
    .i1(\biu/bus_unit/mmu_hwdata [13]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[13]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b14  (
    .i0(\biu/write_data [14]),
    .i1(\biu/bus_unit/mmu_hwdata [14]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[14]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b15  (
    .i0(\biu/write_data [15]),
    .i1(\biu/bus_unit/mmu_hwdata [15]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[15]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b16  (
    .i0(\biu/write_data [16]),
    .i1(\biu/bus_unit/mmu_hwdata [16]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[16]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b17  (
    .i0(\biu/write_data [17]),
    .i1(\biu/bus_unit/mmu_hwdata [17]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[17]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b18  (
    .i0(\biu/write_data [18]),
    .i1(\biu/bus_unit/mmu_hwdata [18]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[18]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b19  (
    .i0(\biu/write_data [19]),
    .i1(\biu/bus_unit/mmu_hwdata [19]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[19]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b2  (
    .i0(\biu/write_data [2]),
    .i1(\biu/bus_unit/mmu_hwdata [2]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[2]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b20  (
    .i0(\biu/write_data [20]),
    .i1(\biu/bus_unit/mmu_hwdata [20]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[20]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b21  (
    .i0(\biu/write_data [21]),
    .i1(\biu/bus_unit/mmu_hwdata [21]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[21]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b22  (
    .i0(\biu/write_data [22]),
    .i1(\biu/bus_unit/mmu_hwdata [22]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[22]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b23  (
    .i0(\biu/write_data [23]),
    .i1(\biu/bus_unit/mmu_hwdata [23]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[23]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b24  (
    .i0(\biu/write_data [24]),
    .i1(\biu/bus_unit/mmu_hwdata [24]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[24]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b25  (
    .i0(\biu/write_data [25]),
    .i1(\biu/bus_unit/mmu_hwdata [25]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[25]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b26  (
    .i0(\biu/write_data [26]),
    .i1(\biu/bus_unit/mmu_hwdata [26]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[26]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b27  (
    .i0(\biu/write_data [27]),
    .i1(\biu/bus_unit/mmu_hwdata [27]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[27]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b28  (
    .i0(\biu/write_data [28]),
    .i1(\biu/bus_unit/mmu_hwdata [28]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[28]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b29  (
    .i0(\biu/write_data [29]),
    .i1(\biu/bus_unit/mmu_hwdata [29]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[29]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b3  (
    .i0(\biu/write_data [3]),
    .i1(\biu/bus_unit/mmu_hwdata [3]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[3]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b30  (
    .i0(\biu/write_data [30]),
    .i1(\biu/bus_unit/mmu_hwdata [30]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[30]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b31  (
    .i0(\biu/write_data [31]),
    .i1(\biu/bus_unit/mmu_hwdata [31]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[31]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b32  (
    .i0(\biu/write_data [32]),
    .i1(\biu/bus_unit/mmu_hwdata [32]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[32]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b33  (
    .i0(\biu/write_data [33]),
    .i1(\biu/bus_unit/mmu_hwdata [33]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[33]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b34  (
    .i0(\biu/write_data [34]),
    .i1(\biu/bus_unit/mmu_hwdata [34]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[34]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b35  (
    .i0(\biu/write_data [35]),
    .i1(\biu/bus_unit/mmu_hwdata [35]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[35]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b36  (
    .i0(\biu/write_data [36]),
    .i1(\biu/bus_unit/mmu_hwdata [36]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[36]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b37  (
    .i0(\biu/write_data [37]),
    .i1(\biu/bus_unit/mmu_hwdata [37]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[37]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b38  (
    .i0(\biu/write_data [38]),
    .i1(\biu/bus_unit/mmu_hwdata [38]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[38]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b39  (
    .i0(\biu/write_data [39]),
    .i1(\biu/bus_unit/mmu_hwdata [39]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[39]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b4  (
    .i0(\biu/write_data [4]),
    .i1(\biu/bus_unit/mmu_hwdata [4]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[4]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b40  (
    .i0(\biu/write_data [40]),
    .i1(\biu/bus_unit/mmu_hwdata [40]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[40]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b41  (
    .i0(\biu/write_data [41]),
    .i1(\biu/bus_unit/mmu_hwdata [41]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[41]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b42  (
    .i0(\biu/write_data [42]),
    .i1(\biu/bus_unit/mmu_hwdata [42]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[42]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b43  (
    .i0(\biu/write_data [43]),
    .i1(\biu/bus_unit/mmu_hwdata [43]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[43]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b44  (
    .i0(\biu/write_data [44]),
    .i1(\biu/bus_unit/mmu_hwdata [44]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[44]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b45  (
    .i0(\biu/write_data [45]),
    .i1(\biu/bus_unit/mmu_hwdata [45]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[45]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b46  (
    .i0(\biu/write_data [46]),
    .i1(\biu/bus_unit/mmu_hwdata [46]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[46]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b47  (
    .i0(\biu/write_data [47]),
    .i1(\biu/bus_unit/mmu_hwdata [47]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[47]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b48  (
    .i0(\biu/write_data [48]),
    .i1(\biu/bus_unit/mmu_hwdata [48]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[48]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b49  (
    .i0(\biu/write_data [49]),
    .i1(\biu/bus_unit/mmu_hwdata [49]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[49]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b5  (
    .i0(\biu/write_data [5]),
    .i1(\biu/bus_unit/mmu_hwdata [5]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[5]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b50  (
    .i0(\biu/write_data [50]),
    .i1(\biu/bus_unit/mmu_hwdata [50]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[50]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b51  (
    .i0(\biu/write_data [51]),
    .i1(\biu/bus_unit/mmu_hwdata [51]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[51]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b52  (
    .i0(\biu/write_data [52]),
    .i1(\biu/bus_unit/mmu_hwdata [52]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[52]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b53  (
    .i0(\biu/write_data [53]),
    .i1(\biu/bus_unit/mmu_hwdata [53]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[53]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b54  (
    .i0(\biu/write_data [54]),
    .i1(\biu/bus_unit/mmu_hwdata [54]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[54]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b55  (
    .i0(\biu/write_data [55]),
    .i1(\biu/bus_unit/mmu_hwdata [55]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[55]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b56  (
    .i0(\biu/write_data [56]),
    .i1(\biu/bus_unit/mmu_hwdata [56]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[56]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b57  (
    .i0(\biu/write_data [57]),
    .i1(\biu/bus_unit/mmu_hwdata [57]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[57]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b58  (
    .i0(\biu/write_data [58]),
    .i1(\biu/bus_unit/mmu_hwdata [58]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[58]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b59  (
    .i0(\biu/write_data [59]),
    .i1(\biu/bus_unit/mmu_hwdata [59]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[59]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b6  (
    .i0(\biu/write_data [6]),
    .i1(\biu/bus_unit/mmu_hwdata [6]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[6]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b60  (
    .i0(\biu/write_data [60]),
    .i1(\biu/bus_unit/mmu_hwdata [60]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[60]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b61  (
    .i0(\biu/write_data [61]),
    .i1(\biu/bus_unit/mmu_hwdata [61]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[61]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b62  (
    .i0(\biu/write_data [62]),
    .i1(\biu/bus_unit/mmu_hwdata [62]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[62]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b63  (
    .i0(\biu/write_data [63]),
    .i1(\biu/bus_unit/mmu_hwdata [63]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[63]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b7  (
    .i0(\biu/write_data [7]),
    .i1(\biu/bus_unit/mmu_hwdata [7]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[7]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b8  (
    .i0(\biu/write_data [8]),
    .i1(\biu/bus_unit/mmu_hwdata [8]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[8]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  binary_mux_s1_w1 \biu/bus_unit/mux29_b9  (
    .i0(\biu/write_data [9]),
    .i1(\biu/bus_unit/mmu_hwdata [9]),
    .sel(\biu/bus_unit/n7 ),
    .o(hwdata[9]));  // ../../RTL/CPU/BIU/bus_unit.v(197)
  AL_MUX \biu/bus_unit/mux2_b0  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\biu/bus_unit/mux2_b0_sel_is_0_o ),
    .o(\biu/bus_unit/n6 [0]));
  and \biu/bus_unit/mux2_b0_sel_is_0  (\biu/bus_unit/mux2_b0_sel_is_0_o , \biu/pa_cov_neg , \biu/bus_unit/n1_neg );
  AL_MUX \biu/bus_unit/mux2_b1  (
    .i0(1'b0),
    .i1(\biu/bus_unit/n3 ),
    .sel(\biu/bus_unit/mux2_b1_sel_is_2_o ),
    .o(\biu/bus_unit/n6 [1]));
  and \biu/bus_unit/mux2_b1_sel_is_2  (\biu/bus_unit/mux2_b1_sel_is_2_o , \biu/pa_cov_neg , \biu/bus_unit/mux1_b1_sel_is_0_o );
  AL_MUX \biu/bus_unit/mux2_b2  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\biu/bus_unit/mux2_b2_sel_is_2_o ),
    .o(\biu/bus_unit/n6 [2]));
  and \biu/bus_unit/mux2_b2_sel_is_2  (\biu/bus_unit/mux2_b2_sel_is_2_o , \biu/pa_cov_neg , \biu/bus_unit/mux1_b2_sel_is_2_o );
  AL_MUX \biu/bus_unit/mux2_b3  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\biu/bus_unit/mux2_b3_sel_is_2_o ),
    .o(\biu/bus_unit/n6 [3]));
  and \biu/bus_unit/mux2_b3_sel_is_2  (\biu/bus_unit/mux2_b3_sel_is_2_o , \biu/pa_cov_neg , \biu/bus_unit/n1 );
  binary_mux_s1_w1 \biu/bus_unit/mux30_b0  (
    .i0(hrdata[0]),
    .i1(\biu/bus_unit/mmu_hwdata [0]),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[0]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b1  (
    .i0(hrdata[1]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[1]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b10  (
    .i0(hrdata[10]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[10]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b11  (
    .i0(hrdata[11]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[11]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b12  (
    .i0(hrdata[12]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[12]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b13  (
    .i0(hrdata[13]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[13]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b14  (
    .i0(hrdata[14]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[14]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b15  (
    .i0(hrdata[15]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[15]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b16  (
    .i0(hrdata[16]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[16]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b17  (
    .i0(hrdata[17]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[17]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b18  (
    .i0(hrdata[18]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[18]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b19  (
    .i0(hrdata[19]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[19]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b2  (
    .i0(hrdata[2]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[2]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b20  (
    .i0(hrdata[20]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[20]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b21  (
    .i0(hrdata[21]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[21]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b22  (
    .i0(hrdata[22]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[22]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b23  (
    .i0(hrdata[23]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[23]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b24  (
    .i0(hrdata[24]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[24]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b25  (
    .i0(hrdata[25]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[25]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b26  (
    .i0(hrdata[26]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[26]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b27  (
    .i0(hrdata[27]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[27]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b28  (
    .i0(hrdata[28]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[28]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b29  (
    .i0(hrdata[29]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[29]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b3  (
    .i0(hrdata[3]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[3]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b30  (
    .i0(hrdata[30]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[30]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b31  (
    .i0(hrdata[31]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[31]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b32  (
    .i0(hrdata[32]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[32]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b33  (
    .i0(hrdata[33]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[33]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b34  (
    .i0(hrdata[34]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[34]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b35  (
    .i0(hrdata[35]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[35]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b36  (
    .i0(hrdata[36]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[36]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b37  (
    .i0(hrdata[37]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[37]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b38  (
    .i0(hrdata[38]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[38]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b39  (
    .i0(hrdata[39]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[39]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b4  (
    .i0(hrdata[4]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[4]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b40  (
    .i0(hrdata[40]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[40]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b41  (
    .i0(hrdata[41]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[41]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b42  (
    .i0(hrdata[42]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[42]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b43  (
    .i0(hrdata[43]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[43]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b44  (
    .i0(hrdata[44]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[44]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b45  (
    .i0(hrdata[45]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[45]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b46  (
    .i0(hrdata[46]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[46]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b47  (
    .i0(hrdata[47]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[47]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b48  (
    .i0(hrdata[48]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[48]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b49  (
    .i0(hrdata[49]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[49]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b5  (
    .i0(hrdata[5]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[5]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b50  (
    .i0(hrdata[50]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[50]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b51  (
    .i0(hrdata[51]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[51]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b52  (
    .i0(hrdata[52]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[52]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b53  (
    .i0(hrdata[53]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[53]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b54  (
    .i0(hrdata[54]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[54]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b55  (
    .i0(hrdata[55]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[55]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b56  (
    .i0(hrdata[56]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[56]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b57  (
    .i0(hrdata[57]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[57]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b58  (
    .i0(hrdata[58]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[58]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b59  (
    .i0(hrdata[59]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[59]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b6  (
    .i0(hrdata[6]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[6]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b60  (
    .i0(hrdata[60]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[60]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b61  (
    .i0(hrdata[61]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[61]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b62  (
    .i0(hrdata[62]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[62]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b63  (
    .i0(hrdata[63]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[63]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b7  (
    .i0(hrdata[7]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[7]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b8  (
    .i0(hrdata[8]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[8]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux30_b9  (
    .i0(hrdata[9]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n7 ),
    .o(uncache_data[9]));  // ../../RTL/CPU/BIU/bus_unit.v(201)
  binary_mux_s1_w1 \biu/bus_unit/mux31_b0  (
    .i0(\biu/bus_unit/last_addr [0]),
    .i1(\biu/bus_unit/addr_counter [0]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/cache_counter [0]));  // ../../RTL/CPU/BIU/bus_unit.v(207)
  binary_mux_s1_w1 \biu/bus_unit/mux31_b1  (
    .i0(\biu/bus_unit/last_addr [1]),
    .i1(\biu/bus_unit/addr_counter [1]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/cache_counter [1]));  // ../../RTL/CPU/BIU/bus_unit.v(207)
  binary_mux_s1_w1 \biu/bus_unit/mux31_b2  (
    .i0(\biu/bus_unit/last_addr [2]),
    .i1(\biu/bus_unit/addr_counter [2]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/cache_counter [2]));  // ../../RTL/CPU/BIU/bus_unit.v(207)
  binary_mux_s1_w1 \biu/bus_unit/mux31_b3  (
    .i0(\biu/bus_unit/last_addr [3]),
    .i1(\biu/bus_unit/addr_counter [3]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/cache_counter [3]));  // ../../RTL/CPU/BIU/bus_unit.v(207)
  binary_mux_s1_w1 \biu/bus_unit/mux31_b4  (
    .i0(\biu/bus_unit/last_addr [4]),
    .i1(\biu/bus_unit/addr_counter [4]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/cache_counter [4]));  // ../../RTL/CPU/BIU/bus_unit.v(207)
  binary_mux_s1_w1 \biu/bus_unit/mux31_b5  (
    .i0(\biu/bus_unit/last_addr [5]),
    .i1(\biu/bus_unit/addr_counter [5]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/cache_counter [5]));  // ../../RTL/CPU/BIU/bus_unit.v(207)
  binary_mux_s1_w1 \biu/bus_unit/mux31_b6  (
    .i0(\biu/bus_unit/last_addr [6]),
    .i1(\biu/bus_unit/addr_counter [6]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/cache_counter [6]));  // ../../RTL/CPU/BIU/bus_unit.v(207)
  binary_mux_s1_w1 \biu/bus_unit/mux31_b7  (
    .i0(\biu/bus_unit/last_addr [7]),
    .i1(\biu/bus_unit/addr_counter [7]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/cache_counter [7]));  // ../../RTL/CPU/BIU/bus_unit.v(207)
  binary_mux_s1_w1 \biu/bus_unit/mux31_b8  (
    .i0(\biu/bus_unit/last_addr [8]),
    .i1(\biu/bus_unit/addr_counter [8]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/cache_counter [8]));  // ../../RTL/CPU/BIU/bus_unit.v(207)
  binary_mux_s1_w1 \biu/bus_unit/mux3_b0  (
    .i0(\biu/bus_unit/n16 ),
    .i1(1'b1),
    .sel(hresp),
    .o(\biu/bus_unit/n17 [0]));  // ../../RTL/CPU/BIU/bus_unit.v(146)
  binary_mux_s1_w1 \biu/bus_unit/mux4_b0  (
    .i0(\biu/bus_unit/n23 [0]),
    .i1(1'b1),
    .sel(hresp),
    .o(\biu/bus_unit/n19 [0]));  // ../../RTL/CPU/BIU/bus_unit.v(149)
  binary_mux_s1_w1 \biu/bus_unit/mux7_b0  (
    .i0(\biu/bus_unit/statu [0]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n25 ),
    .o(\biu/bus_unit/n26 [0]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux7_b1  (
    .i0(\biu/bus_unit/statu [1]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n25 ),
    .o(\biu/bus_unit/n26 [1]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux7_b2  (
    .i0(\biu/bus_unit/statu [2]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n25 ),
    .o(\biu/bus_unit/n26 [2]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux7_b3  (
    .i0(\biu/bus_unit/statu [3]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n25 ),
    .o(\biu/bus_unit/n26 [3]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux7_b4  (
    .i0(\biu/bus_unit/statu [4]),
    .i1(1'b0),
    .sel(\biu/bus_unit/n25 ),
    .o(\biu/bus_unit/n26 [4]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux8_b1  (
    .i0(\biu/bus_unit/n26 [1]),
    .i1(\biu/bus_unit/n19 [0]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/bus_unit/n27 [1]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux8_b2  (
    .i0(\biu/bus_unit/n26 [2]),
    .i1(\biu/bus_unit/mmu/n36 [3]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/bus_unit/n27 [2]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux8_b3  (
    .i0(\biu/bus_unit/n26 [3]),
    .i1(\biu/bus_unit/n19 [0]),
    .sel(\biu/bus_unit/n22 ),
    .o(\biu/bus_unit/n27 [3]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  and \biu/bus_unit/mux9_b0_sel_is_0  (\biu/bus_unit/mux9_b0_sel_is_0_o , \biu/bus_unit/n20_neg , \biu/bus_unit/n22_neg );
  binary_mux_s1_w1 \biu/bus_unit/mux9_b1  (
    .i0(\biu/bus_unit/n27 [1]),
    .i1(\biu/bus_unit/mmu/n36 [3]),
    .sel(\biu/bus_unit/n20 ),
    .o(\biu/bus_unit/n28 [1]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  binary_mux_s1_w1 \biu/bus_unit/mux9_b2  (
    .i0(\biu/bus_unit/n27 [2]),
    .i1(\biu/bus_unit/n19 [0]),
    .sel(\biu/bus_unit/n20 ),
    .o(\biu/bus_unit/n28 [2]));  // ../../RTL/CPU/BIU/bus_unit.v(162)
  not \biu/bus_unit/n0_inv  (\biu/bus_unit/n0_neg , \biu/bus_unit/n0 );
  not \biu/bus_unit/n11_inv  (\biu/bus_unit/n11_neg , \biu/bus_unit/n11 );
  not \biu/bus_unit/n12_inv  (\biu/bus_unit/n12_neg , \biu/bus_unit/n12 );
  not \biu/bus_unit/n13_inv  (\biu/bus_unit/n13_neg , \biu/bus_unit/n13 );
  not \biu/bus_unit/n14_inv  (\biu/bus_unit/n14_neg , \biu/bus_unit/n14 );
  not \biu/bus_unit/n18_inv  (\biu/bus_unit/n18_neg , \biu/bus_unit/n18 );
  not \biu/bus_unit/n1_inv  (\biu/bus_unit/n1_neg , \biu/bus_unit/n1 );
  not \biu/bus_unit/n20_inv  (\biu/bus_unit/n20_neg , \biu/bus_unit/n20 );
  not \biu/bus_unit/n22_inv  (\biu/bus_unit/n22_neg , \biu/bus_unit/n22 );
  not \biu/bus_unit/n2_inv  (\biu/bus_unit/n2_neg , \biu/bus_unit/n2 );
  not \biu/bus_unit/n50_inv  (\biu/bus_unit/n50_neg , \biu/bus_unit/n50 );
  not \biu/bus_unit/n51_inv  (\biu/bus_unit/n51_neg , \biu/bus_unit/n51 );
  not \biu/bus_unit/n56_inv  (\biu/bus_unit/n56_neg , \biu/bus_unit/n56 );
  not \biu/bus_unit/n58_inv  (\biu/bus_unit/n58_neg , \biu/bus_unit/n58 );
  not \biu/bus_unit/n7_inv  (\biu/bus_unit/n7_neg , \biu/bus_unit/n7 );
  reg_sr_ss_w1 \biu/bus_unit/reg0_b0  (
    .clk(clk),
    .d(\biu/bus_unit/n39 [0]),
    .en(\biu/bus_unit/mux19_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/n37 ),
    .set(\biu/bus_unit/n15 ),
    .q(\biu/bus_unit/addr_counter [0]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_ss_w1 \biu/bus_unit/reg0_b1  (
    .clk(clk),
    .d(\biu/bus_unit/n39 [1]),
    .en(\biu/bus_unit/mux19_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/n37 ),
    .set(\biu/bus_unit/n15 ),
    .q(\biu/bus_unit/addr_counter [1]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_ss_w1 \biu/bus_unit/reg0_b2  (
    .clk(clk),
    .d(\biu/bus_unit/n39 [2]),
    .en(\biu/bus_unit/mux19_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/n37 ),
    .set(\biu/bus_unit/n15 ),
    .q(\biu/bus_unit/addr_counter [2]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_ss_w1 \biu/bus_unit/reg0_b3  (
    .clk(clk),
    .d(\biu/bus_unit/n39 [3]),
    .en(\biu/bus_unit/mux19_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/n37 ),
    .set(\biu/bus_unit/n15 ),
    .q(\biu/bus_unit/addr_counter [3]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_ss_w1 \biu/bus_unit/reg0_b4  (
    .clk(clk),
    .d(\biu/bus_unit/n39 [4]),
    .en(\biu/bus_unit/mux19_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/n37 ),
    .set(\biu/bus_unit/n15 ),
    .q(\biu/bus_unit/addr_counter [4]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_ss_w1 \biu/bus_unit/reg0_b5  (
    .clk(clk),
    .d(\biu/bus_unit/n39 [5]),
    .en(\biu/bus_unit/mux19_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/n37 ),
    .set(\biu/bus_unit/n15 ),
    .q(\biu/bus_unit/addr_counter [5]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_ss_w1 \biu/bus_unit/reg0_b6  (
    .clk(clk),
    .d(\biu/bus_unit/n39 [6]),
    .en(\biu/bus_unit/mux19_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/n37 ),
    .set(\biu/bus_unit/n15 ),
    .q(\biu/bus_unit/addr_counter [6]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_ss_w1 \biu/bus_unit/reg0_b7  (
    .clk(clk),
    .d(\biu/bus_unit/n39 [7]),
    .en(\biu/bus_unit/mux19_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/n37 ),
    .set(\biu/bus_unit/n15 ),
    .q(\biu/bus_unit/addr_counter [7]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_ss_w1 \biu/bus_unit/reg0_b8  (
    .clk(clk),
    .d(\biu/bus_unit/n39 [8]),
    .en(\biu/bus_unit/mux19_b0_sel_is_3_o ),
    .reset(\biu/bus_unit/n37 ),
    .set(\biu/bus_unit/n15 ),
    .q(\biu/bus_unit/addr_counter [8]));  // ../../RTL/CPU/BIU/bus_unit.v(177)
  reg_sr_as_w1 \biu/bus_unit/reg1_b0  (
    .clk(clk),
    .d(\biu/bus_unit/n35 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/statu [0]));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  reg_sr_as_w1 \biu/bus_unit/reg1_b1  (
    .clk(clk),
    .d(\biu/bus_unit/n35 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/statu [1]));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  reg_sr_as_w1 \biu/bus_unit/reg1_b2  (
    .clk(clk),
    .d(\biu/bus_unit/n35 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/statu [2]));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  reg_sr_as_w1 \biu/bus_unit/reg1_b3  (
    .clk(clk),
    .d(\biu/bus_unit/n35 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/bus_unit/statu [3]));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  reg_sr_as_w1 \biu/bus_unit/reg1_b4  (
    .clk(clk),
    .d(\biu/bus_unit/n30 [4]),
    .en(1'b1),
    .reset(~\biu/bus_unit/mux17_b4_sel_is_2_o ),
    .set(1'b0),
    .q(\biu/bus_unit/statu [4]));  // ../../RTL/CPU/BIU/bus_unit.v(163)
  add_pu9_mu9_o9 \biu/bus_unit/sub0  (
    .i0(\biu/bus_unit/addr_counter ),
    .i1(9'b000000001),
    .o(\biu/bus_unit/last_addr ));  // ../../RTL/CPU/BIU/bus_unit.v(203)
  or \biu/bus_unit/u10  (\biu/bus_unit/n37 , rst, \biu/bus_unit/n0 );  // ../../RTL/CPU/BIU/bus_unit.v(167)
  or \biu/bus_unit/u11  (\biu/bus_unit/n38 , \biu/bus_unit/n11 , \biu/bus_unit/n14 );  // ../../RTL/CPU/BIU/bus_unit.v(174)
  or \biu/bus_unit/u12  (\biu/bus_unit/n44 , \biu/bus_unit/n20 , \biu/bus_unit/n18 );  // ../../RTL/CPU/BIU/bus_unit.v(181)
  or \biu/bus_unit/u13  (\biu/bus_unit/n46 , \biu/bus_unit/n44 , \biu/bus_unit/n45 );  // ../../RTL/CPU/BIU/bus_unit.v(181)
  or \biu/bus_unit/u14  (\biu/bus_unit/n47 , \biu/bus_unit/n46 , \biu/bus_unit/n22 );  // ../../RTL/CPU/BIU/bus_unit.v(181)
  AL_MUX \biu/bus_unit/u15  (
    .i0(1'b0),
    .i1(hready),
    .sel(\biu/bus_unit/n47 ),
    .o(\biu/bus_unit/n48 ));  // ../../RTL/CPU/BIU/bus_unit.v(181)
  AL_MUX \biu/bus_unit/u16  (
    .i0(\biu/bus_unit/n48 ),
    .i1(\biu/bus_unit/mmu_trans_rdy ),
    .sel(\biu/bus_unit/n7 ),
    .o(\biu/trans_rdy ));  // ../../RTL/CPU/BIU/bus_unit.v(181)
  AL_MUX \biu/bus_unit/u17  (
    .i0(\biu/bus_unit/n25 ),
    .i1(\biu/bus_unit/mmu_acc_fault ),
    .sel(\biu/bus_unit/n7 ),
    .o(\biu/bus_error ));  // ../../RTL/CPU/BIU/bus_unit.v(184)
  AL_MUX \biu/bus_unit/u18  (
    .i0(1'b0),
    .i1(\biu/bus_unit/mmu_page_fault ),
    .sel(\biu/bus_unit/n7 ),
    .o(\biu/page_fault ));  // ../../RTL/CPU/BIU/bus_unit.v(185)
  AL_MUX \biu/bus_unit/u19  (
    .i0(\biu/bus_unit/n12 ),
    .i1(\biu/bus_unit/mmu_hwrite ),
    .sel(\biu/bus_unit/n7 ),
    .o(hwrite));  // ../../RTL/CPU/BIU/bus_unit.v(190)
  not \biu/bus_unit/u2  (\biu/bus_unit/n23 [0], hready);  // ../../RTL/CPU/BIU/bus_unit.v(157)
  and \biu/bus_unit/u20  (\biu/bus_unit/n50 , \biu/bus_unit/n12 , ex_size[0]);  // ../../RTL/CPU/BIU/bus_unit.v(191)
  and \biu/bus_unit/u21  (\biu/bus_unit/n51 , \biu/bus_unit/n12 , ex_size[1]);  // ../../RTL/CPU/BIU/bus_unit.v(191)
  and \biu/bus_unit/u22  (\biu/bus_unit/n52 , \biu/bus_unit/n12 , ex_size[2]);  // ../../RTL/CPU/BIU/bus_unit.v(191)
  not \biu/bus_unit/u23  (\biu/bus_unit/n53 , \biu/bus_unit/n52 );  // ../../RTL/CPU/BIU/bus_unit.v(191)
  or \biu/bus_unit/u24  (\biu/bus_unit/n56 , \biu/bus_unit/n12 , \biu/bus_unit/n13 );  // ../../RTL/CPU/BIU/bus_unit.v(193)
  or \biu/bus_unit/u26  (\biu/bus_unit/n58 , \biu/bus_unit/n56 , \biu/bus_unit/n11 );  // ../../RTL/CPU/BIU/bus_unit.v(195)
  and \biu/bus_unit/u3  (\biu/bus_unit/n1 , \biu/rd , \biu/cache_addr_sel );  // ../../RTL/CPU/BIU/bus_unit.v(127)
  or \biu/bus_unit/u32  (\biu/bus_unit/n60 , \biu/bus_unit/n14 , \biu/bus_unit/n22 );  // ../../RTL/CPU/BIU/bus_unit.v(209)
  AL_MUX \biu/bus_unit/u33  (
    .i0(1'b0),
    .i1(hready),
    .sel(\biu/bus_unit/n60 ),
    .o(\biu/cache_write ));  // ../../RTL/CPU/BIU/bus_unit.v(209)
  and \biu/bus_unit/u4  (\biu/bus_unit/n2 , \biu/rd , \biu/paddr );  // ../../RTL/CPU/BIU/bus_unit.v(127)
  or \biu/bus_unit/u5  (\biu/bus_unit/n3 , \biu/wr , \biu/new_pte_update );  // ../../RTL/CPU/BIU/bus_unit.v(127)
  or \biu/bus_unit/u6  (\biu/bus_unit/n8 , \biu/bus_unit/mmu_acc_fault , \biu/bus_unit/mmu_page_fault );  // ../../RTL/CPU/BIU/bus_unit.v(131)
  or \biu/bus_unit/u7  (\biu/bus_unit/n9 , \biu/bus_unit/n8 , \biu/bus_unit/mmu_trans_rdy );  // ../../RTL/CPU/BIU/bus_unit.v(131)
  not \biu/bus_unit/u8  (\biu/bus_unit/n10 , \biu/bus_unit/n9 );  // ../../RTL/CPU/BIU/bus_unit.v(131)
  and \biu/bus_unit/u9  (\biu/bus_unit/n16 , \biu/bus_unit/n15 , hready);  // ../../RTL/CPU/BIU/bus_unit.v(146)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d00  (
    .addra(\biu/l1d_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [7:0]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n1 ),
    .web(1'b0),
    .doa(\biu/l1d_out [7:0]));  // ../../RTL/CPU/BIU/cache.v(41)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d10  (
    .addra(\biu/l1d_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [15:8]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n3 ),
    .web(1'b0),
    .doa(\biu/l1d_out [15:8]));  // ../../RTL/CPU/BIU/cache.v(43)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d20  (
    .addra(\biu/l1d_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [23:16]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n5 ),
    .web(1'b0),
    .doa(\biu/l1d_out [23:16]));  // ../../RTL/CPU/BIU/cache.v(45)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d30  (
    .addra(\biu/l1d_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [31:24]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n7 ),
    .web(1'b0),
    .doa(\biu/l1d_out [31:24]));  // ../../RTL/CPU/BIU/cache.v(47)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d40  (
    .addra(\biu/l1d_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [39:32]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n9 ),
    .web(1'b0),
    .doa(\biu/l1d_out [39:32]));  // ../../RTL/CPU/BIU/cache.v(49)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d50  (
    .addra(\biu/l1d_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [47:40]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n11 ),
    .web(1'b0),
    .doa(\biu/l1d_out [47:40]));  // ../../RTL/CPU/BIU/cache.v(51)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d60  (
    .addra(\biu/l1d_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [55:48]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n13 ),
    .web(1'b0),
    .doa(\biu/l1d_out [55:48]));  // ../../RTL/CPU/BIU/cache.v(53)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1d70  (
    .addra(\biu/l1d_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [63:56]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n15 ),
    .web(1'b0),
    .doa(\biu/l1d_out [63:56]));  // ../../RTL/CPU/BIU/cache.v(55)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i00  (
    .addra(\biu/l1i_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [7:0]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n17 ),
    .web(1'b0),
    .doa(ins_read[7:0]));  // ../../RTL/CPU/BIU/cache.v(24)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i10  (
    .addra(\biu/l1i_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [15:8]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n19 ),
    .web(1'b0),
    .doa(ins_read[15:8]));  // ../../RTL/CPU/BIU/cache.v(26)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i20  (
    .addra(\biu/l1i_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [23:16]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n21 ),
    .web(1'b0),
    .doa(ins_read[23:16]));  // ../../RTL/CPU/BIU/cache.v(28)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i30  (
    .addra(\biu/l1i_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [31:24]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n23 ),
    .web(1'b0),
    .doa(ins_read[31:24]));  // ../../RTL/CPU/BIU/cache.v(30)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i40  (
    .addra(\biu/l1i_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [39:32]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n25 ),
    .web(1'b0),
    .doa(ins_read[39:32]));  // ../../RTL/CPU/BIU/cache.v(32)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i50  (
    .addra(\biu/l1i_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [47:40]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n27 ),
    .web(1'b0),
    .doa(ins_read[47:40]));  // ../../RTL/CPU/BIU/cache.v(34)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i60  (
    .addra(\biu/l1i_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [55:48]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n29 ),
    .web(1'b0),
    .doa(ins_read[55:48]));  // ../../RTL/CPU/BIU/cache.v(36)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(9),
    .ADDR_WIDTH_B(9),
    .BYTE_A(1),
    .BYTE_B(1),
    .BYTE_ENABLE(0),
    .DATA_DEPTH_A(512),
    .DATA_DEPTH_B(512),
    .DATA_WIDTH_A(8),
    .DATA_WIDTH_B(8),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K"),
    .MODE("SP"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"),
    .WRITEMODE_A("READBEFOREWRITE"),
    .WRITEMODE_B("NORMAL"))
    \biu/cache/ram_l1i70  (
    .addra(\biu/l1i_addr ),
    .addrb(9'b000000000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(clk),
    .clkb(1'b0),
    .dia(\biu/l1i_in [63:56]),
    .dib(8'b00000000),
    .ocea(1'b1),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(\biu/cache/n31 ),
    .web(1'b0),
    .doa(ins_read[63:56]));  // ../../RTL/CPU/BIU/cache.v(38)
  and \biu/cache/u10  (\biu/cache/n13 , \biu/l1d_write , \biu/l1d_bsel [6]);  // ../../RTL/CPU/BIU/cache.v(106)
  and \biu/cache/u11  (\biu/cache/n15 , \biu/l1d_write , \biu/l1d_bsel [7]);  // ../../RTL/CPU/BIU/cache.v(113)
  and \biu/cache/u12  (\biu/cache/n17 , \biu/l1i_write , \biu/l1i_bsel [0]);  // ../../RTL/CPU/BIU/cache.v(123)
  and \biu/cache/u13  (\biu/cache/n19 , \biu/l1i_write , \biu/l1i_bsel [1]);  // ../../RTL/CPU/BIU/cache.v(130)
  and \biu/cache/u14  (\biu/cache/n21 , \biu/l1i_write , \biu/l1i_bsel [2]);  // ../../RTL/CPU/BIU/cache.v(137)
  and \biu/cache/u15  (\biu/cache/n23 , \biu/l1i_write , \biu/l1i_bsel [3]);  // ../../RTL/CPU/BIU/cache.v(144)
  and \biu/cache/u16  (\biu/cache/n25 , \biu/l1i_write , \biu/l1i_bsel [4]);  // ../../RTL/CPU/BIU/cache.v(152)
  and \biu/cache/u17  (\biu/cache/n27 , \biu/l1i_write , \biu/l1i_bsel [5]);  // ../../RTL/CPU/BIU/cache.v(159)
  and \biu/cache/u18  (\biu/cache/n29 , \biu/l1i_write , \biu/l1i_bsel [6]);  // ../../RTL/CPU/BIU/cache.v(166)
  and \biu/cache/u19  (\biu/cache/n31 , \biu/l1i_write , \biu/l1i_bsel [7]);  // ../../RTL/CPU/BIU/cache.v(173)
  and \biu/cache/u4  (\biu/cache/n1 , \biu/l1d_write , \biu/l1d_bsel [0]);  // ../../RTL/CPU/BIU/cache.v(62)
  and \biu/cache/u5  (\biu/cache/n3 , \biu/l1d_write , \biu/l1d_bsel [1]);  // ../../RTL/CPU/BIU/cache.v(70)
  and \biu/cache/u6  (\biu/cache/n5 , \biu/l1d_write , \biu/l1d_bsel [2]);  // ../../RTL/CPU/BIU/cache.v(77)
  and \biu/cache/u7  (\biu/cache/n7 , \biu/l1d_write , \biu/l1d_bsel [3]);  // ../../RTL/CPU/BIU/cache.v(84)
  and \biu/cache/u8  (\biu/cache/n9 , \biu/l1d_write , \biu/l1d_bsel [4]);  // ../../RTL/CPU/BIU/cache.v(92)
  and \biu/cache/u9  (\biu/cache/n11 , \biu/l1d_write , \biu/l1d_bsel [5]);  // ../../RTL/CPU/BIU/cache.v(99)
  add_pu64_pu64_o64 \biu/cache_ctrl_logic/add0  (
    .i0(\biu/cache_ctrl_logic/pa_temp [63:0]),
    .i1({52'b0000000000000000000000000000000000000000000000000000,\biu/cache_ctrl_logic/off }),
    .o(\biu/cache_ctrl_logic/n207 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  add_pu64_pu64_o64 \biu/cache_ctrl_logic/add1  (
    .i0(\biu/cache_ctrl_logic/l1i_pa [63:0]),
    .i1({52'b0000000000000000000000000000000000000000000000000000,\biu/cache_ctrl_logic/off }),
    .o(\biu/cache_ctrl_logic/n209 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  add_pu64_pu64_o64 \biu/cache_ctrl_logic/add2  (
    .i0(\biu/cache_ctrl_logic/l1d_pa [63:0]),
    .i1({52'b0000000000000000000000000000000000000000000000000000,\biu/cache_ctrl_logic/off }),
    .o(\biu/cache_ctrl_logic/n212 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  eq_w52 \biu/cache_ctrl_logic/eq0  (
    .i0(\biu/cache_ctrl_logic/l1i_va [63:12]),
    .i1(addr_ex[63:12]),
    .o(\biu/cache_ctrl_logic/n3 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(187)
  eq_w52 \biu/cache_ctrl_logic/eq1  (
    .i0(\biu/cache_ctrl_logic/l1d_va [63:12]),
    .i1(addr_ex[63:12]),
    .o(\biu/cache_ctrl_logic/n5 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(188)
  eq_w5 \biu/cache_ctrl_logic/eq10  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b00000),
    .o(\biu/cache_ctrl_logic/n55 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(218)
  eq_w5 \biu/cache_ctrl_logic/eq11  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b00011),
    .o(\biu/cache_ctrl_logic/n67 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(243)
  eq_w5 \biu/cache_ctrl_logic/eq12  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b00100),
    .o(\biu/opc [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(249)
  eq_w5 \biu/cache_ctrl_logic/eq13  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b00110),
    .o(\biu/cache_ctrl_logic/l1i_wr_sel ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(253)
  eq_w5 \biu/cache_ctrl_logic/eq14  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b00111),
    .o(\biu/cache_ctrl_logic/n75 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(258)
  eq_w5 \biu/cache_ctrl_logic/eq15  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b01001),
    .o(\biu/cache_ctrl_logic/l1d_wr_sel ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(263)
  eq_w5 \biu/cache_ctrl_logic/eq16  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b01011),
    .o(\biu/wr ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(268)
  eq_w5 \biu/cache_ctrl_logic/eq17  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b01010),
    .o(\biu/ex_data_sel [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(272)
  eq_w5 \biu/cache_ctrl_logic/eq18  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b01111),
    .o(\biu/cache_ctrl_logic/n93 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(276)
  eq_w5 \biu/cache_ctrl_logic/eq19  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b10000),
    .o(\biu/cache_ctrl_logic/n97 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(279)
  eq_w52 \biu/cache_ctrl_logic/eq2  (
    .i0(\biu/cache_ctrl_logic/l1i_va [63:12]),
    .i1(addr_if[63:12]),
    .o(\biu/cache_ctrl_logic/n7 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(189)
  eq_w5 \biu/cache_ctrl_logic/eq20  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b01100),
    .o(\biu/cache_ctrl_logic/n101 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(282)
  eq_w5 \biu/cache_ctrl_logic/eq21  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b01110),
    .o(\biu/cache_ctrl_logic/n102 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(285)
  eq_w5 \biu/cache_ctrl_logic/eq22  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b01101),
    .o(\biu/cache_ctrl_logic/n104 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(288)
  eq_w5 \biu/cache_ctrl_logic/eq23  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b10010),
    .o(\biu/cache_ctrl_logic/n106 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(291)
  eq_w5 \biu/cache_ctrl_logic/eq24  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b10001),
    .o(ins_acc_fault));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(294)
  eq_w5 \biu/cache_ctrl_logic/eq25  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b10100),
    .o(\biu/cache_ctrl_logic/n107 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(297)
  eq_w5 \biu/cache_ctrl_logic/eq26  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b10011),
    .o(store_acc_fault));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(300)
  eq_w5 \biu/cache_ctrl_logic/eq27  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b10101),
    .o(\biu/cache_ctrl_logic/n108 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(303)
  eq_w5 \biu/cache_ctrl_logic/eq28  (
    .i0(\biu/cache_ctrl_logic/statu ),
    .i1(5'b10110),
    .o(load_acc_fault));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(306)
  eq_w9 \biu/cache_ctrl_logic/eq29  (
    .i0(\biu/cache_counter ),
    .i1(9'b111111111),
    .o(\biu/cache_ctrl_logic/n138 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(330)
  eq_w3 \biu/cache_ctrl_logic/eq30  (
    .i0(addr_ex[2:0]),
    .i1(3'b000),
    .o(\biu/cache_ctrl_logic/n172 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(445)
  eq_w4 \biu/cache_ctrl_logic/eq31  (
    .i0(ex_size),
    .i1(4'b0001),
    .o(\biu/cache_ctrl_logic/n173 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(445)
  eq_w4 \biu/cache_ctrl_logic/eq32  (
    .i0(ex_size),
    .i1(4'b0010),
    .o(\biu/cache_ctrl_logic/n174 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(445)
  eq_w4 \biu/cache_ctrl_logic/eq33  (
    .i0(ex_size),
    .i1(4'b0100),
    .o(\biu/cache_ctrl_logic/n176 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(445)
  eq_w4 \biu/cache_ctrl_logic/eq34  (
    .i0(ex_size),
    .i1(4'b1000),
    .o(\biu/cache_ctrl_logic/n178 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(445)
  eq_w3 \biu/cache_ctrl_logic/eq35  (
    .i0(addr_ex[2:0]),
    .i1(3'b001),
    .o(\biu/cache_ctrl_logic/n183 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(447)
  eq_w3 \biu/cache_ctrl_logic/eq36  (
    .i0(addr_ex[2:0]),
    .i1(3'b010),
    .o(\biu/cache_ctrl_logic/n187 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(450)
  eq_w3 \biu/cache_ctrl_logic/eq37  (
    .i0(addr_ex[2:0]),
    .i1(3'b011),
    .o(\biu/cache_ctrl_logic/n191 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(454)
  eq_w3 \biu/cache_ctrl_logic/eq38  (
    .i0(addr_ex[2:0]),
    .i1(3'b100),
    .o(\biu/cache_ctrl_logic/n194 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(459)
  eq_w3 \biu/cache_ctrl_logic/eq39  (
    .i0(addr_ex[2:0]),
    .i1(3'b101),
    .o(\biu/cache_ctrl_logic/n195 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(464)
  eq_w3 \biu/cache_ctrl_logic/eq4  (
    .i0({ex_priv[3],ex_priv[1:0]}),
    .i1(3'b001),
    .o(\biu/cache_ctrl_logic/n12 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(201)
  eq_w3 \biu/cache_ctrl_logic/eq40  (
    .i0(addr_ex[2:0]),
    .i1(3'b110),
    .o(\biu/cache_ctrl_logic/n196 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(469)
  eq_w3 \biu/cache_ctrl_logic/eq41  (
    .i0(addr_ex[2:0]),
    .i1(3'b111),
    .o(\biu/cache_ctrl_logic/n197 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(473)
  eq_w3 \biu/cache_ctrl_logic/eq5  (
    .i0({ex_priv[3],ex_priv[1:0]}),
    .i1(3'b010),
    .o(\biu/cache_ctrl_logic/n20 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(202)
  eq_w3 \biu/cache_ctrl_logic/eq6  (
    .i0({ex_priv[3],ex_priv[1:0]}),
    .i1(3'b100),
    .o(\biu/cache_ctrl_logic/n27 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(203)
  eq_w3 \biu/cache_ctrl_logic/eq7  (
    .i0({priv[3],priv[1:0]}),
    .i1(3'b001),
    .o(\biu/cache_ctrl_logic/n48 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(207)
  eq_w3 \biu/cache_ctrl_logic/eq8  (
    .i0({priv[3],priv[1:0]}),
    .i1(3'b010),
    .o(\biu/cache_ctrl_logic/n50 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(208)
  eq_w3 \biu/cache_ctrl_logic/eq9  (
    .i0({priv[3],priv[1:0]}),
    .i1(3'b100),
    .o(\biu/cache_ctrl_logic/n52 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(209)
  reg_sr_ss_w1 \biu/cache_ctrl_logic/l1d_value_reg  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/l1d_value ),
    .en(1'b1),
    .reset(~\biu/cache_ctrl_logic/u128_sel_is_0_o ),
    .set(\biu/cache_ctrl_logic/n149 ),
    .q(\biu/cache_ctrl_logic/l1d_value ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(394)
  reg_sr_ss_w1 \biu/cache_ctrl_logic/l1i_value_reg  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/l1i_value ),
    .en(1'b1),
    .reset(~\biu/cache_ctrl_logic/u128_sel_is_0_o ),
    .set(\biu/cache_ctrl_logic/n135 ),
    .q(\biu/cache_ctrl_logic/l1i_value ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(347)
  not \biu/cache_ctrl_logic/l1i_wr_sel_inv  (\biu/cache_ctrl_logic/l1i_wr_sel_neg , \biu/cache_ctrl_logic/l1i_wr_sel );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux0_b0  (
    .i0(\biu/cache_ctrl_logic/n60 [0]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n58 ),
    .o(\biu/cache_ctrl_logic/n61 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(223)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux0_b2  (
    .i0(\biu/cache_ctrl_logic/n60 [0]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n58 ),
    .o(\biu/cache_ctrl_logic/n61 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(223)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux0_b3  (
    .i0(\biu/cache_ctrl_logic/n59 ),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n58 ),
    .o(\biu/cache_ctrl_logic/n61 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(223)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux10_b0  (
    .i0(\biu/cache_ctrl_logic/n73 [2]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n89 ),
    .o(\biu/cache_ctrl_logic/n90 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(269)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux11_b0  (
    .i0(\biu/cache_ctrl_logic/n90 [0]),
    .i1(1'b1),
    .sel(\biu/bus_error ),
    .o(\biu/cache_ctrl_logic/n91 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(269)
  AL_MUX \biu/cache_ctrl_logic/mux11_b2  (
    .i0(1'b0),
    .i1(\biu/trans_rdy ),
    .sel(\biu/cache_ctrl_logic/mux11_b2_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n91 [2]));
  and \biu/cache_ctrl_logic/mux11_b2_sel_is_0  (\biu/cache_ctrl_logic/mux11_b2_sel_is_0_o , \biu/bus_error_neg , \biu/cache_ctrl_logic/n89_neg );
  AL_MUX \biu/cache_ctrl_logic/mux11_b3  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/mux11_b2_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n91 [3]));
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux11_b4  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\biu/bus_error ),
    .o(\biu/cache_ctrl_logic/n91 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(269)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux12_b1  (
    .i0(\biu/cache_ctrl_logic/n73 [2]),
    .i1(1'b1),
    .sel(\biu/bus_error ),
    .o(\biu/cache_ctrl_logic/n92 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(273)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux12_b3  (
    .i0(\biu/cache_ctrl_logic/n73 [2]),
    .i1(1'b0),
    .sel(\biu/bus_error ),
    .o(\biu/cache_ctrl_logic/n92 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(273)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux13_b0  (
    .i0(\biu/cache_ctrl_logic/n73 [2]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n94 ),
    .o(\biu/cache_ctrl_logic/n95 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(277)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux13_b1  (
    .i0(\biu/cache_ctrl_logic/n73 [2]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n94 ),
    .o(\biu/cache_ctrl_logic/n95 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(277)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux14_b0  (
    .i0(\biu/cache_ctrl_logic/n95 [0]),
    .i1(1'b1),
    .sel(\biu/bus_error ),
    .o(\biu/cache_ctrl_logic/n96 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(277)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux14_b1  (
    .i0(\biu/cache_ctrl_logic/n95 [1]),
    .i1(1'b1),
    .sel(\biu/bus_error ),
    .o(\biu/cache_ctrl_logic/n96 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(277)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux14_b2  (
    .i0(\biu/cache_ctrl_logic/n95 [1]),
    .i1(1'b0),
    .sel(\biu/bus_error ),
    .o(\biu/cache_ctrl_logic/n96 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(277)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux15_b0  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n98 ),
    .o(\biu/cache_ctrl_logic/n99 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(280)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux15_b4  (
    .i0(\biu/cache_ctrl_logic/n73 [2]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n98 ),
    .o(\biu/cache_ctrl_logic/n99 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(280)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux16_b0  (
    .i0(\biu/cache_ctrl_logic/n99 [0]),
    .i1(1'b1),
    .sel(\biu/bus_error ),
    .o(\biu/cache_ctrl_logic/n100 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(280)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux16_b2  (
    .i0(\biu/cache_ctrl_logic/n99 [0]),
    .i1(1'b0),
    .sel(\biu/bus_error ),
    .o(\biu/cache_ctrl_logic/n100 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(280)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux16_b4  (
    .i0(\biu/cache_ctrl_logic/n99 [4]),
    .i1(1'b1),
    .sel(\biu/bus_error ),
    .o(\biu/cache_ctrl_logic/n100 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(280)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux1_b0  (
    .i0(\biu/cache_ctrl_logic/n69 ),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n68 ),
    .o(\biu/cache_ctrl_logic/n71 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(250)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux1_b2  (
    .i0(\biu/cache_ctrl_logic/n70 [2]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n68 ),
    .o(\biu/cache_ctrl_logic/n71 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(250)
  and \biu/cache_ctrl_logic/mux20_b0_sel_is_0  (\biu/cache_ctrl_logic/mux20_b0_sel_is_0_o , \biu/cache_ctrl_logic/n108_neg , load_acc_fault_neg);
  and \biu/cache_ctrl_logic/mux21_b0_sel_is_2  (\biu/cache_ctrl_logic/mux21_b0_sel_is_2_o , store_acc_fault_neg, \biu/cache_ctrl_logic/mux20_b0_sel_is_0_o );
  and \biu/cache_ctrl_logic/mux22_b0_sel_is_2  (\biu/cache_ctrl_logic/mux22_b0_sel_is_2_o , \biu/cache_ctrl_logic/n107_neg , \biu/cache_ctrl_logic/mux21_b0_sel_is_2_o );
  and \biu/cache_ctrl_logic/mux23_b0_sel_is_2  (\biu/cache_ctrl_logic/mux23_b0_sel_is_2_o , ins_acc_fault_neg, \biu/cache_ctrl_logic/mux22_b0_sel_is_2_o );
  AL_MUX \biu/cache_ctrl_logic/mux24_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/statu [0]),
    .sel(\biu/cache_ctrl_logic/mux24_b0_sel_is_2_o ),
    .o(\biu/cache_ctrl_logic/n114 [0]));
  and \biu/cache_ctrl_logic/mux24_b0_sel_is_2  (\biu/cache_ctrl_logic/mux24_b0_sel_is_2_o , \biu/cache_ctrl_logic/n106_neg , \biu/cache_ctrl_logic/mux23_b0_sel_is_2_o );
  AL_MUX \biu/cache_ctrl_logic/mux24_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/statu [1]),
    .sel(\biu/cache_ctrl_logic/mux24_b0_sel_is_2_o ),
    .o(\biu/cache_ctrl_logic/n114 [1]));
  AL_MUX \biu/cache_ctrl_logic/mux24_b2  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/statu [2]),
    .sel(\biu/cache_ctrl_logic/mux24_b0_sel_is_2_o ),
    .o(\biu/cache_ctrl_logic/n114 [2]));
  AL_MUX \biu/cache_ctrl_logic/mux24_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/statu [3]),
    .sel(\biu/cache_ctrl_logic/mux24_b0_sel_is_2_o ),
    .o(\biu/cache_ctrl_logic/n114 [3]));
  AL_MUX \biu/cache_ctrl_logic/mux24_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/statu [4]),
    .sel(\biu/cache_ctrl_logic/mux24_b0_sel_is_2_o ),
    .o(\biu/cache_ctrl_logic/n114 [4]));
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux25_b0  (
    .i0(\biu/cache_ctrl_logic/n114 [0]),
    .i1(\biu/cache_ctrl_logic/n92 [1]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n115 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux25_b1  (
    .i0(\biu/cache_ctrl_logic/n114 [1]),
    .i1(\biu/cache_ctrl_logic/n91 [4]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n115 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux26_b0  (
    .i0(\biu/cache_ctrl_logic/n115 [0]),
    .i1(\biu/cache_ctrl_logic/n91 [4]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n116 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux26_b1  (
    .i0(\biu/cache_ctrl_logic/n115 [1]),
    .i1(\biu/cache_ctrl_logic/n92 [1]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n116 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  AL_MUX \biu/cache_ctrl_logic/mux26_b2  (
    .i0(\biu/cache_ctrl_logic/n92 [3]),
    .i1(\biu/cache_ctrl_logic/n114 [2]),
    .sel(\biu/cache_ctrl_logic/mux26_b2_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n116 [2]));
  and \biu/cache_ctrl_logic/mux26_b2_sel_is_0  (\biu/cache_ctrl_logic/mux26_b2_sel_is_0_o , \biu/cache_ctrl_logic/n102_neg , \biu/cache_ctrl_logic/n104_neg );
  AL_MUX \biu/cache_ctrl_logic/mux26_b3  (
    .i0(\biu/cache_ctrl_logic/n92 [3]),
    .i1(\biu/cache_ctrl_logic/n114 [3]),
    .sel(\biu/cache_ctrl_logic/mux26_b2_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n116 [3]));
  AL_MUX \biu/cache_ctrl_logic/mux26_b4  (
    .i0(\biu/cache_ctrl_logic/n91 [4]),
    .i1(\biu/cache_ctrl_logic/n114 [4]),
    .sel(\biu/cache_ctrl_logic/mux26_b2_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n116 [4]));
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux27_b0  (
    .i0(\biu/cache_ctrl_logic/n116 [0]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n117 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux27_b1  (
    .i0(\biu/cache_ctrl_logic/n116 [1]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n117 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux27_b2  (
    .i0(\biu/cache_ctrl_logic/n116 [2]),
    .i1(\biu/cache_ctrl_logic/n73 [2]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n117 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux27_b3  (
    .i0(\biu/cache_ctrl_logic/n116 [3]),
    .i1(\biu/cache_ctrl_logic/n73 [2]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n117 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux27_b4  (
    .i0(\biu/cache_ctrl_logic/n116 [4]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n117 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux28_b0  (
    .i0(\biu/cache_ctrl_logic/n117 [0]),
    .i1(\biu/cache_ctrl_logic/n100 [0]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n118 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux28_b1  (
    .i0(\biu/cache_ctrl_logic/n117 [1]),
    .i1(\biu/cache_ctrl_logic/n91 [4]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n118 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux28_b2  (
    .i0(\biu/cache_ctrl_logic/n117 [2]),
    .i1(\biu/cache_ctrl_logic/n100 [2]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n118 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux28_b3  (
    .i0(\biu/cache_ctrl_logic/n117 [3]),
    .i1(\biu/cache_ctrl_logic/n100 [2]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n118 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux28_b4  (
    .i0(\biu/cache_ctrl_logic/n117 [4]),
    .i1(\biu/cache_ctrl_logic/n100 [4]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n118 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux29_b0  (
    .i0(\biu/cache_ctrl_logic/n118 [0]),
    .i1(\biu/cache_ctrl_logic/n96 [0]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n119 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux29_b1  (
    .i0(\biu/cache_ctrl_logic/n118 [1]),
    .i1(\biu/cache_ctrl_logic/n96 [1]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n119 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux29_b2  (
    .i0(\biu/cache_ctrl_logic/n118 [2]),
    .i1(\biu/cache_ctrl_logic/n96 [2]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n119 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux29_b3  (
    .i0(\biu/cache_ctrl_logic/n118 [3]),
    .i1(\biu/cache_ctrl_logic/n96 [2]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n119 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux2_b0  (
    .i0(\biu/cache_ctrl_logic/n71 [0]),
    .i1(1'b0),
    .sel(\biu/page_fault ),
    .o(\biu/cache_ctrl_logic/n72 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(250)
  AL_MUX \biu/cache_ctrl_logic/mux2_b1  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/mux2_b1_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n72 [1]));
  and \biu/cache_ctrl_logic/mux2_b1_sel_is_0  (\biu/cache_ctrl_logic/mux2_b1_sel_is_0_o , \biu/page_fault_neg , \biu/cache_ctrl_logic/n68_neg );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux2_b2  (
    .i0(\biu/cache_ctrl_logic/n71 [2]),
    .i1(1'b0),
    .sel(\biu/page_fault ),
    .o(\biu/cache_ctrl_logic/n72 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(250)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux2_b4  (
    .i0(\biu/cache_ctrl_logic/n71 [0]),
    .i1(1'b1),
    .sel(\biu/page_fault ),
    .o(\biu/cache_ctrl_logic/n72 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(250)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux30_b0  (
    .i0(\biu/cache_ctrl_logic/n119 [0]),
    .i1(1'b0),
    .sel(\biu/ex_data_sel [1]),
    .o(\biu/cache_ctrl_logic/n120 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux30_b1  (
    .i0(\biu/cache_ctrl_logic/n119 [1]),
    .i1(\biu/cache_ctrl_logic/n92 [1]),
    .sel(\biu/ex_data_sel [1]),
    .o(\biu/cache_ctrl_logic/n120 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux30_b2  (
    .i0(\biu/cache_ctrl_logic/n119 [2]),
    .i1(\biu/cache_ctrl_logic/n91 [4]),
    .sel(\biu/ex_data_sel [1]),
    .o(\biu/cache_ctrl_logic/n120 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux30_b3  (
    .i0(\biu/cache_ctrl_logic/n119 [3]),
    .i1(\biu/cache_ctrl_logic/n92 [3]),
    .sel(\biu/ex_data_sel [1]),
    .o(\biu/cache_ctrl_logic/n120 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  and \biu/cache_ctrl_logic/mux30_b4_sel_is_0  (\biu/cache_ctrl_logic/mux30_b4_sel_is_0_o , \biu/ex_data_sel[1]_neg , \biu/cache_ctrl_logic/n93_neg );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux31_b0  (
    .i0(\biu/cache_ctrl_logic/n120 [0]),
    .i1(\biu/cache_ctrl_logic/n91 [0]),
    .sel(\biu/wr ),
    .o(\biu/cache_ctrl_logic/n121 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux31_b1  (
    .i0(\biu/cache_ctrl_logic/n120 [1]),
    .i1(\biu/cache_ctrl_logic/n91 [0]),
    .sel(\biu/wr ),
    .o(\biu/cache_ctrl_logic/n121 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux31_b2  (
    .i0(\biu/cache_ctrl_logic/n120 [2]),
    .i1(\biu/cache_ctrl_logic/n91 [2]),
    .sel(\biu/wr ),
    .o(\biu/cache_ctrl_logic/n121 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux31_b3  (
    .i0(\biu/cache_ctrl_logic/n120 [3]),
    .i1(\biu/cache_ctrl_logic/n91 [3]),
    .sel(\biu/wr ),
    .o(\biu/cache_ctrl_logic/n121 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  AL_MUX \biu/cache_ctrl_logic/mux31_b4  (
    .i0(\biu/cache_ctrl_logic/n91 [4]),
    .i1(\biu/cache_ctrl_logic/n118 [4]),
    .sel(\biu/cache_ctrl_logic/mux31_b4_sel_is_2_o ),
    .o(\biu/cache_ctrl_logic/n121 [4]));
  and \biu/cache_ctrl_logic/mux31_b4_sel_is_2  (\biu/cache_ctrl_logic/mux31_b4_sel_is_2_o , \biu/wr_neg , \biu/cache_ctrl_logic/mux30_b4_sel_is_0_o );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux32_b0  (
    .i0(\biu/cache_ctrl_logic/n121 [0]),
    .i1(\biu/cache_ctrl_logic/n88 [0]),
    .sel(\biu/cache_ctrl_logic/l1d_wr_sel ),
    .o(\biu/cache_ctrl_logic/n122 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux32_b1  (
    .i0(\biu/cache_ctrl_logic/n121 [1]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/l1d_wr_sel ),
    .o(\biu/cache_ctrl_logic/n122 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux32_b2  (
    .i0(\biu/cache_ctrl_logic/n121 [2]),
    .i1(\biu/cache_ctrl_logic/n88 [2]),
    .sel(\biu/cache_ctrl_logic/l1d_wr_sel ),
    .o(\biu/cache_ctrl_logic/n122 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux32_b3  (
    .i0(\biu/cache_ctrl_logic/n121 [3]),
    .i1(\biu/cache_ctrl_logic/n88 [3]),
    .sel(\biu/cache_ctrl_logic/l1d_wr_sel ),
    .o(\biu/cache_ctrl_logic/n122 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux32_b4  (
    .i0(\biu/cache_ctrl_logic/n121 [4]),
    .i1(\biu/cache_ctrl_logic/n88 [2]),
    .sel(\biu/cache_ctrl_logic/l1d_wr_sel ),
    .o(\biu/cache_ctrl_logic/n122 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux33_b0  (
    .i0(\biu/cache_ctrl_logic/n122 [0]),
    .i1(\biu/cache_ctrl_logic/n84 [0]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n123 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux33_b1  (
    .i0(\biu/cache_ctrl_logic/n122 [1]),
    .i1(\biu/cache_ctrl_logic/n84 [1]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n123 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux33_b2  (
    .i0(\biu/cache_ctrl_logic/n122 [2]),
    .i1(\biu/cache_ctrl_logic/n84 [2]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n123 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux33_b3  (
    .i0(\biu/cache_ctrl_logic/n122 [3]),
    .i1(\biu/cache_ctrl_logic/n84 [3]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n123 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux33_b4  (
    .i0(\biu/cache_ctrl_logic/n122 [4]),
    .i1(\biu/cache_ctrl_logic/n84 [4]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n123 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux34_b0  (
    .i0(\biu/cache_ctrl_logic/n123 [0]),
    .i1(\biu/cache_ctrl_logic/n91 [4]),
    .sel(\biu/cache_ctrl_logic/l1i_wr_sel ),
    .o(\biu/cache_ctrl_logic/n124 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux34_b1  (
    .i0(\biu/cache_ctrl_logic/n123 [1]),
    .i1(\biu/cache_ctrl_logic/n92 [3]),
    .sel(\biu/cache_ctrl_logic/l1i_wr_sel ),
    .o(\biu/cache_ctrl_logic/n124 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux34_b2  (
    .i0(\biu/cache_ctrl_logic/n123 [2]),
    .i1(\biu/cache_ctrl_logic/n92 [3]),
    .sel(\biu/cache_ctrl_logic/l1i_wr_sel ),
    .o(\biu/cache_ctrl_logic/n124 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux34_b4  (
    .i0(\biu/cache_ctrl_logic/n123 [4]),
    .i1(\biu/cache_ctrl_logic/n91 [4]),
    .sel(\biu/cache_ctrl_logic/l1i_wr_sel ),
    .o(\biu/cache_ctrl_logic/n124 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux35_b0  (
    .i0(\biu/cache_ctrl_logic/n124 [0]),
    .i1(\biu/cache_ctrl_logic/n72 [0]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n125 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux35_b1  (
    .i0(\biu/cache_ctrl_logic/n124 [1]),
    .i1(\biu/cache_ctrl_logic/n72 [1]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n125 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux35_b2  (
    .i0(\biu/cache_ctrl_logic/n124 [2]),
    .i1(\biu/cache_ctrl_logic/n72 [2]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n125 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  and \biu/cache_ctrl_logic/mux35_b3_sel_is_0  (\biu/cache_ctrl_logic/mux35_b3_sel_is_0_o , \biu/opc[1]_neg , \biu/cache_ctrl_logic/l1i_wr_sel_neg );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux35_b4  (
    .i0(\biu/cache_ctrl_logic/n124 [4]),
    .i1(\biu/cache_ctrl_logic/n72 [4]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n125 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux36_b0  (
    .i0(\biu/cache_ctrl_logic/n125 [0]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n67 ),
    .o(\biu/cache_ctrl_logic/n126 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux36_b1  (
    .i0(\biu/cache_ctrl_logic/n125 [1]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n67 ),
    .o(\biu/cache_ctrl_logic/n126 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux36_b2  (
    .i0(\biu/cache_ctrl_logic/n125 [2]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n67 ),
    .o(\biu/cache_ctrl_logic/n126 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  AL_MUX \biu/cache_ctrl_logic/mux36_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n123 [3]),
    .sel(\biu/cache_ctrl_logic/mux36_b3_sel_is_2_o ),
    .o(\biu/cache_ctrl_logic/n126 [3]));
  and \biu/cache_ctrl_logic/mux36_b3_sel_is_2  (\biu/cache_ctrl_logic/mux36_b3_sel_is_2_o , \biu/cache_ctrl_logic/n67_neg , \biu/cache_ctrl_logic/mux35_b3_sel_is_0_o );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux37_b0  (
    .i0(\biu/cache_ctrl_logic/n126 [0]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n66 ),
    .o(\biu/cache_ctrl_logic/n127 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux37_b1  (
    .i0(\biu/cache_ctrl_logic/n126 [1]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n66 ),
    .o(\biu/cache_ctrl_logic/n127 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux37_b2  (
    .i0(\biu/cache_ctrl_logic/n126 [2]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n66 ),
    .o(\biu/cache_ctrl_logic/n127 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux37_b3  (
    .i0(\biu/cache_ctrl_logic/n126 [3]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n66 ),
    .o(\biu/cache_ctrl_logic/n127 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  AL_MUX \biu/cache_ctrl_logic/mux37_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n125 [4]),
    .sel(\biu/cache_ctrl_logic/mux37_b4_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n127 [4]));
  and \biu/cache_ctrl_logic/mux37_b4_sel_is_0  (\biu/cache_ctrl_logic/mux37_b4_sel_is_0_o , \biu/cache_ctrl_logic/n66_neg , \biu/cache_ctrl_logic/n67_neg );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux38_b1  (
    .i0(\biu/cache_ctrl_logic/n127 [1]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n65 ),
    .o(\biu/cache_ctrl_logic/n128 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux38_b2  (
    .i0(\biu/cache_ctrl_logic/n127 [2]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n65 ),
    .o(\biu/cache_ctrl_logic/n128 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux38_b3  (
    .i0(\biu/cache_ctrl_logic/n127 [3]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n65 ),
    .o(\biu/cache_ctrl_logic/n128 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  AL_MUX \biu/cache_ctrl_logic/mux39_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n127 [0]),
    .sel(\biu/cache_ctrl_logic/mux39_b0_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n129 [0]));
  and \biu/cache_ctrl_logic/mux39_b0_sel_is_0  (\biu/cache_ctrl_logic/mux39_b0_sel_is_0_o , \biu/cache_ctrl_logic/n64_neg , \biu/cache_ctrl_logic/n65_neg );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux39_b1  (
    .i0(\biu/cache_ctrl_logic/n128 [1]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n64 ),
    .o(\biu/cache_ctrl_logic/n129 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux40_b0  (
    .i0(\biu/cache_ctrl_logic/n129 [0]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n63 ),
    .o(\biu/cache_ctrl_logic/n130 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  and \biu/cache_ctrl_logic/mux40_b2_sel_is_0  (\biu/cache_ctrl_logic/mux40_b2_sel_is_0_o , \biu/cache_ctrl_logic/n63_neg , \biu/cache_ctrl_logic/n64_neg );
  AL_MUX \biu/cache_ctrl_logic/mux40_b3  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/n128 [3]),
    .sel(\biu/cache_ctrl_logic/mux40_b2_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n130 [3]));
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux41_b0  (
    .i0(\biu/cache_ctrl_logic/n130 [0]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n62 ),
    .o(\biu/cache_ctrl_logic/n131 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  AL_MUX \biu/cache_ctrl_logic/mux41_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n129 [1]),
    .sel(\biu/cache_ctrl_logic/mux41_b1_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n131 [1]));
  and \biu/cache_ctrl_logic/mux41_b1_sel_is_0  (\biu/cache_ctrl_logic/mux41_b1_sel_is_0_o , \biu/cache_ctrl_logic/n62_neg , \biu/cache_ctrl_logic/n63_neg );
  AL_MUX \biu/cache_ctrl_logic/mux41_b2  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/n128 [2]),
    .sel(\biu/cache_ctrl_logic/mux41_b2_sel_is_2_o ),
    .o(\biu/cache_ctrl_logic/n131 [2]));
  and \biu/cache_ctrl_logic/mux41_b2_sel_is_2  (\biu/cache_ctrl_logic/mux41_b2_sel_is_2_o , \biu/cache_ctrl_logic/n62_neg , \biu/cache_ctrl_logic/mux40_b2_sel_is_0_o );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux41_b3  (
    .i0(\biu/cache_ctrl_logic/n130 [3]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n62 ),
    .o(\biu/cache_ctrl_logic/n131 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux42_b0  (
    .i0(\biu/cache_ctrl_logic/n131 [0]),
    .i1(\biu/cache_ctrl_logic/n61 [0]),
    .sel(\biu/cache_ctrl_logic/n57 ),
    .o(\biu/cache_ctrl_logic/n132 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux42_b2  (
    .i0(\biu/cache_ctrl_logic/n131 [2]),
    .i1(\biu/cache_ctrl_logic/n61 [2]),
    .sel(\biu/cache_ctrl_logic/n57 ),
    .o(\biu/cache_ctrl_logic/n132 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux42_b3  (
    .i0(\biu/cache_ctrl_logic/n131 [3]),
    .i1(\biu/cache_ctrl_logic/n61 [3]),
    .sel(\biu/cache_ctrl_logic/n57 ),
    .o(\biu/cache_ctrl_logic/n132 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(311)
  and \biu/cache_ctrl_logic/mux42_b4_sel_is_2  (\biu/cache_ctrl_logic/mux42_b4_sel_is_2_o , \biu/cache_ctrl_logic/n57_neg , \biu/cache_ctrl_logic/mux41_b2_sel_is_2_o );
  and \biu/cache_ctrl_logic/mux43_b1_sel_is_0  (\biu/cache_ctrl_logic/mux43_b1_sel_is_0_o , \biu/cache_ctrl_logic/n56_neg , \biu/cache_ctrl_logic/n57_neg );
  and \biu/cache_ctrl_logic/mux43_b4_sel_is_2  (\biu/cache_ctrl_logic/mux43_b4_sel_is_2_o , \biu/cache_ctrl_logic/n56_neg , \biu/cache_ctrl_logic/mux42_b4_sel_is_2_o );
  and \biu/cache_ctrl_logic/mux44_b2_sel_is_0  (\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o , rst_neg, \biu/cache_ctrl_logic/n56_neg );
  and \biu/cache_ctrl_logic/mux44_b4_sel_is_2  (\biu/cache_ctrl_logic/mux44_b4_sel_is_2_o , rst_neg, \biu/cache_ctrl_logic/mux43_b4_sel_is_2_o );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux49_b7  (
    .i0(\biu/cache_ctrl_logic/n146 ),
    .i1(\biu/cache_ctrl_logic/pte_temp [7]),
    .sel(\biu/cache_ctrl_logic/n135 ),
    .o(\biu/cache_ctrl_logic/n147 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(361)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux4_b0  (
    .i0(\biu/cache_ctrl_logic/n80 [2]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n78 ),
    .o(\biu/cache_ctrl_logic/n81 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux4_b2  (
    .i0(\biu/cache_ctrl_logic/n80 [2]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n78 ),
    .o(\biu/cache_ctrl_logic/n81 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux4_b3  (
    .i0(\biu/cache_ctrl_logic/n79 ),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n78 ),
    .o(\biu/cache_ctrl_logic/n81 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux55_b7  (
    .i0(\biu/cache_ctrl_logic/n157 ),
    .i1(\biu/cache_ctrl_logic/pte_temp [7]),
    .sel(\biu/cache_ctrl_logic/n149 ),
    .o(\biu/cache_ctrl_logic/n158 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(406)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b0  (
    .i0(\biu/cache_ctrl_logic/pa_temp [0]),
    .i1(\biu/paddress [0]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b1  (
    .i0(\biu/cache_ctrl_logic/pa_temp [1]),
    .i1(\biu/paddress [1]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b10  (
    .i0(\biu/cache_ctrl_logic/pa_temp [10]),
    .i1(\biu/paddress [10]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b11  (
    .i0(\biu/cache_ctrl_logic/pa_temp [11]),
    .i1(\biu/paddress [11]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b12  (
    .i0(\biu/cache_ctrl_logic/pa_temp [12]),
    .i1(\biu/paddress [12]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b13  (
    .i0(\biu/cache_ctrl_logic/pa_temp [13]),
    .i1(\biu/paddress [13]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b14  (
    .i0(\biu/cache_ctrl_logic/pa_temp [14]),
    .i1(\biu/paddress [14]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b15  (
    .i0(\biu/cache_ctrl_logic/pa_temp [15]),
    .i1(\biu/paddress [15]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b16  (
    .i0(\biu/cache_ctrl_logic/pa_temp [16]),
    .i1(\biu/paddress [16]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b17  (
    .i0(\biu/cache_ctrl_logic/pa_temp [17]),
    .i1(\biu/paddress [17]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b18  (
    .i0(\biu/cache_ctrl_logic/pa_temp [18]),
    .i1(\biu/paddress [18]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b19  (
    .i0(\biu/cache_ctrl_logic/pa_temp [19]),
    .i1(\biu/paddress [19]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b2  (
    .i0(\biu/cache_ctrl_logic/pa_temp [2]),
    .i1(\biu/paddress [2]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b20  (
    .i0(\biu/cache_ctrl_logic/pa_temp [20]),
    .i1(\biu/paddress [20]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b21  (
    .i0(\biu/cache_ctrl_logic/pa_temp [21]),
    .i1(\biu/paddress [21]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b22  (
    .i0(\biu/cache_ctrl_logic/pa_temp [22]),
    .i1(\biu/paddress [22]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b23  (
    .i0(\biu/cache_ctrl_logic/pa_temp [23]),
    .i1(\biu/paddress [23]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b24  (
    .i0(\biu/cache_ctrl_logic/pa_temp [24]),
    .i1(\biu/paddress [24]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b25  (
    .i0(\biu/cache_ctrl_logic/pa_temp [25]),
    .i1(\biu/paddress [25]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b26  (
    .i0(\biu/cache_ctrl_logic/pa_temp [26]),
    .i1(\biu/paddress [26]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b27  (
    .i0(\biu/cache_ctrl_logic/pa_temp [27]),
    .i1(\biu/paddress [27]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b28  (
    .i0(\biu/cache_ctrl_logic/pa_temp [28]),
    .i1(\biu/paddress [28]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b29  (
    .i0(\biu/cache_ctrl_logic/pa_temp [29]),
    .i1(\biu/paddress [29]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b3  (
    .i0(\biu/cache_ctrl_logic/pa_temp [3]),
    .i1(\biu/paddress [3]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b30  (
    .i0(\biu/cache_ctrl_logic/pa_temp [30]),
    .i1(\biu/paddress [30]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b31  (
    .i0(\biu/cache_ctrl_logic/pa_temp [31]),
    .i1(\biu/paddress [31]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b32  (
    .i0(\biu/cache_ctrl_logic/pa_temp [32]),
    .i1(\biu/paddress [32]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b33  (
    .i0(\biu/cache_ctrl_logic/pa_temp [33]),
    .i1(\biu/paddress [33]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b34  (
    .i0(\biu/cache_ctrl_logic/pa_temp [34]),
    .i1(\biu/paddress [34]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b35  (
    .i0(\biu/cache_ctrl_logic/pa_temp [35]),
    .i1(\biu/paddress [35]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b36  (
    .i0(\biu/cache_ctrl_logic/pa_temp [36]),
    .i1(\biu/paddress [36]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b37  (
    .i0(\biu/cache_ctrl_logic/pa_temp [37]),
    .i1(\biu/paddress [37]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b38  (
    .i0(\biu/cache_ctrl_logic/pa_temp [38]),
    .i1(\biu/paddress [38]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b39  (
    .i0(\biu/cache_ctrl_logic/pa_temp [39]),
    .i1(\biu/paddress [39]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b4  (
    .i0(\biu/cache_ctrl_logic/pa_temp [4]),
    .i1(\biu/paddress [4]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b40  (
    .i0(\biu/cache_ctrl_logic/pa_temp [40]),
    .i1(\biu/paddress [40]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b41  (
    .i0(\biu/cache_ctrl_logic/pa_temp [41]),
    .i1(\biu/paddress [41]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b42  (
    .i0(\biu/cache_ctrl_logic/pa_temp [42]),
    .i1(\biu/paddress [42]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b43  (
    .i0(\biu/cache_ctrl_logic/pa_temp [43]),
    .i1(\biu/paddress [43]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b44  (
    .i0(\biu/cache_ctrl_logic/pa_temp [44]),
    .i1(\biu/paddress [44]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b45  (
    .i0(\biu/cache_ctrl_logic/pa_temp [45]),
    .i1(\biu/paddress [45]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b46  (
    .i0(\biu/cache_ctrl_logic/pa_temp [46]),
    .i1(\biu/paddress [46]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b47  (
    .i0(\biu/cache_ctrl_logic/pa_temp [47]),
    .i1(\biu/paddress [47]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b48  (
    .i0(\biu/cache_ctrl_logic/pa_temp [48]),
    .i1(\biu/paddress [48]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b49  (
    .i0(\biu/cache_ctrl_logic/pa_temp [49]),
    .i1(\biu/paddress [49]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b5  (
    .i0(\biu/cache_ctrl_logic/pa_temp [5]),
    .i1(\biu/paddress [5]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b50  (
    .i0(\biu/cache_ctrl_logic/pa_temp [50]),
    .i1(\biu/paddress [50]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b51  (
    .i0(\biu/cache_ctrl_logic/pa_temp [51]),
    .i1(\biu/paddress [51]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b52  (
    .i0(\biu/cache_ctrl_logic/pa_temp [52]),
    .i1(\biu/paddress [52]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b53  (
    .i0(\biu/cache_ctrl_logic/pa_temp [53]),
    .i1(\biu/paddress [53]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b54  (
    .i0(\biu/cache_ctrl_logic/pa_temp [54]),
    .i1(\biu/paddress [54]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b55  (
    .i0(\biu/cache_ctrl_logic/pa_temp [55]),
    .i1(\biu/paddress [55]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b56  (
    .i0(\biu/cache_ctrl_logic/pa_temp [56]),
    .i1(\biu/paddress [56]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b57  (
    .i0(\biu/cache_ctrl_logic/pa_temp [57]),
    .i1(\biu/paddress [57]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b58  (
    .i0(\biu/cache_ctrl_logic/pa_temp [58]),
    .i1(\biu/paddress [58]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b59  (
    .i0(\biu/cache_ctrl_logic/pa_temp [59]),
    .i1(\biu/paddress [59]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b6  (
    .i0(\biu/cache_ctrl_logic/pa_temp [6]),
    .i1(\biu/paddress [6]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b60  (
    .i0(\biu/cache_ctrl_logic/pa_temp [60]),
    .i1(\biu/paddress [60]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b61  (
    .i0(\biu/cache_ctrl_logic/pa_temp [61]),
    .i1(\biu/paddress [61]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b62  (
    .i0(\biu/cache_ctrl_logic/pa_temp [62]),
    .i1(\biu/paddress [62]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b63  (
    .i0(\biu/cache_ctrl_logic/pa_temp [63]),
    .i1(\biu/paddress [63]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b7  (
    .i0(\biu/cache_ctrl_logic/pa_temp [7]),
    .i1(\biu/paddress [7]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b8  (
    .i0(\biu/cache_ctrl_logic/pa_temp [8]),
    .i1(\biu/paddress [8]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux57_b9  (
    .i0(\biu/cache_ctrl_logic/pa_temp [9]),
    .i1(\biu/paddress [9]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n164 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux58_b7  (
    .i0(\biu/cache_ctrl_logic/n163 ),
    .i1(uncache_data[7]),
    .sel(\biu/cache_ctrl_logic/n162 ),
    .o(\biu/cache_ctrl_logic/n165 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b0  (
    .i0(\biu/cache_ctrl_logic/n164 [0]),
    .i1(addr_ex[0]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b1  (
    .i0(\biu/cache_ctrl_logic/n164 [1]),
    .i1(addr_ex[1]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b10  (
    .i0(\biu/cache_ctrl_logic/n164 [10]),
    .i1(addr_ex[10]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  and \biu/cache_ctrl_logic/mux59_b100_sel_is_2  (\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o , \biu/cache_ctrl_logic/n161_neg , \biu/cache_ctrl_logic/n162 );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b11  (
    .i0(\biu/cache_ctrl_logic/n164 [11]),
    .i1(addr_ex[11]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b12  (
    .i0(\biu/cache_ctrl_logic/n164 [12]),
    .i1(addr_ex[12]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b13  (
    .i0(\biu/cache_ctrl_logic/n164 [13]),
    .i1(addr_ex[13]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b14  (
    .i0(\biu/cache_ctrl_logic/n164 [14]),
    .i1(addr_ex[14]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b15  (
    .i0(\biu/cache_ctrl_logic/n164 [15]),
    .i1(addr_ex[15]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b16  (
    .i0(\biu/cache_ctrl_logic/n164 [16]),
    .i1(addr_ex[16]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b17  (
    .i0(\biu/cache_ctrl_logic/n164 [17]),
    .i1(addr_ex[17]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b18  (
    .i0(\biu/cache_ctrl_logic/n164 [18]),
    .i1(addr_ex[18]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b19  (
    .i0(\biu/cache_ctrl_logic/n164 [19]),
    .i1(addr_ex[19]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b2  (
    .i0(\biu/cache_ctrl_logic/n164 [2]),
    .i1(addr_ex[2]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b20  (
    .i0(\biu/cache_ctrl_logic/n164 [20]),
    .i1(addr_ex[20]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b21  (
    .i0(\biu/cache_ctrl_logic/n164 [21]),
    .i1(addr_ex[21]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b22  (
    .i0(\biu/cache_ctrl_logic/n164 [22]),
    .i1(addr_ex[22]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b23  (
    .i0(\biu/cache_ctrl_logic/n164 [23]),
    .i1(addr_ex[23]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b24  (
    .i0(\biu/cache_ctrl_logic/n164 [24]),
    .i1(addr_ex[24]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b25  (
    .i0(\biu/cache_ctrl_logic/n164 [25]),
    .i1(addr_ex[25]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b26  (
    .i0(\biu/cache_ctrl_logic/n164 [26]),
    .i1(addr_ex[26]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b27  (
    .i0(\biu/cache_ctrl_logic/n164 [27]),
    .i1(addr_ex[27]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b28  (
    .i0(\biu/cache_ctrl_logic/n164 [28]),
    .i1(addr_ex[28]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b29  (
    .i0(\biu/cache_ctrl_logic/n164 [29]),
    .i1(addr_ex[29]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b3  (
    .i0(\biu/cache_ctrl_logic/n164 [3]),
    .i1(addr_ex[3]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b30  (
    .i0(\biu/cache_ctrl_logic/n164 [30]),
    .i1(addr_ex[30]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b31  (
    .i0(\biu/cache_ctrl_logic/n164 [31]),
    .i1(addr_ex[31]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b32  (
    .i0(\biu/cache_ctrl_logic/n164 [32]),
    .i1(addr_ex[32]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b33  (
    .i0(\biu/cache_ctrl_logic/n164 [33]),
    .i1(addr_ex[33]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b34  (
    .i0(\biu/cache_ctrl_logic/n164 [34]),
    .i1(addr_ex[34]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b35  (
    .i0(\biu/cache_ctrl_logic/n164 [35]),
    .i1(addr_ex[35]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b36  (
    .i0(\biu/cache_ctrl_logic/n164 [36]),
    .i1(addr_ex[36]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b37  (
    .i0(\biu/cache_ctrl_logic/n164 [37]),
    .i1(addr_ex[37]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b38  (
    .i0(\biu/cache_ctrl_logic/n164 [38]),
    .i1(addr_ex[38]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b39  (
    .i0(\biu/cache_ctrl_logic/n164 [39]),
    .i1(addr_ex[39]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b4  (
    .i0(\biu/cache_ctrl_logic/n164 [4]),
    .i1(addr_ex[4]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b40  (
    .i0(\biu/cache_ctrl_logic/n164 [40]),
    .i1(addr_ex[40]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b41  (
    .i0(\biu/cache_ctrl_logic/n164 [41]),
    .i1(addr_ex[41]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b42  (
    .i0(\biu/cache_ctrl_logic/n164 [42]),
    .i1(addr_ex[42]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b43  (
    .i0(\biu/cache_ctrl_logic/n164 [43]),
    .i1(addr_ex[43]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b44  (
    .i0(\biu/cache_ctrl_logic/n164 [44]),
    .i1(addr_ex[44]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b45  (
    .i0(\biu/cache_ctrl_logic/n164 [45]),
    .i1(addr_ex[45]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b46  (
    .i0(\biu/cache_ctrl_logic/n164 [46]),
    .i1(addr_ex[46]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b47  (
    .i0(\biu/cache_ctrl_logic/n164 [47]),
    .i1(addr_ex[47]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b48  (
    .i0(\biu/cache_ctrl_logic/n164 [48]),
    .i1(addr_ex[48]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b49  (
    .i0(\biu/cache_ctrl_logic/n164 [49]),
    .i1(addr_ex[49]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b5  (
    .i0(\biu/cache_ctrl_logic/n164 [5]),
    .i1(addr_ex[5]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b50  (
    .i0(\biu/cache_ctrl_logic/n164 [50]),
    .i1(addr_ex[50]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b51  (
    .i0(\biu/cache_ctrl_logic/n164 [51]),
    .i1(addr_ex[51]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b52  (
    .i0(\biu/cache_ctrl_logic/n164 [52]),
    .i1(addr_ex[52]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b53  (
    .i0(\biu/cache_ctrl_logic/n164 [53]),
    .i1(addr_ex[53]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b54  (
    .i0(\biu/cache_ctrl_logic/n164 [54]),
    .i1(addr_ex[54]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b55  (
    .i0(\biu/cache_ctrl_logic/n164 [55]),
    .i1(addr_ex[55]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b56  (
    .i0(\biu/cache_ctrl_logic/n164 [56]),
    .i1(addr_ex[56]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b57  (
    .i0(\biu/cache_ctrl_logic/n164 [57]),
    .i1(addr_ex[57]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b58  (
    .i0(\biu/cache_ctrl_logic/n164 [58]),
    .i1(addr_ex[58]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b59  (
    .i0(\biu/cache_ctrl_logic/n164 [59]),
    .i1(addr_ex[59]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b6  (
    .i0(\biu/cache_ctrl_logic/n164 [6]),
    .i1(addr_ex[6]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b60  (
    .i0(\biu/cache_ctrl_logic/n164 [60]),
    .i1(addr_ex[60]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b61  (
    .i0(\biu/cache_ctrl_logic/n164 [61]),
    .i1(addr_ex[61]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b62  (
    .i0(\biu/cache_ctrl_logic/n164 [62]),
    .i1(addr_ex[62]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b63  (
    .i0(\biu/cache_ctrl_logic/n164 [63]),
    .i1(addr_ex[63]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b7  (
    .i0(\biu/cache_ctrl_logic/n164 [7]),
    .i1(addr_ex[7]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b8  (
    .i0(\biu/cache_ctrl_logic/n164 [8]),
    .i1(addr_ex[8]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux59_b9  (
    .i0(\biu/cache_ctrl_logic/n164 [9]),
    .i1(addr_ex[9]),
    .sel(\biu/cache_ctrl_logic/n161 ),
    .o(\biu/cache_ctrl_logic/n166 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux5_b0  (
    .i0(\biu/cache_ctrl_logic/n81 [0]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n68 ),
    .o(\biu/cache_ctrl_logic/n82 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux63_b0  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [0]),
    .sel(\biu/cache_ctrl_logic/n170 ),
    .o(\biu/l1i_bsel [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(440)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux63_b1  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [1]),
    .sel(\biu/cache_ctrl_logic/n170 ),
    .o(\biu/l1i_bsel [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(440)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux63_b2  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [2]),
    .sel(\biu/cache_ctrl_logic/n170 ),
    .o(\biu/l1i_bsel [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(440)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux63_b3  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [3]),
    .sel(\biu/cache_ctrl_logic/n170 ),
    .o(\biu/l1i_bsel [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(440)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux63_b4  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [4]),
    .sel(\biu/cache_ctrl_logic/n170 ),
    .o(\biu/l1i_bsel [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(440)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux63_b5  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [5]),
    .sel(\biu/cache_ctrl_logic/n170 ),
    .o(\biu/l1i_bsel [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(440)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux63_b6  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [6]),
    .sel(\biu/cache_ctrl_logic/n170 ),
    .o(\biu/l1i_bsel [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(440)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux63_b7  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [7]),
    .sel(\biu/cache_ctrl_logic/n170 ),
    .o(\biu/l1i_bsel [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(440)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux64_b0  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [0]),
    .sel(\biu/cache_ctrl_logic/n171 ),
    .o(\biu/l1d_bsel [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(442)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux64_b1  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [1]),
    .sel(\biu/cache_ctrl_logic/n171 ),
    .o(\biu/l1d_bsel [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(442)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux64_b2  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [2]),
    .sel(\biu/cache_ctrl_logic/n171 ),
    .o(\biu/l1d_bsel [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(442)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux64_b3  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [3]),
    .sel(\biu/cache_ctrl_logic/n171 ),
    .o(\biu/l1d_bsel [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(442)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux64_b4  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [4]),
    .sel(\biu/cache_ctrl_logic/n171 ),
    .o(\biu/l1d_bsel [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(442)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux64_b5  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [5]),
    .sel(\biu/cache_ctrl_logic/n171 ),
    .o(\biu/l1d_bsel [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(442)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux64_b6  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [6]),
    .sel(\biu/cache_ctrl_logic/n171 ),
    .o(\biu/l1d_bsel [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(442)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux64_b7  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/ex_bsel [7]),
    .sel(\biu/cache_ctrl_logic/n171 ),
    .o(\biu/l1d_bsel [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(442)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux65_b0  (
    .i0(ex_priv[0]),
    .i1(priv[0]),
    .sel(\biu/opc [1]),
    .o(\biu/priv [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(499)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux65_b1  (
    .i0(ex_priv[1]),
    .i1(priv[1]),
    .sel(\biu/opc [1]),
    .o(\biu/priv [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(499)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux65_b3  (
    .i0(ex_priv[3]),
    .i1(priv[3]),
    .sel(\biu/opc [1]),
    .o(\biu/priv [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(499)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [0]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [1]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b10  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [10]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b11  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [11]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b12  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [12]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b13  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [13]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b14  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [14]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b15  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [15]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b16  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [16]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b17  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [17]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b18  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [18]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b19  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [19]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b2  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [2]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b20  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [20]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b21  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [21]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b22  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [22]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b23  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [23]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b24  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [24]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b25  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [25]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b26  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [26]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b27  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [27]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b28  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [28]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b29  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [29]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [3]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b30  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [30]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b31  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [31]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b32  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [32]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b33  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [33]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b34  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [34]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b35  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [35]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b36  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [36]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b37  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [37]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b38  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [38]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b39  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [39]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [4]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b40  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [40]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b41  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [41]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b42  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [42]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b43  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [43]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b44  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [44]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b45  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [45]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b46  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [46]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b47  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [47]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b48  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [48]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b49  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [49]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b5  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [5]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b50  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [50]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b51  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [51]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b52  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [52]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b53  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [53]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b54  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [54]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b55  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [55]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b56  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [56]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b57  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [57]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b58  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [58]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b59  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [59]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b6  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [6]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b60  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [60]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b61  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [61]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b62  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [62]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b63  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [63]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b7  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [7]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b8  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [8]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux66_b9  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n207 [9]),
    .sel(\biu/cache_ctrl_logic/n206 ),
    .o(\biu/cache_ctrl_logic/n208 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [0]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [1]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b10  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [10]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b11  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [11]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b12  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [12]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b13  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [13]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b14  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [14]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b15  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [15]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b16  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [16]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b17  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [17]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b18  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [18]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b19  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [19]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b2  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [2]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b20  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [20]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b21  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [21]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b22  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [22]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b23  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [23]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b24  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [24]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b25  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [25]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b26  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [26]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b27  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [27]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b28  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [28]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b29  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [29]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [3]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b30  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [30]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b31  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [31]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b32  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [32]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b33  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [33]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b34  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [34]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b35  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [35]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b36  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [36]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b37  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [37]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b38  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [38]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b39  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [39]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [4]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b40  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [40]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b41  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [41]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b42  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [42]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b43  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [43]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b44  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [44]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b45  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [45]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b46  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [46]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b47  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [47]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b48  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [48]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b49  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [49]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b5  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [5]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b50  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [50]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b51  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [51]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b52  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [52]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b53  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [53]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b54  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [54]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b55  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [55]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b56  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [56]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b57  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [57]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b58  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [58]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b59  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [59]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b6  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [6]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b60  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [60]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b61  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [61]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b62  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [62]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b63  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [63]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b7  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [7]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b8  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [8]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux67_b9  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n209 [9]),
    .sel(\biu/cache_ctrl_logic/n93 ),
    .o(\biu/cache_ctrl_logic/n210 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [0]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [1]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b10  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [10]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b11  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [11]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b12  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [12]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b13  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [13]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b14  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [14]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b15  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [15]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b16  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [16]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b17  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [17]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b18  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [18]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b19  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [19]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b2  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [2]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b20  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [20]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b21  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [21]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b22  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [22]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b23  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [23]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b24  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [24]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b25  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [25]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b26  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [26]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b27  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [27]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b28  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [28]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b29  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [29]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [3]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b30  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [30]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b31  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [31]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b32  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [32]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b33  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [33]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b34  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [34]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b35  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [35]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b36  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [36]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b37  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [37]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b38  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [38]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b39  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [39]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [4]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b40  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [40]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b41  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [41]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b42  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [42]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b43  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [43]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b44  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [44]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b45  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [45]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b46  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [46]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b47  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [47]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b48  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [48]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b49  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [49]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b5  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [5]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b50  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [50]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b51  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [51]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b52  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [52]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b53  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [53]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b54  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [54]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b55  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [55]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b56  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [56]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b57  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [57]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b58  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [58]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b59  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [59]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b6  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [6]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b60  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [60]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b61  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [61]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b62  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [62]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b63  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [63]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b7  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [7]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b8  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [8]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux68_b9  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n212 [9]),
    .sel(\biu/cache_ctrl_logic/n97 ),
    .o(\biu/cache_ctrl_logic/n213 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b0  (
    .i0(1'b0),
    .i1(addr_ex[0]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b1  (
    .i0(1'b0),
    .i1(addr_ex[1]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b10  (
    .i0(1'b0),
    .i1(addr_ex[10]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b11  (
    .i0(1'b0),
    .i1(addr_ex[11]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b12  (
    .i0(1'b0),
    .i1(addr_ex[12]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b13  (
    .i0(1'b0),
    .i1(addr_ex[13]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b14  (
    .i0(1'b0),
    .i1(addr_ex[14]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b15  (
    .i0(1'b0),
    .i1(addr_ex[15]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b16  (
    .i0(1'b0),
    .i1(addr_ex[16]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b17  (
    .i0(1'b0),
    .i1(addr_ex[17]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b18  (
    .i0(1'b0),
    .i1(addr_ex[18]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b19  (
    .i0(1'b0),
    .i1(addr_ex[19]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b2  (
    .i0(1'b0),
    .i1(addr_ex[2]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b20  (
    .i0(1'b0),
    .i1(addr_ex[20]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b21  (
    .i0(1'b0),
    .i1(addr_ex[21]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b22  (
    .i0(1'b0),
    .i1(addr_ex[22]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b23  (
    .i0(1'b0),
    .i1(addr_ex[23]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b24  (
    .i0(1'b0),
    .i1(addr_ex[24]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b25  (
    .i0(1'b0),
    .i1(addr_ex[25]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b26  (
    .i0(1'b0),
    .i1(addr_ex[26]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b27  (
    .i0(1'b0),
    .i1(addr_ex[27]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b28  (
    .i0(1'b0),
    .i1(addr_ex[28]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b29  (
    .i0(1'b0),
    .i1(addr_ex[29]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b3  (
    .i0(1'b0),
    .i1(addr_ex[3]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b30  (
    .i0(1'b0),
    .i1(addr_ex[30]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b31  (
    .i0(1'b0),
    .i1(addr_ex[31]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b32  (
    .i0(1'b0),
    .i1(addr_ex[32]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b33  (
    .i0(1'b0),
    .i1(addr_ex[33]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b34  (
    .i0(1'b0),
    .i1(addr_ex[34]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b35  (
    .i0(1'b0),
    .i1(addr_ex[35]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b36  (
    .i0(1'b0),
    .i1(addr_ex[36]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b37  (
    .i0(1'b0),
    .i1(addr_ex[37]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b38  (
    .i0(1'b0),
    .i1(addr_ex[38]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b39  (
    .i0(1'b0),
    .i1(addr_ex[39]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b4  (
    .i0(1'b0),
    .i1(addr_ex[4]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b40  (
    .i0(1'b0),
    .i1(addr_ex[40]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b41  (
    .i0(1'b0),
    .i1(addr_ex[41]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b42  (
    .i0(1'b0),
    .i1(addr_ex[42]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b43  (
    .i0(1'b0),
    .i1(addr_ex[43]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b44  (
    .i0(1'b0),
    .i1(addr_ex[44]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b45  (
    .i0(1'b0),
    .i1(addr_ex[45]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b46  (
    .i0(1'b0),
    .i1(addr_ex[46]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b47  (
    .i0(1'b0),
    .i1(addr_ex[47]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b48  (
    .i0(1'b0),
    .i1(addr_ex[48]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b49  (
    .i0(1'b0),
    .i1(addr_ex[49]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b5  (
    .i0(1'b0),
    .i1(addr_ex[5]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b50  (
    .i0(1'b0),
    .i1(addr_ex[50]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b51  (
    .i0(1'b0),
    .i1(addr_ex[51]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b52  (
    .i0(1'b0),
    .i1(addr_ex[52]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b53  (
    .i0(1'b0),
    .i1(addr_ex[53]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b54  (
    .i0(1'b0),
    .i1(addr_ex[54]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b55  (
    .i0(1'b0),
    .i1(addr_ex[55]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b56  (
    .i0(1'b0),
    .i1(addr_ex[56]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b57  (
    .i0(1'b0),
    .i1(addr_ex[57]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b58  (
    .i0(1'b0),
    .i1(addr_ex[58]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b59  (
    .i0(1'b0),
    .i1(addr_ex[59]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b6  (
    .i0(1'b0),
    .i1(addr_ex[6]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b60  (
    .i0(1'b0),
    .i1(addr_ex[60]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b61  (
    .i0(1'b0),
    .i1(addr_ex[61]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b62  (
    .i0(1'b0),
    .i1(addr_ex[62]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b63  (
    .i0(1'b0),
    .i1(addr_ex[63]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b7  (
    .i0(1'b0),
    .i1(addr_ex[7]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b8  (
    .i0(1'b0),
    .i1(addr_ex[8]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux69_b9  (
    .i0(1'b0),
    .i1(addr_ex[9]),
    .sel(\biu/cache_ctrl_logic/n75 ),
    .o(\biu/cache_ctrl_logic/n215 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux6_b0  (
    .i0(\biu/cache_ctrl_logic/n82 [0]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n77 ),
    .o(\biu/cache_ctrl_logic/n83 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  and \biu/cache_ctrl_logic/mux6_b2_sel_is_0  (\biu/cache_ctrl_logic/mux6_b2_sel_is_0_o , \biu/cache_ctrl_logic/n77_neg , \biu/cache_ctrl_logic/n68_neg );
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b0  (
    .i0(1'b0),
    .i1(addr_if[0]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b1  (
    .i0(1'b0),
    .i1(addr_if[1]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b10  (
    .i0(1'b0),
    .i1(addr_if[10]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b11  (
    .i0(1'b0),
    .i1(addr_if[11]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b12  (
    .i0(1'b0),
    .i1(addr_if[12]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b13  (
    .i0(1'b0),
    .i1(addr_if[13]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b14  (
    .i0(1'b0),
    .i1(addr_if[14]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b15  (
    .i0(1'b0),
    .i1(addr_if[15]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b16  (
    .i0(1'b0),
    .i1(addr_if[16]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b17  (
    .i0(1'b0),
    .i1(addr_if[17]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b18  (
    .i0(1'b0),
    .i1(addr_if[18]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b19  (
    .i0(1'b0),
    .i1(addr_if[19]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b2  (
    .i0(1'b0),
    .i1(addr_if[2]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b20  (
    .i0(1'b0),
    .i1(addr_if[20]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b21  (
    .i0(1'b0),
    .i1(addr_if[21]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b22  (
    .i0(1'b0),
    .i1(addr_if[22]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b23  (
    .i0(1'b0),
    .i1(addr_if[23]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b24  (
    .i0(1'b0),
    .i1(addr_if[24]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b25  (
    .i0(1'b0),
    .i1(addr_if[25]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b26  (
    .i0(1'b0),
    .i1(addr_if[26]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b27  (
    .i0(1'b0),
    .i1(addr_if[27]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b28  (
    .i0(1'b0),
    .i1(addr_if[28]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b29  (
    .i0(1'b0),
    .i1(addr_if[29]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b3  (
    .i0(1'b0),
    .i1(addr_if[3]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b30  (
    .i0(1'b0),
    .i1(addr_if[30]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b31  (
    .i0(1'b0),
    .i1(addr_if[31]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b32  (
    .i0(1'b0),
    .i1(addr_if[32]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b33  (
    .i0(1'b0),
    .i1(addr_if[33]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b34  (
    .i0(1'b0),
    .i1(addr_if[34]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b35  (
    .i0(1'b0),
    .i1(addr_if[35]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b36  (
    .i0(1'b0),
    .i1(addr_if[36]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b37  (
    .i0(1'b0),
    .i1(addr_if[37]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b38  (
    .i0(1'b0),
    .i1(addr_if[38]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b39  (
    .i0(1'b0),
    .i1(addr_if[39]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b4  (
    .i0(1'b0),
    .i1(addr_if[4]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b40  (
    .i0(1'b0),
    .i1(addr_if[40]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b41  (
    .i0(1'b0),
    .i1(addr_if[41]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b42  (
    .i0(1'b0),
    .i1(addr_if[42]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b43  (
    .i0(1'b0),
    .i1(addr_if[43]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b44  (
    .i0(1'b0),
    .i1(addr_if[44]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b45  (
    .i0(1'b0),
    .i1(addr_if[45]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b46  (
    .i0(1'b0),
    .i1(addr_if[46]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b47  (
    .i0(1'b0),
    .i1(addr_if[47]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b48  (
    .i0(1'b0),
    .i1(addr_if[48]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b49  (
    .i0(1'b0),
    .i1(addr_if[49]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b5  (
    .i0(1'b0),
    .i1(addr_if[5]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b50  (
    .i0(1'b0),
    .i1(addr_if[50]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b51  (
    .i0(1'b0),
    .i1(addr_if[51]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b52  (
    .i0(1'b0),
    .i1(addr_if[52]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b53  (
    .i0(1'b0),
    .i1(addr_if[53]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b54  (
    .i0(1'b0),
    .i1(addr_if[54]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b55  (
    .i0(1'b0),
    .i1(addr_if[55]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b56  (
    .i0(1'b0),
    .i1(addr_if[56]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b57  (
    .i0(1'b0),
    .i1(addr_if[57]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b58  (
    .i0(1'b0),
    .i1(addr_if[58]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b59  (
    .i0(1'b0),
    .i1(addr_if[59]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b6  (
    .i0(1'b0),
    .i1(addr_if[6]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b60  (
    .i0(1'b0),
    .i1(addr_if[60]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b61  (
    .i0(1'b0),
    .i1(addr_if[61]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b62  (
    .i0(1'b0),
    .i1(addr_if[62]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b63  (
    .i0(1'b0),
    .i1(addr_if[63]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b7  (
    .i0(1'b0),
    .i1(addr_if[7]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b8  (
    .i0(1'b0),
    .i1(addr_if[8]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux70_b9  (
    .i0(1'b0),
    .i1(addr_if[9]),
    .sel(\biu/opc [1]),
    .o(\biu/cache_ctrl_logic/n217 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [64]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [65]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b10  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [74]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b11  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [75]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b12  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [76]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b13  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [77]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b14  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [78]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b15  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [79]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b16  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [80]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b17  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [81]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b18  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [82]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b19  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [83]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b2  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [66]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b20  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [84]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b21  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [85]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b22  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [86]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b23  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [87]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b24  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [88]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b25  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [89]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b26  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [90]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b27  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [91]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b28  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [92]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b29  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [93]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [67]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b30  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [94]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b31  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [95]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b32  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [96]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b33  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [97]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b34  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [98]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b35  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [99]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b36  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [100]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b37  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [101]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b38  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [102]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b39  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [103]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [68]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b40  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [104]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b41  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [105]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b42  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [106]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b43  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [107]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b44  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [108]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b45  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [109]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b46  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [110]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b47  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [111]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b48  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [112]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b49  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [113]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b5  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [69]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b50  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [114]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b51  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [115]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b52  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [116]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b53  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [117]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b54  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [118]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b55  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [119]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b56  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [120]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b57  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [121]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b58  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [122]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b59  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [123]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b6  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [70]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b60  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [124]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b61  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [125]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b62  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [126]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b63  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [127]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b7  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [71]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b8  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [72]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux71_b9  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pa [73]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n219 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [64]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [65]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b10  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [74]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b11  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [75]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b12  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [76]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b13  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [77]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b14  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [78]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b15  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [79]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b16  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [80]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b17  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [81]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b18  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [82]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b19  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [83]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b2  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [66]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b20  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [84]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b21  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [85]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b22  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [86]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b23  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [87]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b24  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [88]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b25  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [89]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b26  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [90]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b27  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [91]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b28  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [92]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b29  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [93]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [67]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b30  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [94]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b31  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [95]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b32  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [96]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b33  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [97]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b34  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [98]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b35  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [99]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b36  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [100]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b37  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [101]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b38  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [102]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b39  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [103]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [68]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b40  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [104]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b41  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [105]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b42  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [106]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b43  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [107]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b44  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [108]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b45  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [109]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b46  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [110]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b47  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [111]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b48  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [112]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b49  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [113]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b5  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [69]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b50  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [114]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b51  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [115]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b52  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [116]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b53  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [117]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b54  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [118]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b55  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [119]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b56  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [120]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b57  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [121]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b58  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [122]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b59  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [123]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b6  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [70]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b60  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [124]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b61  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [125]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b62  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [126]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b63  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [127]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b7  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [71]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b8  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [72]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux72_b9  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pa [73]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n221 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [64]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [65]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b10  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [74]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b11  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [75]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b12  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [76]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b13  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [77]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b14  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [78]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b15  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [79]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b16  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [80]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b17  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [81]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b18  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [82]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b19  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [83]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b2  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [66]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b20  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [84]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b21  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [85]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b22  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [86]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b23  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [87]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b24  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [88]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b25  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [89]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b26  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [90]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b27  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [91]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b28  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [92]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b29  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [93]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [67]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b30  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [94]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b31  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [95]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b32  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [96]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b33  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [97]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b34  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [98]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b35  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [99]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b36  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [100]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b37  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [101]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b38  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [102]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b39  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [103]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [68]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b40  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [104]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b41  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [105]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b42  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [106]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b43  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [107]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b44  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [108]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b45  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [109]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b46  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [110]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b47  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [111]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b48  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [112]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b49  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [113]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b5  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [69]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b50  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [114]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b51  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [115]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b52  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [116]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b53  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [117]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b54  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [118]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b55  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [119]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b56  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [120]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b57  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [121]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b58  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [122]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b59  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [123]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b6  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [70]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b60  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [124]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b61  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [125]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b62  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [126]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b63  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [127]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b7  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [71]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b8  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [72]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux73_b9  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pa_temp [73]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n223 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b0  (
    .i0(1'b0),
    .i1(addr_ex[0]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b1  (
    .i0(1'b0),
    .i1(addr_ex[1]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b10  (
    .i0(1'b0),
    .i1(addr_ex[10]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b11  (
    .i0(1'b0),
    .i1(addr_ex[11]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b2  (
    .i0(1'b0),
    .i1(addr_ex[2]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b3  (
    .i0(1'b0),
    .i1(addr_ex[3]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b4  (
    .i0(1'b0),
    .i1(addr_ex[4]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b5  (
    .i0(1'b0),
    .i1(addr_ex[5]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b6  (
    .i0(1'b0),
    .i1(addr_ex[6]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b7  (
    .i0(1'b0),
    .i1(addr_ex[7]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b8  (
    .i0(1'b0),
    .i1(addr_ex[8]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux74_b9  (
    .i0(1'b0),
    .i1(addr_ex[9]),
    .sel(\biu/cache_ctrl_logic/n225 ),
    .o(\biu/cache_ctrl_logic/off [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b0  (
    .i0(1'b0),
    .i1(\exu/lsu/n1 [0]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b1  (
    .i0(1'b0),
    .i1(\exu/lsu/n1 [1]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b10  (
    .i0(1'b0),
    .i1(\exu/lsu/n4 [10]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b11  (
    .i0(1'b0),
    .i1(\exu/lsu/n4 [11]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b12  (
    .i0(1'b0),
    .i1(\exu/lsu/n4 [12]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b13  (
    .i0(1'b0),
    .i1(\exu/lsu/n4 [13]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b14  (
    .i0(1'b0),
    .i1(\exu/lsu/n4 [14]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b15  (
    .i0(1'b0),
    .i1(\exu/lsu/n4 [15]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b16  (
    .i0(1'b0),
    .i1(\exu/lsu/n7 [16]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b17  (
    .i0(1'b0),
    .i1(\exu/lsu/n7 [17]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b18  (
    .i0(1'b0),
    .i1(\exu/lsu/n7 [18]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b19  (
    .i0(1'b0),
    .i1(\exu/lsu/n7 [19]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b2  (
    .i0(1'b0),
    .i1(\exu/lsu/n1 [2]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b20  (
    .i0(1'b0),
    .i1(\exu/lsu/n7 [20]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b21  (
    .i0(1'b0),
    .i1(\exu/lsu/n7 [21]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b22  (
    .i0(1'b0),
    .i1(\exu/lsu/n7 [22]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b23  (
    .i0(1'b0),
    .i1(\exu/lsu/n7 [23]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b24  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [24]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b25  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [25]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b26  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [26]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b27  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [27]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b28  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [28]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b29  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [29]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b3  (
    .i0(1'b0),
    .i1(\exu/lsu/n1 [3]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b30  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [30]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b31  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [31]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b32  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [32]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b33  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [33]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b34  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [34]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b35  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [35]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b36  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [36]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b37  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [37]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b38  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [38]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b39  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [39]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b4  (
    .i0(1'b0),
    .i1(\exu/lsu/n1 [4]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b40  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [40]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b41  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [41]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b42  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [42]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b43  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [43]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b44  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [44]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b45  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [45]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b46  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [46]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b47  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [47]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b48  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [48]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b49  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [49]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b5  (
    .i0(1'b0),
    .i1(\exu/lsu/n1 [5]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b50  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [50]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b51  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [51]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b52  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [52]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b53  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [53]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b54  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [54]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b55  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [55]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b56  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [56]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b57  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [57]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b58  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [58]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b59  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [59]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b6  (
    .i0(1'b0),
    .i1(\exu/lsu/n1 [6]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b60  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [60]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b61  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [61]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b62  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [62]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b63  (
    .i0(1'b0),
    .i1(\exu/lsu/n10 [63]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b7  (
    .i0(1'b0),
    .i1(\exu/lsu/n1 [7]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b8  (
    .i0(1'b0),
    .i1(\exu/lsu/n4 [8]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux75_b9  (
    .i0(1'b0),
    .i1(\exu/lsu/n4 [9]),
    .sel(\biu/cache_ctrl_logic/n227 ),
    .o(\biu/cache_ctrl_logic/n228 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [0]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [1]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b10  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [10]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b11  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [11]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b12  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [12]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b13  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [13]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b14  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [14]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b15  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [15]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b16  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [16]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b17  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [17]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b18  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [18]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b19  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [19]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b2  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [2]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b20  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [20]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b21  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [21]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b22  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [22]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b23  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [23]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b24  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [24]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b25  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [25]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b26  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [26]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b27  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [27]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b28  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [28]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b29  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [29]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [3]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b30  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [30]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b31  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [31]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b32  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [32]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b33  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [33]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b34  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [34]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b35  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [35]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b36  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [36]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b37  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [37]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b38  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [38]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b39  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [39]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [4]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b40  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [40]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b41  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [41]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b42  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [42]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b43  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [43]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b44  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [44]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b45  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [45]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b46  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [46]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b47  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [47]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b48  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [48]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b49  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [49]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b5  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [5]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b50  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [50]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b51  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [51]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b52  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [52]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b53  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [53]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b54  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [54]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b55  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [55]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b56  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [56]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b57  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [57]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b58  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [58]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b59  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [59]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b6  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [6]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b60  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [60]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b61  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [61]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b62  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [62]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b63  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [63]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b7  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [7]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b8  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [8]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux76_b9  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/pte_temp [9]),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n229 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [0]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [1]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b10  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [10]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b11  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [11]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b12  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [12]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b13  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [13]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b14  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [14]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b15  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [15]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b16  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [16]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b17  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [17]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b18  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [18]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b19  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [19]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b2  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [2]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b20  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [20]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b21  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [21]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b22  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [22]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b23  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [23]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b24  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [24]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b25  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [25]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b26  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [26]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b27  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [27]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b28  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [28]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b29  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [29]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [3]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b30  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [30]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b31  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [31]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b32  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [32]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b33  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [33]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b34  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [34]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b35  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [35]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b36  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [36]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b37  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [37]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b38  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [38]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b39  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [39]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [4]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b40  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [40]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b41  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [41]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b42  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [42]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b43  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [43]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b44  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [44]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b45  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [45]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b46  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [46]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b47  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [47]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b48  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [48]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b49  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [49]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b5  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [5]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b50  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [50]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b51  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [51]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b52  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [52]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b53  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [53]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b54  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [54]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b55  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [55]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b56  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [56]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b57  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [57]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b58  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [58]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b59  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [59]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b6  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [6]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b60  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [60]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b61  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [61]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b62  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [62]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b63  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [63]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b7  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [7]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b8  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [8]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux77_b9  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1i_pte [9]),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n231 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b0  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [0]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b1  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [1]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b10  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [10]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b11  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [11]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b12  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [12]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b13  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [13]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b14  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [14]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b15  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [15]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b16  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [16]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b17  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [17]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b18  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [18]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b19  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [19]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b2  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [2]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b20  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [20]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b21  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [21]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b22  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [22]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b23  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [23]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b24  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [24]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b25  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [25]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b26  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [26]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b27  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [27]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b28  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [28]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b29  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [29]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [3]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b30  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [30]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b31  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [31]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b32  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [32]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b33  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [33]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b34  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [34]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b35  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [35]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b36  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [36]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b37  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [37]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b38  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [38]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b39  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [39]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b4  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [4]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b40  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [40]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b41  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [41]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b42  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [42]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b43  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [43]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b44  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [44]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b45  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [45]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b46  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [46]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b47  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [47]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b48  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [48]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b49  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [49]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b5  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [5]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b50  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [50]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b51  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [51]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b52  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [52]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b53  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [53]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b54  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [54]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b55  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [55]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b56  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [56]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b57  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [57]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b58  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [58]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b59  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [59]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b6  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [6]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b60  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [60]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b61  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [61]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b62  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [62]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b63  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [63]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b7  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [7]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b8  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [8]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux78_b9  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/l1d_pte [9]),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n233 [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux7_b0  (
    .i0(\biu/cache_ctrl_logic/n83 [0]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n76 ),
    .o(\biu/cache_ctrl_logic/n84 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  AL_MUX \biu/cache_ctrl_logic/mux7_b1  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/mux7_b1_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n84 [1]));
  and \biu/cache_ctrl_logic/mux7_b1_sel_is_0  (\biu/cache_ctrl_logic/mux7_b1_sel_is_0_o , \biu/cache_ctrl_logic/n76_neg , \biu/cache_ctrl_logic/n77_neg );
  AL_MUX \biu/cache_ctrl_logic/mux7_b2  (
    .i0(1'b1),
    .i1(\biu/cache_ctrl_logic/n81 [2]),
    .sel(\biu/cache_ctrl_logic/mux7_b2_sel_is_2_o ),
    .o(\biu/cache_ctrl_logic/n84 [2]));
  and \biu/cache_ctrl_logic/mux7_b2_sel_is_2  (\biu/cache_ctrl_logic/mux7_b2_sel_is_2_o , \biu/cache_ctrl_logic/n76_neg , \biu/cache_ctrl_logic/mux6_b2_sel_is_0_o );
  AL_MUX \biu/cache_ctrl_logic/mux7_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n81 [3]),
    .sel(\biu/cache_ctrl_logic/mux7_b2_sel_is_2_o ),
    .o(\biu/cache_ctrl_logic/n84 [3]));
  AL_MUX \biu/cache_ctrl_logic/mux7_b4  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/mux7_b1_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n84 [4]));
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux8_b0  (
    .i0(\biu/cache_ctrl_logic/n73 [2]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n86 ),
    .o(\biu/cache_ctrl_logic/n87 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(264)
  binary_mux_s1_w1 \biu/cache_ctrl_logic/mux9_b0  (
    .i0(\biu/cache_ctrl_logic/n87 [0]),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/n85 ),
    .o(\biu/cache_ctrl_logic/n88 [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(264)
  AL_MUX \biu/cache_ctrl_logic/mux9_b2  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\biu/cache_ctrl_logic/mux9_b2_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n88 [2]));
  and \biu/cache_ctrl_logic/mux9_b2_sel_is_0  (\biu/cache_ctrl_logic/mux9_b2_sel_is_0_o , \biu/cache_ctrl_logic/n85_neg , \biu/cache_ctrl_logic/n86_neg );
  AL_MUX \biu/cache_ctrl_logic/mux9_b3  (
    .i0(1'b0),
    .i1(\biu/cache_ctrl_logic/n73 [2]),
    .sel(\biu/cache_ctrl_logic/mux9_b2_sel_is_0_o ),
    .o(\biu/cache_ctrl_logic/n88 [3]));
  not \biu/cache_ctrl_logic/n102_inv  (\biu/cache_ctrl_logic/n102_neg , \biu/cache_ctrl_logic/n102 );
  not \biu/cache_ctrl_logic/n104_inv  (\biu/cache_ctrl_logic/n104_neg , \biu/cache_ctrl_logic/n104 );
  not \biu/cache_ctrl_logic/n106_inv  (\biu/cache_ctrl_logic/n106_neg , \biu/cache_ctrl_logic/n106 );
  not \biu/cache_ctrl_logic/n107_inv  (\biu/cache_ctrl_logic/n107_neg , \biu/cache_ctrl_logic/n107 );
  not \biu/cache_ctrl_logic/n108_inv  (\biu/cache_ctrl_logic/n108_neg , \biu/cache_ctrl_logic/n108 );
  not \biu/cache_ctrl_logic/n161_inv  (\biu/cache_ctrl_logic/n161_neg , \biu/cache_ctrl_logic/n161 );
  not \biu/cache_ctrl_logic/n56_inv  (\biu/cache_ctrl_logic/n56_neg , \biu/cache_ctrl_logic/n56 );
  not \biu/cache_ctrl_logic/n57_inv  (\biu/cache_ctrl_logic/n57_neg , \biu/cache_ctrl_logic/n57 );
  not \biu/cache_ctrl_logic/n62_inv  (\biu/cache_ctrl_logic/n62_neg , \biu/cache_ctrl_logic/n62 );
  not \biu/cache_ctrl_logic/n63_inv  (\biu/cache_ctrl_logic/n63_neg , \biu/cache_ctrl_logic/n63 );
  not \biu/cache_ctrl_logic/n64_inv  (\biu/cache_ctrl_logic/n64_neg , \biu/cache_ctrl_logic/n64 );
  not \biu/cache_ctrl_logic/n65_inv  (\biu/cache_ctrl_logic/n65_neg , \biu/cache_ctrl_logic/n65 );
  not \biu/cache_ctrl_logic/n66_inv  (\biu/cache_ctrl_logic/n66_neg , \biu/cache_ctrl_logic/n66 );
  not \biu/cache_ctrl_logic/n67_inv  (\biu/cache_ctrl_logic/n67_neg , \biu/cache_ctrl_logic/n67 );
  not \biu/cache_ctrl_logic/n68_inv  (\biu/cache_ctrl_logic/n68_neg , \biu/cache_ctrl_logic/n68 );
  not \biu/cache_ctrl_logic/n76_inv  (\biu/cache_ctrl_logic/n76_neg , \biu/cache_ctrl_logic/n76 );
  not \biu/cache_ctrl_logic/n77_inv  (\biu/cache_ctrl_logic/n77_neg , \biu/cache_ctrl_logic/n77 );
  not \biu/cache_ctrl_logic/n85_inv  (\biu/cache_ctrl_logic/n85_neg , \biu/cache_ctrl_logic/n85 );
  not \biu/cache_ctrl_logic/n86_inv  (\biu/cache_ctrl_logic/n86_neg , \biu/cache_ctrl_logic/n86 );
  not \biu/cache_ctrl_logic/n89_inv  (\biu/cache_ctrl_logic/n89_neg , \biu/cache_ctrl_logic/n89 );
  not \biu/cache_ctrl_logic/n93_inv  (\biu/cache_ctrl_logic/n93_neg , \biu/cache_ctrl_logic/n93 );
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b12  (
    .clk(clk),
    .d(addr_if[12]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b13  (
    .clk(clk),
    .d(addr_if[13]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b14  (
    .clk(clk),
    .d(addr_if[14]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b15  (
    .clk(clk),
    .d(addr_if[15]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b16  (
    .clk(clk),
    .d(addr_if[16]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b17  (
    .clk(clk),
    .d(addr_if[17]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b18  (
    .clk(clk),
    .d(addr_if[18]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b19  (
    .clk(clk),
    .d(addr_if[19]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b20  (
    .clk(clk),
    .d(addr_if[20]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b21  (
    .clk(clk),
    .d(addr_if[21]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b22  (
    .clk(clk),
    .d(addr_if[22]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b23  (
    .clk(clk),
    .d(addr_if[23]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b24  (
    .clk(clk),
    .d(addr_if[24]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b25  (
    .clk(clk),
    .d(addr_if[25]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b26  (
    .clk(clk),
    .d(addr_if[26]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b27  (
    .clk(clk),
    .d(addr_if[27]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b28  (
    .clk(clk),
    .d(addr_if[28]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b29  (
    .clk(clk),
    .d(addr_if[29]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b30  (
    .clk(clk),
    .d(addr_if[30]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b31  (
    .clk(clk),
    .d(addr_if[31]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b32  (
    .clk(clk),
    .d(addr_if[32]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b33  (
    .clk(clk),
    .d(addr_if[33]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b34  (
    .clk(clk),
    .d(addr_if[34]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b35  (
    .clk(clk),
    .d(addr_if[35]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b36  (
    .clk(clk),
    .d(addr_if[36]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b37  (
    .clk(clk),
    .d(addr_if[37]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b38  (
    .clk(clk),
    .d(addr_if[38]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b39  (
    .clk(clk),
    .d(addr_if[39]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b40  (
    .clk(clk),
    .d(addr_if[40]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b41  (
    .clk(clk),
    .d(addr_if[41]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b42  (
    .clk(clk),
    .d(addr_if[42]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b43  (
    .clk(clk),
    .d(addr_if[43]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b44  (
    .clk(clk),
    .d(addr_if[44]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b45  (
    .clk(clk),
    .d(addr_if[45]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b46  (
    .clk(clk),
    .d(addr_if[46]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b47  (
    .clk(clk),
    .d(addr_if[47]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b48  (
    .clk(clk),
    .d(addr_if[48]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b49  (
    .clk(clk),
    .d(addr_if[49]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b50  (
    .clk(clk),
    .d(addr_if[50]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b51  (
    .clk(clk),
    .d(addr_if[51]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b52  (
    .clk(clk),
    .d(addr_if[52]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b53  (
    .clk(clk),
    .d(addr_if[53]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b54  (
    .clk(clk),
    .d(addr_if[54]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b55  (
    .clk(clk),
    .d(addr_if[55]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b56  (
    .clk(clk),
    .d(addr_if[56]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b57  (
    .clk(clk),
    .d(addr_if[57]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b58  (
    .clk(clk),
    .d(addr_if[58]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b59  (
    .clk(clk),
    .d(addr_if[59]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b60  (
    .clk(clk),
    .d(addr_if[60]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b61  (
    .clk(clk),
    .d(addr_if[61]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b62  (
    .clk(clk),
    .d(addr_if[62]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg0_b63  (
    .clk(clk),
    .d(addr_if[63]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_va [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(323)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b0  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [0]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b1  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [1]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b10  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [10]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b100  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [100]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [100]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b101  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [101]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [101]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b102  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [102]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [102]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b103  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [103]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [103]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b104  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [104]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [104]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b105  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [105]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [105]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b106  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [106]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [106]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b107  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [107]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [107]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b108  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [108]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [108]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b109  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [109]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [109]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b11  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [11]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b110  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [110]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [110]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b111  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [111]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [111]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b112  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [112]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [112]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b113  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [113]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [113]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b114  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [114]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [114]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b115  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [115]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [115]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b116  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [116]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [116]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b117  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [117]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [117]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b118  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [118]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [118]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b119  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [119]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [119]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b12  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [12]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b120  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [120]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [120]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b121  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [121]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [121]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b122  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [122]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [122]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b123  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [123]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [123]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b124  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [124]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [124]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b125  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [125]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [125]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b126  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [126]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [126]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b127  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [127]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [127]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b13  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [13]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b14  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [14]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b15  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [15]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b16  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [16]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b17  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [17]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b18  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [18]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b19  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [19]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b2  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [2]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b20  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [20]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b21  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [21]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b22  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [22]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b23  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [23]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b24  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [24]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b25  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [25]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b26  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [26]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b27  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [27]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b28  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [28]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b29  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [29]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b3  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [3]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b30  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [30]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b31  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [31]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b32  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [32]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b33  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [33]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b34  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [34]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b35  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [35]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b36  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [36]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b37  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [37]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b38  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [38]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b39  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [39]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b4  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [4]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b40  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [40]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b41  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [41]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b42  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [42]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b43  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [43]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b44  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [44]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b45  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [45]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b46  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [46]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b47  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [47]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b48  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [48]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b49  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [49]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b5  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [5]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b50  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [50]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b51  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [51]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b52  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [52]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b53  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [53]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b54  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [54]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b55  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [55]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b56  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [56]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b57  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [57]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b58  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [58]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b59  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [59]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b6  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [6]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b60  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [60]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b61  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [61]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b62  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [62]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b63  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [63]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b64  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [64]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [64]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b65  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [65]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [65]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b66  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [66]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [66]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b67  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [67]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [67]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b68  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [68]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [68]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b69  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [69]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [69]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b7  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [7]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b70  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [70]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [70]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b71  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [71]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [71]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b72  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [72]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [72]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b73  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [73]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [73]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b74  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [74]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [74]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b75  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [75]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [75]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b76  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [76]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [76]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b77  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [77]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [77]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b78  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [78]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [78]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b79  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [79]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [79]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b8  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [8]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b80  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [80]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [80]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b81  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [81]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [81]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b82  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [82]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [82]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b83  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [83]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [83]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b84  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [84]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [84]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b85  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [85]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [85]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b86  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [86]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [86]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b87  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [87]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [87]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b88  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [88]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [88]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b89  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [89]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [89]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b9  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [9]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b90  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [90]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [90]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b91  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [91]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [91]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b92  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [92]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [92]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b93  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [93]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [93]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b94  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [94]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [94]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b95  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [95]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [95]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b96  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [96]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [96]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b97  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [97]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [97]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b98  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [98]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [98]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg1_b99  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [99]),
    .en(\biu/cache_ctrl_logic/n140 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pa [99]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(333)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b0  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [0]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b1  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [1]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b10  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [10]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b11  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [11]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b12  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [12]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b13  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [13]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b14  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [14]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b15  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [15]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b16  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [16]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b17  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [17]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b18  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [18]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b19  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [19]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b2  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [2]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b20  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [20]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b21  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [21]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b22  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [22]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b23  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [23]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b24  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [24]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b25  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [25]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b26  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [26]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b27  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [27]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b28  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [28]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b29  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [29]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b3  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [3]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b30  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [30]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b31  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [31]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b32  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [32]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b33  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [33]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b34  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [34]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b35  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [35]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b36  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [36]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b37  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [37]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b38  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [38]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b39  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [39]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b4  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [4]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b40  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [40]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b41  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [41]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b42  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [42]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b43  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [43]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b44  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [44]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b45  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [45]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b46  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [46]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b47  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [47]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b48  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [48]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b49  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [49]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b5  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [5]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b50  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [50]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b51  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [51]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b52  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [52]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b53  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [53]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b54  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [54]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b55  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [55]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b56  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [56]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b57  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [57]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b58  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [58]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b59  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [59]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b6  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [6]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b60  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [60]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b61  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [61]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b62  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [62]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b63  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [63]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b7  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n147 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b8  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [8]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg2_b9  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [9]),
    .en(\biu/cache_ctrl_logic/n135 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1i_pte [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(362)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b12  (
    .clk(clk),
    .d(addr_ex[12]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b13  (
    .clk(clk),
    .d(addr_ex[13]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b14  (
    .clk(clk),
    .d(addr_ex[14]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b15  (
    .clk(clk),
    .d(addr_ex[15]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b16  (
    .clk(clk),
    .d(addr_ex[16]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b17  (
    .clk(clk),
    .d(addr_ex[17]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b18  (
    .clk(clk),
    .d(addr_ex[18]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b19  (
    .clk(clk),
    .d(addr_ex[19]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b20  (
    .clk(clk),
    .d(addr_ex[20]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b21  (
    .clk(clk),
    .d(addr_ex[21]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b22  (
    .clk(clk),
    .d(addr_ex[22]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b23  (
    .clk(clk),
    .d(addr_ex[23]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b24  (
    .clk(clk),
    .d(addr_ex[24]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b25  (
    .clk(clk),
    .d(addr_ex[25]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b26  (
    .clk(clk),
    .d(addr_ex[26]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b27  (
    .clk(clk),
    .d(addr_ex[27]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b28  (
    .clk(clk),
    .d(addr_ex[28]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b29  (
    .clk(clk),
    .d(addr_ex[29]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b30  (
    .clk(clk),
    .d(addr_ex[30]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b31  (
    .clk(clk),
    .d(addr_ex[31]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b32  (
    .clk(clk),
    .d(addr_ex[32]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b33  (
    .clk(clk),
    .d(addr_ex[33]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b34  (
    .clk(clk),
    .d(addr_ex[34]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b35  (
    .clk(clk),
    .d(addr_ex[35]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b36  (
    .clk(clk),
    .d(addr_ex[36]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b37  (
    .clk(clk),
    .d(addr_ex[37]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b38  (
    .clk(clk),
    .d(addr_ex[38]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b39  (
    .clk(clk),
    .d(addr_ex[39]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b40  (
    .clk(clk),
    .d(addr_ex[40]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b41  (
    .clk(clk),
    .d(addr_ex[41]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b42  (
    .clk(clk),
    .d(addr_ex[42]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b43  (
    .clk(clk),
    .d(addr_ex[43]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b44  (
    .clk(clk),
    .d(addr_ex[44]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b45  (
    .clk(clk),
    .d(addr_ex[45]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b46  (
    .clk(clk),
    .d(addr_ex[46]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b47  (
    .clk(clk),
    .d(addr_ex[47]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b48  (
    .clk(clk),
    .d(addr_ex[48]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b49  (
    .clk(clk),
    .d(addr_ex[49]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b50  (
    .clk(clk),
    .d(addr_ex[50]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b51  (
    .clk(clk),
    .d(addr_ex[51]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b52  (
    .clk(clk),
    .d(addr_ex[52]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b53  (
    .clk(clk),
    .d(addr_ex[53]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b54  (
    .clk(clk),
    .d(addr_ex[54]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b55  (
    .clk(clk),
    .d(addr_ex[55]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b56  (
    .clk(clk),
    .d(addr_ex[56]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b57  (
    .clk(clk),
    .d(addr_ex[57]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b58  (
    .clk(clk),
    .d(addr_ex[58]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b59  (
    .clk(clk),
    .d(addr_ex[59]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b60  (
    .clk(clk),
    .d(addr_ex[60]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b61  (
    .clk(clk),
    .d(addr_ex[61]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b62  (
    .clk(clk),
    .d(addr_ex[62]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg3_b63  (
    .clk(clk),
    .d(addr_ex[63]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_va [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(372)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b0  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [0]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b1  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [1]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b10  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [10]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b100  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [100]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [100]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b101  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [101]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [101]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b102  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [102]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [102]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b103  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [103]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [103]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b104  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [104]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [104]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b105  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [105]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [105]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b106  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [106]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [106]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b107  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [107]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [107]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b108  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [108]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [108]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b109  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [109]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [109]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b11  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [11]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b110  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [110]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [110]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b111  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [111]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [111]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b112  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [112]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [112]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b113  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [113]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [113]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b114  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [114]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [114]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b115  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [115]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [115]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b116  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [116]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [116]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b117  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [117]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [117]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b118  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [118]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [118]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b119  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [119]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [119]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b12  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [12]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b120  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [120]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [120]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b121  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [121]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [121]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b122  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [122]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [122]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b123  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [123]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [123]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b124  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [124]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [124]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b125  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [125]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [125]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b126  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [126]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [126]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b127  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [127]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [127]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b13  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [13]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b14  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [14]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b15  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [15]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b16  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [16]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b17  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [17]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b18  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [18]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b19  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [19]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b2  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [2]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b20  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [20]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b21  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [21]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b22  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [22]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b23  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [23]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b24  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [24]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b25  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [25]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b26  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [26]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b27  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [27]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b28  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [28]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b29  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [29]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b3  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [3]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b30  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [30]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b31  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [31]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b32  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [32]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b33  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [33]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b34  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [34]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b35  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [35]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b36  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [36]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b37  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [37]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b38  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [38]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b39  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [39]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b4  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [4]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b40  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [40]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b41  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [41]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b42  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [42]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b43  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [43]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b44  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [44]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b45  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [45]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b46  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [46]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b47  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [47]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b48  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [48]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b49  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [49]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b5  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [5]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b50  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [50]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b51  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [51]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b52  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [52]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b53  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [53]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b54  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [54]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b55  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [55]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b56  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [56]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b57  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [57]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b58  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [58]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b59  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [59]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b6  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [6]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b60  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [60]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b61  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [61]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b62  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [62]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b63  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [63]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b64  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [64]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [64]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b65  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [65]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [65]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b66  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [66]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [66]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b67  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [67]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [67]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b68  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [68]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [68]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b69  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [69]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [69]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b7  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [7]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b70  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [70]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [70]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b71  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [71]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [71]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b72  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [72]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [72]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b73  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [73]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [73]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b74  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [74]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [74]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b75  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [75]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [75]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b76  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [76]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [76]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b77  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [77]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [77]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b78  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [78]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [78]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b79  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [79]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [79]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b8  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [8]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b80  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [80]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [80]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b81  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [81]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [81]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b82  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [82]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [82]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b83  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [83]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [83]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b84  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [84]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [84]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b85  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [85]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [85]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b86  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [86]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [86]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b87  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [87]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [87]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b88  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [88]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [88]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b89  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [89]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [89]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b9  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [9]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b90  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [90]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [90]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b91  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [91]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [91]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b92  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [92]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [92]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b93  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [93]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [93]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b94  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [94]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [94]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b95  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [95]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [95]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b96  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [96]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [96]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b97  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [97]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [97]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b98  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [98]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [98]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg4_b99  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pa_temp [99]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pa [99]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(382)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b0  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [0]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b1  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [1]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b10  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [10]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b11  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [11]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b12  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [12]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b13  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [13]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b14  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [14]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b15  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [15]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b16  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [16]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b17  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [17]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b18  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [18]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b19  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [19]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b2  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [2]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b20  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [20]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b21  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [21]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b22  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [22]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b23  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [23]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b24  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [24]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b25  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [25]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b26  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [26]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b27  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [27]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b28  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [28]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b29  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [29]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b3  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [3]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b30  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [30]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b31  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [31]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b32  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [32]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b33  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [33]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b34  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [34]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b35  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [35]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b36  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [36]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b37  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [37]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b38  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [38]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b39  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [39]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b4  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [4]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b40  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [40]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b41  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [41]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b42  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [42]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b43  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [43]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b44  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [44]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b45  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [45]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b46  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [46]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b47  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [47]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b48  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [48]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b49  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [49]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b5  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [5]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b50  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [50]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b51  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [51]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b52  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [52]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b53  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [53]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b54  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [54]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b55  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [55]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b56  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [56]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b57  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [57]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b58  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [58]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b59  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [59]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b6  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [6]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b60  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [60]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b61  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [61]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b62  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [62]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b63  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [63]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b7  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n158 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b8  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [8]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg5_b9  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/pte_temp [9]),
    .en(\biu/cache_ctrl_logic/n149 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/l1d_pte [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(407)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b0  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b1  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b10  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b100  (
    .clk(clk),
    .d(\biu/paddress [100]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [100]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b101  (
    .clk(clk),
    .d(\biu/paddress [101]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [101]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b102  (
    .clk(clk),
    .d(\biu/paddress [102]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [102]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b103  (
    .clk(clk),
    .d(\biu/paddress [103]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [103]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b104  (
    .clk(clk),
    .d(\biu/paddress [104]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [104]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b105  (
    .clk(clk),
    .d(\biu/paddress [105]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [105]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b106  (
    .clk(clk),
    .d(\biu/paddress [106]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [106]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b107  (
    .clk(clk),
    .d(\biu/paddress [107]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [107]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b108  (
    .clk(clk),
    .d(\biu/paddress [108]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [108]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b109  (
    .clk(clk),
    .d(\biu/paddress [109]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [109]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b11  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b110  (
    .clk(clk),
    .d(\biu/paddress [110]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [110]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b111  (
    .clk(clk),
    .d(\biu/paddress [111]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [111]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b112  (
    .clk(clk),
    .d(\biu/paddress [112]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [112]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b113  (
    .clk(clk),
    .d(\biu/paddress [113]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [113]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b114  (
    .clk(clk),
    .d(\biu/paddress [114]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [114]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b115  (
    .clk(clk),
    .d(\biu/paddress [115]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [115]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b116  (
    .clk(clk),
    .d(\biu/paddress [116]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [116]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b117  (
    .clk(clk),
    .d(\biu/paddress [117]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [117]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b118  (
    .clk(clk),
    .d(\biu/paddress [118]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [118]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b119  (
    .clk(clk),
    .d(\biu/paddress [119]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [119]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b12  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b120  (
    .clk(clk),
    .d(\biu/paddress [120]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [120]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b121  (
    .clk(clk),
    .d(\biu/paddress [121]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [121]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b122  (
    .clk(clk),
    .d(\biu/paddress [122]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [122]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b123  (
    .clk(clk),
    .d(\biu/paddress [123]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [123]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b124  (
    .clk(clk),
    .d(\biu/paddress [124]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [124]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b125  (
    .clk(clk),
    .d(\biu/paddress [125]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [125]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b126  (
    .clk(clk),
    .d(\biu/paddress [126]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [126]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b127  (
    .clk(clk),
    .d(\biu/paddress [127]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [127]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b13  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b14  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b15  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b16  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b17  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b18  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b19  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b2  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b20  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b21  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b22  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b23  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b24  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b25  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b26  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b27  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b28  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b29  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b3  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b30  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b31  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b32  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b33  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b34  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b35  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b36  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b37  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b38  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b39  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b4  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b40  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b41  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b42  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b43  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b44  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b45  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b46  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b47  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b48  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b49  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b5  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b50  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b51  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b52  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b53  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b54  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b55  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b56  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b57  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b58  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b59  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b6  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b60  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b61  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b62  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b63  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b64  (
    .clk(clk),
    .d(\biu/paddress [64]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [64]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b65  (
    .clk(clk),
    .d(\biu/paddress [65]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [65]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b66  (
    .clk(clk),
    .d(\biu/paddress [66]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [66]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b67  (
    .clk(clk),
    .d(\biu/paddress [67]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [67]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b68  (
    .clk(clk),
    .d(\biu/paddress [68]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [68]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b69  (
    .clk(clk),
    .d(\biu/paddress [69]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [69]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b7  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b70  (
    .clk(clk),
    .d(\biu/paddress [70]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [70]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b71  (
    .clk(clk),
    .d(\biu/paddress [71]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [71]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b72  (
    .clk(clk),
    .d(\biu/paddress [72]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [72]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b73  (
    .clk(clk),
    .d(\biu/paddress [73]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [73]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b74  (
    .clk(clk),
    .d(\biu/paddress [74]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [74]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b75  (
    .clk(clk),
    .d(\biu/paddress [75]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [75]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b76  (
    .clk(clk),
    .d(\biu/paddress [76]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [76]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b77  (
    .clk(clk),
    .d(\biu/paddress [77]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [77]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b78  (
    .clk(clk),
    .d(\biu/paddress [78]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [78]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b79  (
    .clk(clk),
    .d(\biu/paddress [79]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [79]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b8  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b80  (
    .clk(clk),
    .d(\biu/paddress [80]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [80]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b81  (
    .clk(clk),
    .d(\biu/paddress [81]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [81]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b82  (
    .clk(clk),
    .d(\biu/paddress [82]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [82]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b83  (
    .clk(clk),
    .d(\biu/paddress [83]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [83]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b84  (
    .clk(clk),
    .d(\biu/paddress [84]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [84]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b85  (
    .clk(clk),
    .d(\biu/paddress [85]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [85]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b86  (
    .clk(clk),
    .d(\biu/paddress [86]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [86]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b87  (
    .clk(clk),
    .d(\biu/paddress [87]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [87]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b88  (
    .clk(clk),
    .d(\biu/paddress [88]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [88]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b89  (
    .clk(clk),
    .d(\biu/paddress [89]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [89]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b9  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n166 [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b90  (
    .clk(clk),
    .d(\biu/paddress [90]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [90]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b91  (
    .clk(clk),
    .d(\biu/paddress [91]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [91]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b92  (
    .clk(clk),
    .d(\biu/paddress [92]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [92]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b93  (
    .clk(clk),
    .d(\biu/paddress [93]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [93]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b94  (
    .clk(clk),
    .d(\biu/paddress [94]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [94]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b95  (
    .clk(clk),
    .d(\biu/paddress [95]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [95]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b96  (
    .clk(clk),
    .d(\biu/paddress [96]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [96]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b97  (
    .clk(clk),
    .d(\biu/paddress [97]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [97]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b98  (
    .clk(clk),
    .d(\biu/paddress [98]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [98]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg6_b99  (
    .clk(clk),
    .d(\biu/paddress [99]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pa_temp [99]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b0  (
    .clk(clk),
    .d(uncache_data[0]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b1  (
    .clk(clk),
    .d(uncache_data[1]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b10  (
    .clk(clk),
    .d(uncache_data[10]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [10]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b11  (
    .clk(clk),
    .d(uncache_data[11]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [11]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b12  (
    .clk(clk),
    .d(uncache_data[12]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [12]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b13  (
    .clk(clk),
    .d(uncache_data[13]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [13]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b14  (
    .clk(clk),
    .d(uncache_data[14]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [14]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b15  (
    .clk(clk),
    .d(uncache_data[15]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [15]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b16  (
    .clk(clk),
    .d(uncache_data[16]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [16]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b17  (
    .clk(clk),
    .d(uncache_data[17]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [17]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b18  (
    .clk(clk),
    .d(uncache_data[18]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [18]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b19  (
    .clk(clk),
    .d(uncache_data[19]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [19]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b2  (
    .clk(clk),
    .d(uncache_data[2]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b20  (
    .clk(clk),
    .d(uncache_data[20]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [20]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b21  (
    .clk(clk),
    .d(uncache_data[21]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [21]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b22  (
    .clk(clk),
    .d(uncache_data[22]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [22]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b23  (
    .clk(clk),
    .d(uncache_data[23]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [23]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b24  (
    .clk(clk),
    .d(uncache_data[24]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [24]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b25  (
    .clk(clk),
    .d(uncache_data[25]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [25]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b26  (
    .clk(clk),
    .d(uncache_data[26]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [26]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b27  (
    .clk(clk),
    .d(uncache_data[27]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [27]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b28  (
    .clk(clk),
    .d(uncache_data[28]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [28]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b29  (
    .clk(clk),
    .d(uncache_data[29]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [29]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b3  (
    .clk(clk),
    .d(uncache_data[3]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b30  (
    .clk(clk),
    .d(uncache_data[30]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [30]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b31  (
    .clk(clk),
    .d(uncache_data[31]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [31]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b32  (
    .clk(clk),
    .d(uncache_data[32]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [32]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b33  (
    .clk(clk),
    .d(uncache_data[33]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [33]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b34  (
    .clk(clk),
    .d(uncache_data[34]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [34]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b35  (
    .clk(clk),
    .d(uncache_data[35]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [35]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b36  (
    .clk(clk),
    .d(uncache_data[36]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [36]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b37  (
    .clk(clk),
    .d(uncache_data[37]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [37]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b38  (
    .clk(clk),
    .d(uncache_data[38]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [38]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b39  (
    .clk(clk),
    .d(uncache_data[39]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [39]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b4  (
    .clk(clk),
    .d(uncache_data[4]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b40  (
    .clk(clk),
    .d(uncache_data[40]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [40]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b41  (
    .clk(clk),
    .d(uncache_data[41]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [41]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b42  (
    .clk(clk),
    .d(uncache_data[42]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [42]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b43  (
    .clk(clk),
    .d(uncache_data[43]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [43]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b44  (
    .clk(clk),
    .d(uncache_data[44]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [44]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b45  (
    .clk(clk),
    .d(uncache_data[45]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [45]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b46  (
    .clk(clk),
    .d(uncache_data[46]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [46]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b47  (
    .clk(clk),
    .d(uncache_data[47]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [47]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b48  (
    .clk(clk),
    .d(uncache_data[48]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [48]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b49  (
    .clk(clk),
    .d(uncache_data[49]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [49]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b5  (
    .clk(clk),
    .d(uncache_data[5]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [5]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b50  (
    .clk(clk),
    .d(uncache_data[50]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [50]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b51  (
    .clk(clk),
    .d(uncache_data[51]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [51]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b52  (
    .clk(clk),
    .d(uncache_data[52]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [52]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b53  (
    .clk(clk),
    .d(uncache_data[53]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [53]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b54  (
    .clk(clk),
    .d(uncache_data[54]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [54]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b55  (
    .clk(clk),
    .d(uncache_data[55]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [55]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b56  (
    .clk(clk),
    .d(uncache_data[56]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [56]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b57  (
    .clk(clk),
    .d(uncache_data[57]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [57]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b58  (
    .clk(clk),
    .d(uncache_data[58]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [58]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b59  (
    .clk(clk),
    .d(uncache_data[59]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [59]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b6  (
    .clk(clk),
    .d(uncache_data[6]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [6]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b60  (
    .clk(clk),
    .d(uncache_data[60]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [60]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b61  (
    .clk(clk),
    .d(uncache_data[61]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [61]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b62  (
    .clk(clk),
    .d(uncache_data[62]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [62]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b63  (
    .clk(clk),
    .d(uncache_data[63]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [63]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b7  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n165 [7]),
    .en(~\biu/cache_ctrl_logic/n161 ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [7]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b8  (
    .clk(clk),
    .d(uncache_data[8]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [8]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg7_b9  (
    .clk(clk),
    .d(uncache_data[9]),
    .en(\biu/cache_ctrl_logic/mux59_b100_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/pte_temp [9]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(429)
  reg_sr_ss_w1 \biu/cache_ctrl_logic/reg8_b0  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n132 [0]),
    .en(1'b1),
    .reset(rst),
    .set(\biu/cache_ctrl_logic/n56 ),
    .q(\biu/cache_ctrl_logic/statu [0]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  reg_sr_ss_w1 \biu/cache_ctrl_logic/reg8_b1  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n131 [1]),
    .en(1'b1),
    .reset(rst),
    .set(~\biu/cache_ctrl_logic/mux43_b1_sel_is_0_o ),
    .q(\biu/cache_ctrl_logic/statu [1]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg8_b2  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n132 [2]),
    .en(1'b1),
    .reset(~\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/statu [2]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  reg_sr_as_w1 \biu/cache_ctrl_logic/reg8_b3  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n132 [3]),
    .en(1'b1),
    .reset(~\biu/cache_ctrl_logic/mux44_b2_sel_is_0_o ),
    .set(1'b0),
    .q(\biu/cache_ctrl_logic/statu [3]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  reg_sr_ss_w1 \biu/cache_ctrl_logic/reg8_b4  (
    .clk(clk),
    .d(\biu/cache_ctrl_logic/n127 [4]),
    .en(1'b1),
    .reset(~\biu/cache_ctrl_logic/mux44_b4_sel_is_2_o ),
    .set(\biu/cache_ctrl_logic/n65 ),
    .q(\biu/cache_ctrl_logic/statu [4]));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(312)
  or \biu/cache_ctrl_logic/u10  (\biu/cache_ctrl_logic/n232 [17], \biu/cache_ctrl_logic/n230 [17], \biu/cache_ctrl_logic/n231 [17]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u100  (\biu/cache_ctrl_logic/n78 , \biu/trans_rdy , write);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  and \biu/cache_ctrl_logic/u101  (\biu/cache_ctrl_logic/n79 , \biu/trans_rdy , read);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  or \biu/cache_ctrl_logic/u102  (\biu/write_data [58], \biu/cache_ctrl_logic/n232 [58], \biu/cache_ctrl_logic/n233 [58]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u103  (\biu/cache_ctrl_logic/n85 , \biu/bus_error , write);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(264)
  and \biu/cache_ctrl_logic/u104  (\biu/cache_ctrl_logic/n86 , \biu/bus_error , read);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(264)
  or \biu/cache_ctrl_logic/u105  (\biu/write_data [57], \biu/cache_ctrl_logic/n232 [57], \biu/cache_ctrl_logic/n233 [57]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u106  (\biu/cache_ctrl_logic/n89 , \biu/trans_rdy , \biu/cache_ctrl_logic/pte_temp [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(269)
  or \biu/cache_ctrl_logic/u107  (\biu/write_data [56], \biu/cache_ctrl_logic/n232 [56], \biu/cache_ctrl_logic/n233 [56]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u108  (\biu/write_data [55], \biu/cache_ctrl_logic/n232 [55], \biu/cache_ctrl_logic/n233 [55]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u109  (\biu/write_data [54], \biu/cache_ctrl_logic/n232 [54], \biu/cache_ctrl_logic/n233 [54]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u11  (\biu/cache_ctrl_logic/n232 [16], \biu/cache_ctrl_logic/n230 [16], \biu/cache_ctrl_logic/n231 [16]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u110  (\biu/cache_ctrl_logic/n94 , \biu/trans_rdy , \biu/cache_ctrl_logic/n0 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(277)
  or \biu/cache_ctrl_logic/u111  (\biu/write_data [53], \biu/cache_ctrl_logic/n232 [53], \biu/cache_ctrl_logic/n233 [53]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u112  (\biu/write_data [52], \biu/cache_ctrl_logic/n232 [52], \biu/cache_ctrl_logic/n233 [52]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u113  (\biu/cache_ctrl_logic/n98 , \biu/trans_rdy , \biu/cache_ctrl_logic/n1 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(280)
  or \biu/cache_ctrl_logic/u114  (\biu/write_data [51], \biu/cache_ctrl_logic/n232 [51], \biu/cache_ctrl_logic/n233 [51]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u115  (\biu/write_data [50], \biu/cache_ctrl_logic/n232 [50], \biu/cache_ctrl_logic/n233 [50]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u116  (\biu/write_data [49], \biu/cache_ctrl_logic/n232 [49], \biu/cache_ctrl_logic/n233 [49]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u117  (\biu/cache_ctrl_logic/n232 [19], \biu/cache_ctrl_logic/n230 [19], \biu/cache_ctrl_logic/n231 [19]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u118  (\biu/write_data [48], \biu/cache_ctrl_logic/n232 [48], \biu/cache_ctrl_logic/n233 [48]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u119  (\biu/cache_ctrl_logic/n135 , \biu/cache_ctrl_logic/l1i_wr_sel , \biu/trans_rdy );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(320)
  or \biu/cache_ctrl_logic/u12  (\biu/cache_ctrl_logic/n2 , read, write);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(187)
  or \biu/cache_ctrl_logic/u120  (\biu/write_data [47], \biu/cache_ctrl_logic/n232 [47], \biu/cache_ctrl_logic/n233 [47]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u121  (\biu/cache_ctrl_logic/n139 , \biu/cache_ctrl_logic/l1d_wr_sel , \biu/cache_ctrl_logic/n138 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(330)
  and \biu/cache_ctrl_logic/u122  (\biu/cache_ctrl_logic/n140 , \biu/cache_ctrl_logic/n139 , \biu/trans_rdy );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(330)
  or \biu/cache_ctrl_logic/u123  (\biu/write_data [46], \biu/cache_ctrl_logic/n232 [46], \biu/cache_ctrl_logic/n233 [46]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u124  (\biu/write_data [45], \biu/cache_ctrl_logic/n232 [45], \biu/cache_ctrl_logic/n233 [45]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u125  (\biu/write_data [44], \biu/cache_ctrl_logic/n232 [44], \biu/cache_ctrl_logic/n233 [44]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u128_sel_is_0  (\biu/cache_ctrl_logic/u128_sel_is_0_o , rst_neg, \biu/cache_ctrl_logic/n67_neg );
  or \biu/cache_ctrl_logic/u129  (\biu/write_data [43], \biu/cache_ctrl_logic/n232 [43], \biu/cache_ctrl_logic/n233 [43]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u13  (\biu/cache_ctrl_logic/n4 , \biu/cache_ctrl_logic/n2 , \biu/cache_ctrl_logic/n3 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(187)
  or \biu/cache_ctrl_logic/u130  (\biu/write_data [42], \biu/cache_ctrl_logic/n232 [42], \biu/cache_ctrl_logic/n233 [42]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u131  (\biu/write_data [41], \biu/cache_ctrl_logic/n232 [41], \biu/cache_ctrl_logic/n233 [41]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  AL_MUX \biu/cache_ctrl_logic/u132  (
    .i0(\biu/cache_ctrl_logic/l1i_pte [7]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n102 ),
    .o(\biu/cache_ctrl_logic/n146 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(361)
  or \biu/cache_ctrl_logic/u133  (\biu/write_data [40], \biu/cache_ctrl_logic/n232 [40], \biu/cache_ctrl_logic/n233 [40]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u134  (\biu/cache_ctrl_logic/n149 , \biu/cache_ctrl_logic/l1d_wr_sel , \biu/trans_rdy );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(369)
  or \biu/cache_ctrl_logic/u135  (\biu/write_data [39], \biu/cache_ctrl_logic/n232 [39], \biu/cache_ctrl_logic/n233 [39]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u136  (\biu/write_data [38], \biu/cache_ctrl_logic/n232 [38], \biu/cache_ctrl_logic/n233 [38]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u137  (\biu/write_data [37], \biu/cache_ctrl_logic/n232 [37], \biu/cache_ctrl_logic/n233 [37]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u138  (\biu/write_data [36], \biu/cache_ctrl_logic/n232 [36], \biu/cache_ctrl_logic/n233 [36]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u139  (\biu/write_data [35], \biu/cache_ctrl_logic/n232 [35], \biu/cache_ctrl_logic/n233 [35]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u14  (\biu/cache_ctrl_logic/ex_l1i_hit , \biu/cache_ctrl_logic/n4 , \biu/cache_ctrl_logic/l1i_value );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(187)
  or \biu/cache_ctrl_logic/u143  (\biu/write_data [34], \biu/cache_ctrl_logic/n232 [34], \biu/cache_ctrl_logic/n233 [34]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u144  (\biu/write_data [33], \biu/cache_ctrl_logic/n232 [33], \biu/cache_ctrl_logic/n233 [33]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u145  (\biu/write_data [32], \biu/cache_ctrl_logic/n232 [32], \biu/cache_ctrl_logic/n233 [32]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  AL_MUX \biu/cache_ctrl_logic/u146  (
    .i0(\biu/cache_ctrl_logic/l1d_pte [7]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n104 ),
    .o(\biu/cache_ctrl_logic/n157 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(406)
  or \biu/cache_ctrl_logic/u147  (\biu/write_data [31], \biu/cache_ctrl_logic/n232 [31], \biu/cache_ctrl_logic/n233 [31]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u148  (\biu/cache_ctrl_logic/n160 , \biu/cache_ctrl_logic/n55 , unpage);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(418)
  or \biu/cache_ctrl_logic/u149  (\biu/write_data [30], \biu/cache_ctrl_logic/n232 [30], \biu/cache_ctrl_logic/n233 [30]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u15  (\biu/cache_ctrl_logic/n232 [15], \biu/cache_ctrl_logic/n230 [15], \biu/cache_ctrl_logic/n231 [15]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u150  (\biu/cache_ctrl_logic/n161 , \biu/cache_ctrl_logic/n160 , \biu/cache_ctrl_logic/n2 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(418)
  or \biu/cache_ctrl_logic/u151  (\biu/write_data [29], \biu/cache_ctrl_logic/n232 [29], \biu/cache_ctrl_logic/n233 [29]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u152  (\biu/write_data [28], \biu/cache_ctrl_logic/n232 [28], \biu/cache_ctrl_logic/n233 [28]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u153  (\biu/pa_cov , \biu/opc [1], \biu/cache_ctrl_logic/n75 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(421)
  and \biu/cache_ctrl_logic/u154  (\biu/cache_ctrl_logic/n162 , \biu/pa_cov , \biu/trans_rdy );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(421)
  or \biu/cache_ctrl_logic/u155  (\biu/write_data [27], \biu/cache_ctrl_logic/n232 [27], \biu/cache_ctrl_logic/n233 [27]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  AL_MUX \biu/cache_ctrl_logic/u156  (
    .i0(\biu/cache_ctrl_logic/pte_temp [7]),
    .i1(1'b1),
    .sel(\biu/cache_ctrl_logic/n101 ),
    .o(\biu/cache_ctrl_logic/n163 ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(428)
  or \biu/cache_ctrl_logic/u157  (\biu/write_data [26], \biu/cache_ctrl_logic/n232 [26], \biu/cache_ctrl_logic/n233 [26]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u158  (\biu/write_data [25], \biu/cache_ctrl_logic/n232 [25], \biu/cache_ctrl_logic/n233 [25]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u159  (\biu/write_data [24], \biu/cache_ctrl_logic/n232 [24], \biu/cache_ctrl_logic/n233 [24]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u16  (\biu/cache_ctrl_logic/n6 , \biu/cache_ctrl_logic/n2 , \biu/cache_ctrl_logic/n5 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(188)
  or \biu/cache_ctrl_logic/u160  (\biu/write_data [23], \biu/cache_ctrl_logic/n232 [23], \biu/cache_ctrl_logic/n233 [23]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u161  (\biu/cache_addr_sel , \biu/cache_ctrl_logic/l1i_wr_sel , \biu/cache_ctrl_logic/l1d_wr_sel );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(436)
  or \biu/cache_ctrl_logic/u162  (\biu/write_data [22], \biu/cache_ctrl_logic/n232 [22], \biu/cache_ctrl_logic/n233 [22]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u163  (\biu/write_data [21], \biu/cache_ctrl_logic/n232 [21], \biu/cache_ctrl_logic/n233 [21]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u164  (\biu/cache_ctrl_logic/ex_bsel [1], \biu/cache_ctrl_logic/n182 [7], \biu/cache_ctrl_logic/n182 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(473)
  or \biu/cache_ctrl_logic/u165  (\biu/write_data [20], \biu/cache_ctrl_logic/n232 [20], \biu/cache_ctrl_logic/n233 [20]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u166  (\biu/cache_ctrl_logic/n170 , \biu/cache_ctrl_logic/n55 , \biu/cache_ctrl_logic/ex_l1i_hit );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(440)
  or \biu/cache_ctrl_logic/u167  (\biu/write_data [19], \biu/cache_ctrl_logic/n232 [19], \biu/cache_ctrl_logic/n233 [19]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u168  (\biu/cache_ctrl_logic/n171 , \biu/cache_ctrl_logic/n55 , \biu/cache_ctrl_logic/ex_l1d_hit );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(442)
  or \biu/cache_ctrl_logic/u169  (\biu/cache_ctrl_logic/n175 , \biu/cache_ctrl_logic/n173 , \biu/cache_ctrl_logic/n174 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(445)
  and \biu/cache_ctrl_logic/u17  (\biu/cache_ctrl_logic/ex_l1d_hit , \biu/cache_ctrl_logic/n6 , \biu/cache_ctrl_logic/l1d_value );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(188)
  or \biu/cache_ctrl_logic/u170  (\biu/cache_ctrl_logic/n177 , \biu/cache_ctrl_logic/n175 , \biu/cache_ctrl_logic/n176 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(445)
  or \biu/cache_ctrl_logic/u171  (\biu/cache_ctrl_logic/n179 , \biu/cache_ctrl_logic/n177 , \biu/cache_ctrl_logic/n178 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(445)
  and \biu/cache_ctrl_logic/u172  (\biu/cache_ctrl_logic/ex_bsel [0], \biu/cache_ctrl_logic/n172 , \biu/cache_ctrl_logic/n179 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(445)
  or \biu/cache_ctrl_logic/u173  (\biu/write_data [18], \biu/cache_ctrl_logic/n232 [18], \biu/cache_ctrl_logic/n233 [18]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u174  (\biu/write_data [17], \biu/cache_ctrl_logic/n232 [17], \biu/cache_ctrl_logic/n233 [17]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u175  (\biu/write_data [16], \biu/cache_ctrl_logic/n232 [16], \biu/cache_ctrl_logic/n233 [16]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u176  (\biu/write_data [15], \biu/cache_ctrl_logic/n232 [15], \biu/cache_ctrl_logic/n233 [15]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u177  (\biu/write_data [14], \biu/cache_ctrl_logic/n232 [14], \biu/cache_ctrl_logic/n233 [14]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u18  (\biu/cache_ctrl_logic/n8 , rd_ins, \biu/cache_ctrl_logic/n7 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(189)
  or \biu/cache_ctrl_logic/u180  (\biu/write_data [13], \biu/cache_ctrl_logic/n232 [13], \biu/cache_ctrl_logic/n233 [13]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u181  (\biu/write_data [12], \biu/cache_ctrl_logic/n232 [12], \biu/cache_ctrl_logic/n233 [12]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u182  (\biu/write_data [11], \biu/cache_ctrl_logic/n232 [11], \biu/cache_ctrl_logic/n233 [11]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u183  (\biu/write_data [10], \biu/cache_ctrl_logic/n232 [10], \biu/cache_ctrl_logic/n233 [10]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u184  (\biu/write_data [9], \biu/cache_ctrl_logic/n232 [9], \biu/cache_ctrl_logic/n233 [9]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u185  (\biu/cache_ctrl_logic/n232 [24], \biu/cache_ctrl_logic/n230 [24], \biu/cache_ctrl_logic/n231 [24]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u186  (\biu/cache_ctrl_logic/n232 [62], \biu/cache_ctrl_logic/n230 [62], \biu/cache_ctrl_logic/n231 [62]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u187  (\biu/write_data [8], \biu/cache_ctrl_logic/n232 [8], \biu/cache_ctrl_logic/n233 [8]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u188  (\biu/write_data [7], \biu/cache_ctrl_logic/n232 [7], \biu/cache_ctrl_logic/n233 [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u189  (\biu/write_data [6], \biu/cache_ctrl_logic/n232 [6], \biu/cache_ctrl_logic/n233 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  and \biu/cache_ctrl_logic/u19  (\biu/cache_ctrl_logic/if_l1i_hit , \biu/cache_ctrl_logic/n8 , \biu/cache_ctrl_logic/l1i_value );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(189)
  or \biu/cache_ctrl_logic/u190  (\biu/cache_ctrl_logic/n184 [3], \biu/cache_ctrl_logic/n174 , \biu/cache_ctrl_logic/n176 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(448)
  and \biu/cache_ctrl_logic/u191  (\biu/cache_ctrl_logic/n182 [0], \biu/cache_ctrl_logic/n183 , \biu/cache_ctrl_logic/n177 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(446)
  or \biu/cache_ctrl_logic/u192  (\biu/write_data [5], \biu/cache_ctrl_logic/n232 [5], \biu/cache_ctrl_logic/n233 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u193  (\biu/write_data [4], \biu/cache_ctrl_logic/n232 [4], \biu/cache_ctrl_logic/n233 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u194  (\biu/write_data [3], \biu/cache_ctrl_logic/n232 [3], \biu/cache_ctrl_logic/n233 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u195  (\biu/cache_ctrl_logic/n232 [28], \biu/cache_ctrl_logic/n230 [28], \biu/cache_ctrl_logic/n231 [28]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u196  (\biu/cache_ctrl_logic/n232 [34], \biu/cache_ctrl_logic/n230 [34], \biu/cache_ctrl_logic/n231 [34]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u197  (\biu/cache_ctrl_logic/n232 [56], \biu/cache_ctrl_logic/n230 [56], \biu/cache_ctrl_logic/n231 [56]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u198  (\biu/write_data [2], \biu/cache_ctrl_logic/n232 [2], \biu/cache_ctrl_logic/n233 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u199  (\biu/write_data [1], \biu/cache_ctrl_logic/n232 [1], \biu/cache_ctrl_logic/n233 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  not \biu/cache_ctrl_logic/u2  (\biu/cache_ctrl_logic/n60 [0], \biu/cache_ctrl_logic/n59 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(223)
  not \biu/cache_ctrl_logic/u20  (\biu/cache_ctrl_logic/n9 , \biu/cache_ctrl_logic/if_l1i_hit );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(192)
  or \biu/cache_ctrl_logic/u203  (\biu/cache_ctrl_logic/n232 [23], \biu/cache_ctrl_logic/n230 [23], \biu/cache_ctrl_logic/n231 [23]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u204  (\biu/cache_ctrl_logic/n232 [61], \biu/cache_ctrl_logic/n230 [61], \biu/cache_ctrl_logic/n231 [61]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u208  (\biu/cache_ctrl_logic/n188 , \biu/cache_ctrl_logic/n176 , \biu/cache_ctrl_logic/n178 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(451)
  or \biu/cache_ctrl_logic/u209  (\biu/cache_ctrl_logic/n232 [42], \biu/cache_ctrl_logic/n230 [42], \biu/cache_ctrl_logic/n231 [42]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u21  (\biu/cache_ctrl_logic/l1i_miss , rd_ins, \biu/cache_ctrl_logic/n9 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(192)
  or \biu/cache_ctrl_logic/u212  (\biu/cache_ctrl_logic/n232 [47], \biu/cache_ctrl_logic/n230 [47], \biu/cache_ctrl_logic/n231 [47]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u213  (\biu/cache_ctrl_logic/n232 [51], \biu/cache_ctrl_logic/n230 [51], \biu/cache_ctrl_logic/n231 [51]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u217  (\biu/cache_ctrl_logic/n232 [27], \biu/cache_ctrl_logic/n230 [27], \biu/cache_ctrl_logic/n231 [27]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u218  (\biu/cache_ctrl_logic/n232 [33], \biu/cache_ctrl_logic/n230 [33], \biu/cache_ctrl_logic/n231 [33]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u219  (\biu/cache_ctrl_logic/n232 [55], \biu/cache_ctrl_logic/n230 [55], \biu/cache_ctrl_logic/n231 [55]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u22  (\biu/cache_ctrl_logic/n232 [14], \biu/cache_ctrl_logic/n230 [14], \biu/cache_ctrl_logic/n231 [14]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u225  (\biu/cache_ctrl_logic/n232 [22], \biu/cache_ctrl_logic/n230 [22], \biu/cache_ctrl_logic/n231 [22]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u226  (\biu/cache_ctrl_logic/n232 [60], \biu/cache_ctrl_logic/n230 [60], \biu/cache_ctrl_logic/n231 [60]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u229  (\biu/cache_ctrl_logic/n232 [36], \biu/cache_ctrl_logic/n230 [36], \biu/cache_ctrl_logic/n231 [36]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  not \biu/cache_ctrl_logic/u23  (\biu/cache_ctrl_logic/n10 , \biu/cache_ctrl_logic/ex_l1d_hit );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(193)
  or \biu/cache_ctrl_logic/u232  (\biu/cache_ctrl_logic/n232 [39], \biu/cache_ctrl_logic/n230 [39], \biu/cache_ctrl_logic/n231 [39]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u233  (\biu/cache_ctrl_logic/n232 [41], \biu/cache_ctrl_logic/n230 [41], \biu/cache_ctrl_logic/n231 [41]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u236  (\biu/cache_ctrl_logic/n232 [46], \biu/cache_ctrl_logic/n230 [46], \biu/cache_ctrl_logic/n231 [46]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u237  (\biu/cache_ctrl_logic/n232 [50], \biu/cache_ctrl_logic/n230 [50], \biu/cache_ctrl_logic/n231 [50]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u24  (\biu/cache_ctrl_logic/n11 , \biu/cache_ctrl_logic/n2 , \biu/cache_ctrl_logic/n10 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(193)
  or \biu/cache_ctrl_logic/u241  (\biu/cache_ctrl_logic/n232 [26], \biu/cache_ctrl_logic/n230 [26], \biu/cache_ctrl_logic/n231 [26]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u242  (\biu/cache_ctrl_logic/n232 [32], \biu/cache_ctrl_logic/n230 [32], \biu/cache_ctrl_logic/n231 [32]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u243  (\biu/cache_ctrl_logic/n232 [54], \biu/cache_ctrl_logic/n230 [54], \biu/cache_ctrl_logic/n231 [54]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u249  (\biu/cache_ctrl_logic/n232 [21], \biu/cache_ctrl_logic/n230 [21], \biu/cache_ctrl_logic/n231 [21]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u25  (\biu/cache_ctrl_logic/n232 [13], \biu/cache_ctrl_logic/n230 [13], \biu/cache_ctrl_logic/n231 [13]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u250  (\biu/cache_ctrl_logic/n232 [59], \biu/cache_ctrl_logic/n230 [59], \biu/cache_ctrl_logic/n231 [59]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u253  (\biu/cache_ctrl_logic/n232 [35], \biu/cache_ctrl_logic/n230 [35], \biu/cache_ctrl_logic/n231 [35]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u256  (\biu/cache_ctrl_logic/n232 [38], \biu/cache_ctrl_logic/n230 [38], \biu/cache_ctrl_logic/n231 [38]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u257  (\biu/cache_ctrl_logic/n232 [40], \biu/cache_ctrl_logic/n230 [40], \biu/cache_ctrl_logic/n231 [40]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u26  (\biu/cache_ctrl_logic/l1d_miss , \biu/cache_ctrl_logic/n11 , \biu/cache_ctrl_logic/n10 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(193)
  or \biu/cache_ctrl_logic/u260  (\biu/cache_ctrl_logic/n232 [45], \biu/cache_ctrl_logic/n230 [45], \biu/cache_ctrl_logic/n231 [45]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u261  (\biu/cache_ctrl_logic/n232 [49], \biu/cache_ctrl_logic/n230 [49], \biu/cache_ctrl_logic/n231 [49]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u265  (\biu/cache_ctrl_logic/n232 [25], \biu/cache_ctrl_logic/n230 [25], \biu/cache_ctrl_logic/n231 [25]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u266  (\biu/cache_ctrl_logic/n232 [31], \biu/cache_ctrl_logic/n230 [31], \biu/cache_ctrl_logic/n231 [31]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u267  (\biu/cache_ctrl_logic/n232 [53], \biu/cache_ctrl_logic/n230 [53], \biu/cache_ctrl_logic/n231 [53]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u27  (\biu/cache_ctrl_logic/n13 , \biu/cache_ctrl_logic/n12 , \biu/cache_ctrl_logic/l1i_pte [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(201)
  or \biu/cache_ctrl_logic/u271  (\biu/cache_ctrl_logic/n232 [20], \biu/cache_ctrl_logic/n230 [20], \biu/cache_ctrl_logic/n231 [20]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u272  (\biu/cache_ctrl_logic/n232 [58], \biu/cache_ctrl_logic/n230 [58], \biu/cache_ctrl_logic/n231 [58]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u275  (\biu/cache_ctrl_logic/n192 [0], \biu/cache_ctrl_logic/n183 , \biu/cache_ctrl_logic/n176 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(465)
  or \biu/cache_ctrl_logic/u278  (\biu/cache_ctrl_logic/n232 [37], \biu/cache_ctrl_logic/n230 [37], \biu/cache_ctrl_logic/n231 [37]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u279  (\biu/cache_ctrl_logic/n185 [0], \biu/cache_ctrl_logic/n183 , \biu/cache_ctrl_logic/n184 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(448)
  and \biu/cache_ctrl_logic/u28  (\biu/cache_ctrl_logic/n14 , write, \biu/cache_ctrl_logic/l1i_pte [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(201)
  or \biu/cache_ctrl_logic/u282  (\biu/cache_ctrl_logic/n232 [44], \biu/cache_ctrl_logic/n230 [44], \biu/cache_ctrl_logic/n231 [44]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u283  (\biu/cache_ctrl_logic/n232 [48], \biu/cache_ctrl_logic/n230 [48], \biu/cache_ctrl_logic/n231 [48]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u286  (\biu/cache_ctrl_logic/n232 [30], \biu/cache_ctrl_logic/n230 [30], \biu/cache_ctrl_logic/n231 [30]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u287  (\biu/cache_ctrl_logic/n232 [52], \biu/cache_ctrl_logic/n230 [52], \biu/cache_ctrl_logic/n231 [52]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u29  (\biu/cache_ctrl_logic/n15 , mxr, \biu/cache_ctrl_logic/l1i_pte [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(201)
  or \biu/cache_ctrl_logic/u292  (\biu/cache_ctrl_logic/n232 [57], \biu/cache_ctrl_logic/n230 [57], \biu/cache_ctrl_logic/n231 [57]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u298  (\biu/cache_ctrl_logic/n232 [43], \biu/cache_ctrl_logic/n230 [43], \biu/cache_ctrl_logic/n231 [43]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u3  (\biu/cache_ctrl_logic/n232 [18], \biu/cache_ctrl_logic/n230 [18], \biu/cache_ctrl_logic/n231 [18]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u30  (\biu/cache_ctrl_logic/n16 , \biu/cache_ctrl_logic/l1i_pte [1], \biu/cache_ctrl_logic/n15 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(201)
  or \biu/cache_ctrl_logic/u302  (\biu/cache_ctrl_logic/n232 [29], \biu/cache_ctrl_logic/n230 [29], \biu/cache_ctrl_logic/n231 [29]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u303  (\biu/cache_ctrl_logic/n193 [0], \biu/cache_ctrl_logic/n189 [6], \biu/cache_ctrl_logic/n192 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(466)
  or \biu/cache_ctrl_logic/u306  (\biu/cache_ctrl_logic/n190 [0], \biu/cache_ctrl_logic/n189 [5], \biu/cache_ctrl_logic/n192 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(471)
  AL_MUX \biu/cache_ctrl_logic/u308  (
    .i0(\biu/cache_ctrl_logic/l1i_write_through ),
    .i1(\biu/cache_ctrl_logic/l1i_write_burst ),
    .sel(\biu/cache_ctrl_logic/l1i_wr_sel ),
    .o(\biu/l1i_write ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(477)
  and \biu/cache_ctrl_logic/u31  (\biu/cache_ctrl_logic/n17 , read, \biu/cache_ctrl_logic/n16 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(201)
  AL_MUX \biu/cache_ctrl_logic/u310  (
    .i0(\biu/cache_ctrl_logic/l1d_write_through ),
    .i1(\biu/cache_ctrl_logic/l1d_write_burst ),
    .sel(\biu/cache_ctrl_logic/l1d_wr_sel ),
    .o(\biu/l1d_write ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(478)
  AL_MUX \biu/cache_ctrl_logic/u312  (
    .i0(1'b0),
    .i1(\biu/cache_write ),
    .sel(\biu/cache_ctrl_logic/l1d_wr_sel ),
    .o(\biu/cache_ctrl_logic/l1d_write_burst ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(479)
  AL_MUX \biu/cache_ctrl_logic/u314  (
    .i0(1'b0),
    .i1(\biu/cache_write ),
    .sel(\biu/cache_ctrl_logic/l1i_wr_sel ),
    .o(\biu/cache_ctrl_logic/l1i_write_burst ));  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(480)
  not \biu/cache_ctrl_logic/u315  (\biu/cache_ctrl_logic/n198 , \biu/cache_ctrl_logic/ex_l1d_chkok );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(482)
  and \biu/cache_ctrl_logic/u316  (\biu/ex_data_sel [0], \biu/cache_ctrl_logic/ex_l1i_chkok , \biu/cache_ctrl_logic/n198 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(482)
  or \biu/cache_ctrl_logic/u32  (\biu/cache_ctrl_logic/n18 , \biu/cache_ctrl_logic/n14 , \biu/cache_ctrl_logic/n17 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(201)
  or \biu/cache_ctrl_logic/u321  (\biu/rd , \biu/cache_addr_sel , \biu/ex_data_sel [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(486)
  or \biu/cache_ctrl_logic/u327  (\biu/cache_ctrl_logic/n199 , \biu/cache_addr_sel , \biu/cache_ctrl_logic/n101 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(488)
  or \biu/cache_ctrl_logic/u329  (\biu/cache_ctrl_logic/n200 , \biu/cache_ctrl_logic/n199 , \biu/cache_ctrl_logic/n102 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(488)
  and \biu/cache_ctrl_logic/u33  (\biu/cache_ctrl_logic/n19 , \biu/cache_ctrl_logic/n13 , \biu/cache_ctrl_logic/n18 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(201)
  or \biu/cache_ctrl_logic/u331  (\biu/cache_ctrl_logic/n201 , \biu/cache_ctrl_logic/n200 , \biu/cache_ctrl_logic/n104 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(488)
  or \biu/cache_ctrl_logic/u333  (\biu/cache_ctrl_logic/n202 , \biu/cache_ctrl_logic/n201 , \biu/cache_ctrl_logic/n93 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(488)
  or \biu/cache_ctrl_logic/u335  (\biu/paddr , \biu/cache_ctrl_logic/n202 , \biu/cache_ctrl_logic/n97 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(488)
  and \biu/cache_ctrl_logic/u34  (\biu/cache_ctrl_logic/n21 , sum, \biu/cache_ctrl_logic/l1i_pte [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(202)
  or \biu/cache_ctrl_logic/u344  (\biu/cache_ctrl_logic/n203 , \biu/cache_ctrl_logic/n102 , \biu/cache_ctrl_logic/n104 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(493)
  or \biu/cache_ctrl_logic/u346  (\biu/new_pte_update , \biu/cache_ctrl_logic/n203 , \biu/cache_ctrl_logic/n101 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(493)
  and \biu/cache_ctrl_logic/u349  (\biu/opc [0], \biu/cache_ctrl_logic/n75 , write);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(497)
  not \biu/cache_ctrl_logic/u35  (\biu/cache_ctrl_logic/n22 , \biu/cache_ctrl_logic/l1i_pte [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(202)
  or \biu/cache_ctrl_logic/u353  (\biu/cache_ctrl_logic/n204 , \biu/wr , \biu/ex_data_sel [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  or \biu/cache_ctrl_logic/u355  (\biu/cache_ctrl_logic/n205 , \biu/cache_ctrl_logic/n204 , \biu/cache_ctrl_logic/l1i_wr_sel );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  or \biu/cache_ctrl_logic/u357  (\biu/cache_ctrl_logic/n206 , \biu/cache_ctrl_logic/n205 , \biu/cache_ctrl_logic/l1d_wr_sel );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(503)
  or \biu/cache_ctrl_logic/u359  (\biu/cache_ctrl_logic/n186 [0], \biu/cache_ctrl_logic/n189 [5], \biu/cache_ctrl_logic/n185 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(472)
  or \biu/cache_ctrl_logic/u36  (\biu/cache_ctrl_logic/n23 , \biu/cache_ctrl_logic/n21 , \biu/cache_ctrl_logic/n22 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(202)
  or \biu/cache_ctrl_logic/u361  (\biu/cache_ctrl_logic/n211 [0], \biu/cache_ctrl_logic/n208 [0], \biu/cache_ctrl_logic/n210 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u363  (\biu/cache_ctrl_logic/n214 [0], \biu/cache_ctrl_logic/n211 [0], \biu/cache_ctrl_logic/n213 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u365  (\biu/cache_ctrl_logic/n216 [0], \biu/cache_ctrl_logic/n214 [0], \biu/cache_ctrl_logic/n215 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u367  (\biu/cache_ctrl_logic/n218 [0], \biu/cache_ctrl_logic/n216 [0], \biu/cache_ctrl_logic/n217 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u369  (\biu/cache_ctrl_logic/n220 [0], \biu/cache_ctrl_logic/n218 [0], \biu/cache_ctrl_logic/n219 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  and \biu/cache_ctrl_logic/u37  (\biu/cache_ctrl_logic/n24 , \biu/cache_ctrl_logic/n20 , \biu/cache_ctrl_logic/n23 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(202)
  or \biu/cache_ctrl_logic/u371  (\biu/cache_ctrl_logic/n222 [0], \biu/cache_ctrl_logic/n220 [0], \biu/cache_ctrl_logic/n221 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u376  (\biu/cache_ctrl_logic/n224 , \biu/cache_ctrl_logic/n204 , \biu/cache_ctrl_logic/n97 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  or \biu/cache_ctrl_logic/u378  (\biu/cache_ctrl_logic/n225 , \biu/cache_ctrl_logic/n224 , \biu/cache_ctrl_logic/n93 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(514)
  or \biu/cache_ctrl_logic/u38  (\biu/cache_ctrl_logic/n232 [12], \biu/cache_ctrl_logic/n230 [12], \biu/cache_ctrl_logic/n231 [12]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u381  (\biu/cache_ctrl_logic/n226 , \biu/wr , \biu/cache_ctrl_logic/n93 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  or \biu/cache_ctrl_logic/u383  (\biu/cache_ctrl_logic/n227 , \biu/cache_ctrl_logic/n226 , \biu/cache_ctrl_logic/n97 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(517)
  or \biu/cache_ctrl_logic/u385  (\biu/maddress [0], \biu/cache_ctrl_logic/n222 [0], \biu/cache_ctrl_logic/n223 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u387  (\biu/cache_ctrl_logic/n230 [0], \biu/cache_ctrl_logic/n228 [0], \biu/cache_ctrl_logic/n229 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u389  (\biu/cache_ctrl_logic/n232 [0], \biu/cache_ctrl_logic/n230 [0], \biu/cache_ctrl_logic/n231 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u39  (\biu/cache_ctrl_logic/n232 [11], \biu/cache_ctrl_logic/n230 [11], \biu/cache_ctrl_logic/n231 [11]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u390  (\biu/write_data [0], \biu/cache_ctrl_logic/n232 [0], \biu/cache_ctrl_logic/n233 [0]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  not \biu/cache_ctrl_logic/u394  (\biu/cache_ctrl_logic/n234 , \biu/cache_ctrl_logic/pte_l1i_upd );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(530)
  not \biu/cache_ctrl_logic/u395  (\biu/cache_ctrl_logic/n235 , \biu/cache_ctrl_logic/pte_l1d_upd );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(530)
  or \biu/cache_ctrl_logic/u396  (\biu/cache_ctrl_logic/n236 , \biu/cache_ctrl_logic/n234 , \biu/cache_ctrl_logic/n235 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(530)
  not \biu/cache_ctrl_logic/u397  (\biu/cache_ctrl_logic/n237 , \biu/cache_ctrl_logic/l1i_write_through );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(530)
  or \biu/cache_ctrl_logic/u398  (\biu/cache_ctrl_logic/n238 , \biu/cache_ctrl_logic/n236 , \biu/cache_ctrl_logic/n237 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(530)
  not \biu/cache_ctrl_logic/u399  (\biu/cache_ctrl_logic/n239 , \biu/cache_ctrl_logic/l1d_write_through );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(530)
  and \biu/cache_ctrl_logic/u4  (\biu/cache_ctrl_logic/l1i_write_through , \biu/cache_ctrl_logic/ex_l1i_chkok , write);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(180)
  or \biu/cache_ctrl_logic/u40  (\biu/cache_ctrl_logic/n232 [10], \biu/cache_ctrl_logic/n230 [10], \biu/cache_ctrl_logic/n231 [10]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u400  (\biu/cache_ctrl_logic/n240 , \biu/cache_ctrl_logic/n238 , \biu/cache_ctrl_logic/n239 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(530)
  and \biu/cache_ctrl_logic/u401  (\biu/cache_ctrl_logic/n241 , \biu/cache_ctrl_logic/n55 , \biu/cache_ctrl_logic/n240 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(530)
  and \biu/cache_ctrl_logic/u407  (\biu/cache_ctrl_logic/n242 , \biu/cache_ctrl_logic/n227 , \biu/trans_rdy );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(531)
  or \biu/cache_ctrl_logic/u408  (\biu/cache_ctrl_logic/n243 , \biu/cache_ctrl_logic/n241 , \biu/cache_ctrl_logic/n242 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(531)
  or \biu/cache_ctrl_logic/u41  (\biu/cache_ctrl_logic/n232 [9], \biu/cache_ctrl_logic/n230 [9], \biu/cache_ctrl_logic/n231 [9]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u412  (\biu/cache_ctrl_logic/n244 , \biu/cache_ctrl_logic/n203 , \biu/trans_rdy );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(532)
  or \biu/cache_ctrl_logic/u413  (\biu/cache_ctrl_logic/n245 , \biu/cache_ctrl_logic/n243 , \biu/cache_ctrl_logic/n244 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(532)
  or \biu/cache_ctrl_logic/u415  (cache_ready_ex, \biu/cache_ctrl_logic/n245 , \biu/cache_ctrl_logic/n67 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(533)
  and \biu/cache_ctrl_logic/u417  (uncache_data_rdy, \biu/ex_data_sel [1], \biu/trans_rdy );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(535)
  or \biu/cache_ctrl_logic/u42  (\biu/cache_ctrl_logic/n232 [8], \biu/cache_ctrl_logic/n230 [8], \biu/cache_ctrl_logic/n231 [8]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  and \biu/cache_ctrl_logic/u420  (\biu/cache_ctrl_logic/n246 , \biu/cache_ctrl_logic/n55 , \biu/cache_ctrl_logic/if_l1i_chkok );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(539)
  not \biu/cache_ctrl_logic/u421  (\biu/cache_ctrl_logic/n247 , \biu/cache_ctrl_logic/ex_l1i_chkok );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(539)
  and \biu/cache_ctrl_logic/u422  (cache_ready_if, \biu/cache_ctrl_logic/n246 , \biu/cache_ctrl_logic/n247 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(539)
  not \biu/cache_ctrl_logic/u425  (\biu/cache_ctrl_logic/n248 , \biu/cache_ctrl_logic/if_l1i_chkok );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(543)
  and \biu/cache_ctrl_logic/u426  (\biu/cache_ctrl_logic/n249 , \biu/cache_ctrl_logic/if_l1i_hit , \biu/cache_ctrl_logic/n248 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(543)
  or \biu/cache_ctrl_logic/u427  (ins_page_fault, \biu/cache_ctrl_logic/n106 , \biu/cache_ctrl_logic/n249 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(543)
  and \biu/cache_ctrl_logic/u43  (\biu/cache_ctrl_logic/n25 , \biu/cache_ctrl_logic/n24 , \biu/cache_ctrl_logic/n18 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(202)
  and \biu/cache_ctrl_logic/u431  (\biu/cache_ctrl_logic/n250 , \biu/cache_ctrl_logic/ex_l1i_hit , \biu/cache_ctrl_logic/n247 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(546)
  or \biu/cache_ctrl_logic/u432  (\biu/cache_ctrl_logic/n251 , \biu/cache_ctrl_logic/n107 , \biu/cache_ctrl_logic/n250 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(546)
  and \biu/cache_ctrl_logic/u434  (\biu/cache_ctrl_logic/n252 , \biu/cache_ctrl_logic/ex_l1d_hit , \biu/cache_ctrl_logic/n198 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(546)
  or \biu/cache_ctrl_logic/u435  (store_page_fault, \biu/cache_ctrl_logic/n251 , \biu/cache_ctrl_logic/n252 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(546)
  or \biu/cache_ctrl_logic/u44  (\biu/cache_ctrl_logic/n26 , \biu/cache_ctrl_logic/n19 , \biu/cache_ctrl_logic/n25 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(202)
  or \biu/cache_ctrl_logic/u440  (\biu/cache_ctrl_logic/n253 , \biu/cache_ctrl_logic/n108 , \biu/cache_ctrl_logic/n250 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(549)
  or \biu/cache_ctrl_logic/u443  (load_page_fault, \biu/cache_ctrl_logic/n253 , \biu/cache_ctrl_logic/n252 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(549)
  or \biu/cache_ctrl_logic/u444  (\biu/cache_ctrl_logic/n232 [63], \biu/cache_ctrl_logic/n230 [63], \biu/cache_ctrl_logic/n231 [63]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u445  (\biu/cache_ctrl_logic/n230 [1], \biu/cache_ctrl_logic/n228 [1], \biu/cache_ctrl_logic/n229 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u446  (\biu/cache_ctrl_logic/n230 [2], \biu/cache_ctrl_logic/n228 [2], \biu/cache_ctrl_logic/n229 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u447  (\biu/cache_ctrl_logic/n230 [3], \biu/cache_ctrl_logic/n228 [3], \biu/cache_ctrl_logic/n229 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u448  (\biu/cache_ctrl_logic/n230 [4], \biu/cache_ctrl_logic/n228 [4], \biu/cache_ctrl_logic/n229 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u449  (\biu/cache_ctrl_logic/n230 [5], \biu/cache_ctrl_logic/n228 [5], \biu/cache_ctrl_logic/n229 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u45  (\biu/cache_ctrl_logic/n28 , \biu/cache_ctrl_logic/n26 , \biu/cache_ctrl_logic/n27 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(203)
  or \biu/cache_ctrl_logic/u450  (\biu/cache_ctrl_logic/n230 [6], \biu/cache_ctrl_logic/n228 [6], \biu/cache_ctrl_logic/n229 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u451  (\biu/cache_ctrl_logic/n230 [7], \biu/cache_ctrl_logic/n228 [7], \biu/cache_ctrl_logic/n229 [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u452  (\biu/cache_ctrl_logic/n230 [8], \biu/cache_ctrl_logic/n228 [8], \biu/cache_ctrl_logic/n229 [8]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u453  (\biu/cache_ctrl_logic/n230 [9], \biu/cache_ctrl_logic/n228 [9], \biu/cache_ctrl_logic/n229 [9]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u454  (\biu/cache_ctrl_logic/n230 [10], \biu/cache_ctrl_logic/n228 [10], \biu/cache_ctrl_logic/n229 [10]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u455  (\biu/cache_ctrl_logic/n230 [11], \biu/cache_ctrl_logic/n228 [11], \biu/cache_ctrl_logic/n229 [11]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u456  (\biu/cache_ctrl_logic/n230 [12], \biu/cache_ctrl_logic/n228 [12], \biu/cache_ctrl_logic/n229 [12]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u457  (\biu/cache_ctrl_logic/n230 [13], \biu/cache_ctrl_logic/n228 [13], \biu/cache_ctrl_logic/n229 [13]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u458  (\biu/cache_ctrl_logic/n230 [14], \biu/cache_ctrl_logic/n228 [14], \biu/cache_ctrl_logic/n229 [14]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u459  (\biu/cache_ctrl_logic/n230 [15], \biu/cache_ctrl_logic/n228 [15], \biu/cache_ctrl_logic/n229 [15]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u46  (\biu/cache_ctrl_logic/n29 , \biu/cache_ctrl_logic/n28 , \biu/bus_unit/mmu/n31 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(203)
  or \biu/cache_ctrl_logic/u460  (\biu/cache_ctrl_logic/n230 [16], \biu/cache_ctrl_logic/n228 [16], \biu/cache_ctrl_logic/n229 [16]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u461  (\biu/cache_ctrl_logic/n230 [17], \biu/cache_ctrl_logic/n228 [17], \biu/cache_ctrl_logic/n229 [17]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u462  (\biu/cache_ctrl_logic/n230 [18], \biu/cache_ctrl_logic/n228 [18], \biu/cache_ctrl_logic/n229 [18]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u463  (\biu/cache_ctrl_logic/n230 [19], \biu/cache_ctrl_logic/n228 [19], \biu/cache_ctrl_logic/n229 [19]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u464  (\biu/cache_ctrl_logic/n230 [20], \biu/cache_ctrl_logic/n228 [20], \biu/cache_ctrl_logic/n229 [20]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u465  (\biu/cache_ctrl_logic/n230 [21], \biu/cache_ctrl_logic/n228 [21], \biu/cache_ctrl_logic/n229 [21]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u466  (\biu/cache_ctrl_logic/n230 [22], \biu/cache_ctrl_logic/n228 [22], \biu/cache_ctrl_logic/n229 [22]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u467  (\biu/cache_ctrl_logic/n230 [23], \biu/cache_ctrl_logic/n228 [23], \biu/cache_ctrl_logic/n229 [23]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u468  (\biu/cache_ctrl_logic/n230 [24], \biu/cache_ctrl_logic/n228 [24], \biu/cache_ctrl_logic/n229 [24]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u469  (\biu/cache_ctrl_logic/n230 [25], \biu/cache_ctrl_logic/n228 [25], \biu/cache_ctrl_logic/n229 [25]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  and \biu/cache_ctrl_logic/u47  (\biu/cache_ctrl_logic/ex_l1i_chkok , \biu/cache_ctrl_logic/ex_l1i_hit , \biu/cache_ctrl_logic/n29 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(203)
  or \biu/cache_ctrl_logic/u470  (\biu/cache_ctrl_logic/n230 [26], \biu/cache_ctrl_logic/n228 [26], \biu/cache_ctrl_logic/n229 [26]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u471  (\biu/cache_ctrl_logic/n230 [27], \biu/cache_ctrl_logic/n228 [27], \biu/cache_ctrl_logic/n229 [27]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u472  (\biu/cache_ctrl_logic/n230 [28], \biu/cache_ctrl_logic/n228 [28], \biu/cache_ctrl_logic/n229 [28]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u473  (\biu/cache_ctrl_logic/n230 [29], \biu/cache_ctrl_logic/n228 [29], \biu/cache_ctrl_logic/n229 [29]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u474  (\biu/cache_ctrl_logic/n230 [30], \biu/cache_ctrl_logic/n228 [30], \biu/cache_ctrl_logic/n229 [30]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u475  (\biu/cache_ctrl_logic/n230 [31], \biu/cache_ctrl_logic/n228 [31], \biu/cache_ctrl_logic/n229 [31]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u476  (\biu/cache_ctrl_logic/n230 [32], \biu/cache_ctrl_logic/n228 [32], \biu/cache_ctrl_logic/n229 [32]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u477  (\biu/cache_ctrl_logic/n230 [33], \biu/cache_ctrl_logic/n228 [33], \biu/cache_ctrl_logic/n229 [33]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u478  (\biu/cache_ctrl_logic/n230 [34], \biu/cache_ctrl_logic/n228 [34], \biu/cache_ctrl_logic/n229 [34]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u479  (\biu/cache_ctrl_logic/n230 [35], \biu/cache_ctrl_logic/n228 [35], \biu/cache_ctrl_logic/n229 [35]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u48  (\biu/cache_ctrl_logic/n232 [7], \biu/cache_ctrl_logic/n230 [7], \biu/cache_ctrl_logic/n231 [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u480  (\biu/cache_ctrl_logic/n230 [36], \biu/cache_ctrl_logic/n228 [36], \biu/cache_ctrl_logic/n229 [36]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u481  (\biu/cache_ctrl_logic/n230 [37], \biu/cache_ctrl_logic/n228 [37], \biu/cache_ctrl_logic/n229 [37]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u482  (\biu/cache_ctrl_logic/n230 [38], \biu/cache_ctrl_logic/n228 [38], \biu/cache_ctrl_logic/n229 [38]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u483  (\biu/cache_ctrl_logic/n230 [39], \biu/cache_ctrl_logic/n228 [39], \biu/cache_ctrl_logic/n229 [39]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u484  (\biu/cache_ctrl_logic/n230 [40], \biu/cache_ctrl_logic/n228 [40], \biu/cache_ctrl_logic/n229 [40]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u485  (\biu/cache_ctrl_logic/n230 [41], \biu/cache_ctrl_logic/n228 [41], \biu/cache_ctrl_logic/n229 [41]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u486  (\biu/cache_ctrl_logic/n230 [42], \biu/cache_ctrl_logic/n228 [42], \biu/cache_ctrl_logic/n229 [42]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u487  (\biu/cache_ctrl_logic/n230 [43], \biu/cache_ctrl_logic/n228 [43], \biu/cache_ctrl_logic/n229 [43]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u488  (\biu/cache_ctrl_logic/n230 [44], \biu/cache_ctrl_logic/n228 [44], \biu/cache_ctrl_logic/n229 [44]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u489  (\biu/cache_ctrl_logic/n230 [45], \biu/cache_ctrl_logic/n228 [45], \biu/cache_ctrl_logic/n229 [45]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  and \biu/cache_ctrl_logic/u49  (\biu/cache_ctrl_logic/n30 , \biu/cache_ctrl_logic/n12 , \biu/cache_ctrl_logic/l1d_pte [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(204)
  or \biu/cache_ctrl_logic/u490  (\biu/cache_ctrl_logic/n230 [46], \biu/cache_ctrl_logic/n228 [46], \biu/cache_ctrl_logic/n229 [46]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u491  (\biu/cache_ctrl_logic/n230 [47], \biu/cache_ctrl_logic/n228 [47], \biu/cache_ctrl_logic/n229 [47]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u492  (\biu/cache_ctrl_logic/n230 [48], \biu/cache_ctrl_logic/n228 [48], \biu/cache_ctrl_logic/n229 [48]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u493  (\biu/cache_ctrl_logic/n230 [49], \biu/cache_ctrl_logic/n228 [49], \biu/cache_ctrl_logic/n229 [49]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u494  (\biu/cache_ctrl_logic/n230 [50], \biu/cache_ctrl_logic/n228 [50], \biu/cache_ctrl_logic/n229 [50]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u495  (\biu/cache_ctrl_logic/n230 [51], \biu/cache_ctrl_logic/n228 [51], \biu/cache_ctrl_logic/n229 [51]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u496  (\biu/cache_ctrl_logic/n230 [52], \biu/cache_ctrl_logic/n228 [52], \biu/cache_ctrl_logic/n229 [52]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u497  (\biu/cache_ctrl_logic/n230 [53], \biu/cache_ctrl_logic/n228 [53], \biu/cache_ctrl_logic/n229 [53]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u498  (\biu/cache_ctrl_logic/n230 [54], \biu/cache_ctrl_logic/n228 [54], \biu/cache_ctrl_logic/n229 [54]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u499  (\biu/cache_ctrl_logic/n230 [55], \biu/cache_ctrl_logic/n228 [55], \biu/cache_ctrl_logic/n229 [55]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  not \biu/cache_ctrl_logic/u5  (\biu/cache_ctrl_logic/n0 , \biu/cache_ctrl_logic/l1i_pte [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(180)
  and \biu/cache_ctrl_logic/u50  (\biu/cache_ctrl_logic/n31 , write, \biu/cache_ctrl_logic/l1d_pte [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(204)
  or \biu/cache_ctrl_logic/u500  (\biu/cache_ctrl_logic/n230 [56], \biu/cache_ctrl_logic/n228 [56], \biu/cache_ctrl_logic/n229 [56]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u501  (\biu/cache_ctrl_logic/n230 [57], \biu/cache_ctrl_logic/n228 [57], \biu/cache_ctrl_logic/n229 [57]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u502  (\biu/cache_ctrl_logic/n230 [58], \biu/cache_ctrl_logic/n228 [58], \biu/cache_ctrl_logic/n229 [58]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u503  (\biu/cache_ctrl_logic/n230 [59], \biu/cache_ctrl_logic/n228 [59], \biu/cache_ctrl_logic/n229 [59]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u504  (\biu/cache_ctrl_logic/n230 [60], \biu/cache_ctrl_logic/n228 [60], \biu/cache_ctrl_logic/n229 [60]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u505  (\biu/cache_ctrl_logic/n230 [61], \biu/cache_ctrl_logic/n228 [61], \biu/cache_ctrl_logic/n229 [61]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u506  (\biu/cache_ctrl_logic/n230 [62], \biu/cache_ctrl_logic/n228 [62], \biu/cache_ctrl_logic/n229 [62]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u507  (\biu/cache_ctrl_logic/n230 [63], \biu/cache_ctrl_logic/n228 [63], \biu/cache_ctrl_logic/n229 [63]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(518)
  or \biu/cache_ctrl_logic/u508  (\biu/maddress [1], \biu/cache_ctrl_logic/n222 [1], \biu/cache_ctrl_logic/n223 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u509  (\biu/maddress [2], \biu/cache_ctrl_logic/n222 [2], \biu/cache_ctrl_logic/n223 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  and \biu/cache_ctrl_logic/u51  (\biu/cache_ctrl_logic/n32 , mxr, \biu/cache_ctrl_logic/l1d_pte [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(204)
  or \biu/cache_ctrl_logic/u510  (\biu/maddress [3], \biu/cache_ctrl_logic/n222 [3], \biu/cache_ctrl_logic/n223 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u511  (\biu/maddress [4], \biu/cache_ctrl_logic/n222 [4], \biu/cache_ctrl_logic/n223 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u512  (\biu/maddress [5], \biu/cache_ctrl_logic/n222 [5], \biu/cache_ctrl_logic/n223 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u513  (\biu/maddress [6], \biu/cache_ctrl_logic/n222 [6], \biu/cache_ctrl_logic/n223 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u514  (\biu/maddress [7], \biu/cache_ctrl_logic/n222 [7], \biu/cache_ctrl_logic/n223 [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u515  (\biu/maddress [8], \biu/cache_ctrl_logic/n222 [8], \biu/cache_ctrl_logic/n223 [8]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u516  (\biu/maddress [9], \biu/cache_ctrl_logic/n222 [9], \biu/cache_ctrl_logic/n223 [9]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u517  (\biu/maddress [10], \biu/cache_ctrl_logic/n222 [10], \biu/cache_ctrl_logic/n223 [10]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u518  (\biu/maddress [11], \biu/cache_ctrl_logic/n222 [11], \biu/cache_ctrl_logic/n223 [11]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u519  (\biu/maddress [12], \biu/cache_ctrl_logic/n222 [12], \biu/cache_ctrl_logic/n223 [12]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u52  (\biu/cache_ctrl_logic/n33 , \biu/cache_ctrl_logic/l1d_pte [1], \biu/cache_ctrl_logic/n32 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(204)
  or \biu/cache_ctrl_logic/u520  (\biu/maddress [13], \biu/cache_ctrl_logic/n222 [13], \biu/cache_ctrl_logic/n223 [13]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u521  (\biu/maddress [14], \biu/cache_ctrl_logic/n222 [14], \biu/cache_ctrl_logic/n223 [14]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u522  (\biu/maddress [15], \biu/cache_ctrl_logic/n222 [15], \biu/cache_ctrl_logic/n223 [15]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u523  (\biu/maddress [16], \biu/cache_ctrl_logic/n222 [16], \biu/cache_ctrl_logic/n223 [16]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u524  (\biu/maddress [17], \biu/cache_ctrl_logic/n222 [17], \biu/cache_ctrl_logic/n223 [17]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u525  (\biu/maddress [18], \biu/cache_ctrl_logic/n222 [18], \biu/cache_ctrl_logic/n223 [18]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u526  (\biu/maddress [19], \biu/cache_ctrl_logic/n222 [19], \biu/cache_ctrl_logic/n223 [19]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u527  (\biu/maddress [20], \biu/cache_ctrl_logic/n222 [20], \biu/cache_ctrl_logic/n223 [20]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u528  (\biu/maddress [21], \biu/cache_ctrl_logic/n222 [21], \biu/cache_ctrl_logic/n223 [21]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u529  (\biu/maddress [22], \biu/cache_ctrl_logic/n222 [22], \biu/cache_ctrl_logic/n223 [22]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  and \biu/cache_ctrl_logic/u53  (\biu/cache_ctrl_logic/n34 , read, \biu/cache_ctrl_logic/n33 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(204)
  or \biu/cache_ctrl_logic/u530  (\biu/maddress [23], \biu/cache_ctrl_logic/n222 [23], \biu/cache_ctrl_logic/n223 [23]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u531  (\biu/maddress [24], \biu/cache_ctrl_logic/n222 [24], \biu/cache_ctrl_logic/n223 [24]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u532  (\biu/maddress [25], \biu/cache_ctrl_logic/n222 [25], \biu/cache_ctrl_logic/n223 [25]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u533  (\biu/maddress [26], \biu/cache_ctrl_logic/n222 [26], \biu/cache_ctrl_logic/n223 [26]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u534  (\biu/maddress [27], \biu/cache_ctrl_logic/n222 [27], \biu/cache_ctrl_logic/n223 [27]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u535  (\biu/maddress [28], \biu/cache_ctrl_logic/n222 [28], \biu/cache_ctrl_logic/n223 [28]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u536  (\biu/maddress [29], \biu/cache_ctrl_logic/n222 [29], \biu/cache_ctrl_logic/n223 [29]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u537  (\biu/maddress [30], \biu/cache_ctrl_logic/n222 [30], \biu/cache_ctrl_logic/n223 [30]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u538  (\biu/maddress [31], \biu/cache_ctrl_logic/n222 [31], \biu/cache_ctrl_logic/n223 [31]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u539  (\biu/maddress [32], \biu/cache_ctrl_logic/n222 [32], \biu/cache_ctrl_logic/n223 [32]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u54  (\biu/cache_ctrl_logic/n35 , \biu/cache_ctrl_logic/n31 , \biu/cache_ctrl_logic/n34 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(204)
  or \biu/cache_ctrl_logic/u540  (\biu/maddress [33], \biu/cache_ctrl_logic/n222 [33], \biu/cache_ctrl_logic/n223 [33]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u541  (\biu/maddress [34], \biu/cache_ctrl_logic/n222 [34], \biu/cache_ctrl_logic/n223 [34]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u542  (\biu/maddress [35], \biu/cache_ctrl_logic/n222 [35], \biu/cache_ctrl_logic/n223 [35]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u543  (\biu/maddress [36], \biu/cache_ctrl_logic/n222 [36], \biu/cache_ctrl_logic/n223 [36]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u544  (\biu/maddress [37], \biu/cache_ctrl_logic/n222 [37], \biu/cache_ctrl_logic/n223 [37]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u545  (\biu/maddress [38], \biu/cache_ctrl_logic/n222 [38], \biu/cache_ctrl_logic/n223 [38]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u546  (\biu/maddress [39], \biu/cache_ctrl_logic/n222 [39], \biu/cache_ctrl_logic/n223 [39]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u547  (\biu/maddress [40], \biu/cache_ctrl_logic/n222 [40], \biu/cache_ctrl_logic/n223 [40]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u548  (\biu/maddress [41], \biu/cache_ctrl_logic/n222 [41], \biu/cache_ctrl_logic/n223 [41]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u549  (\biu/maddress [42], \biu/cache_ctrl_logic/n222 [42], \biu/cache_ctrl_logic/n223 [42]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  and \biu/cache_ctrl_logic/u55  (\biu/cache_ctrl_logic/n36 , \biu/cache_ctrl_logic/n30 , \biu/cache_ctrl_logic/n35 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(204)
  or \biu/cache_ctrl_logic/u550  (\biu/maddress [43], \biu/cache_ctrl_logic/n222 [43], \biu/cache_ctrl_logic/n223 [43]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u551  (\biu/maddress [44], \biu/cache_ctrl_logic/n222 [44], \biu/cache_ctrl_logic/n223 [44]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u552  (\biu/maddress [45], \biu/cache_ctrl_logic/n222 [45], \biu/cache_ctrl_logic/n223 [45]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u553  (\biu/maddress [46], \biu/cache_ctrl_logic/n222 [46], \biu/cache_ctrl_logic/n223 [46]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u554  (\biu/maddress [47], \biu/cache_ctrl_logic/n222 [47], \biu/cache_ctrl_logic/n223 [47]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u555  (\biu/maddress [48], \biu/cache_ctrl_logic/n222 [48], \biu/cache_ctrl_logic/n223 [48]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u556  (\biu/maddress [49], \biu/cache_ctrl_logic/n222 [49], \biu/cache_ctrl_logic/n223 [49]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u557  (\biu/maddress [50], \biu/cache_ctrl_logic/n222 [50], \biu/cache_ctrl_logic/n223 [50]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u558  (\biu/maddress [51], \biu/cache_ctrl_logic/n222 [51], \biu/cache_ctrl_logic/n223 [51]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u559  (\biu/maddress [52], \biu/cache_ctrl_logic/n222 [52], \biu/cache_ctrl_logic/n223 [52]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u56  (\biu/cache_ctrl_logic/n232 [6], \biu/cache_ctrl_logic/n230 [6], \biu/cache_ctrl_logic/n231 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u560  (\biu/maddress [53], \biu/cache_ctrl_logic/n222 [53], \biu/cache_ctrl_logic/n223 [53]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u561  (\biu/maddress [54], \biu/cache_ctrl_logic/n222 [54], \biu/cache_ctrl_logic/n223 [54]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u562  (\biu/maddress [55], \biu/cache_ctrl_logic/n222 [55], \biu/cache_ctrl_logic/n223 [55]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u563  (\biu/maddress [56], \biu/cache_ctrl_logic/n222 [56], \biu/cache_ctrl_logic/n223 [56]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u564  (\biu/maddress [57], \biu/cache_ctrl_logic/n222 [57], \biu/cache_ctrl_logic/n223 [57]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u565  (\biu/maddress [58], \biu/cache_ctrl_logic/n222 [58], \biu/cache_ctrl_logic/n223 [58]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u566  (\biu/maddress [59], \biu/cache_ctrl_logic/n222 [59], \biu/cache_ctrl_logic/n223 [59]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u567  (\biu/maddress [60], \biu/cache_ctrl_logic/n222 [60], \biu/cache_ctrl_logic/n223 [60]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u568  (\biu/maddress [61], \biu/cache_ctrl_logic/n222 [61], \biu/cache_ctrl_logic/n223 [61]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u569  (\biu/maddress [62], \biu/cache_ctrl_logic/n222 [62], \biu/cache_ctrl_logic/n223 [62]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  and \biu/cache_ctrl_logic/u57  (\biu/cache_ctrl_logic/n37 , sum, \biu/cache_ctrl_logic/l1d_pte [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(205)
  or \biu/cache_ctrl_logic/u570  (\biu/maddress [63], \biu/cache_ctrl_logic/n222 [63], \biu/cache_ctrl_logic/n223 [63]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(510)
  or \biu/cache_ctrl_logic/u571  (\biu/cache_ctrl_logic/n222 [1], \biu/cache_ctrl_logic/n220 [1], \biu/cache_ctrl_logic/n221 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u572  (\biu/cache_ctrl_logic/n222 [2], \biu/cache_ctrl_logic/n220 [2], \biu/cache_ctrl_logic/n221 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u573  (\biu/cache_ctrl_logic/n222 [3], \biu/cache_ctrl_logic/n220 [3], \biu/cache_ctrl_logic/n221 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u574  (\biu/cache_ctrl_logic/n222 [4], \biu/cache_ctrl_logic/n220 [4], \biu/cache_ctrl_logic/n221 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u575  (\biu/cache_ctrl_logic/n222 [5], \biu/cache_ctrl_logic/n220 [5], \biu/cache_ctrl_logic/n221 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u576  (\biu/cache_ctrl_logic/n222 [6], \biu/cache_ctrl_logic/n220 [6], \biu/cache_ctrl_logic/n221 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u577  (\biu/cache_ctrl_logic/n222 [7], \biu/cache_ctrl_logic/n220 [7], \biu/cache_ctrl_logic/n221 [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u578  (\biu/cache_ctrl_logic/n222 [8], \biu/cache_ctrl_logic/n220 [8], \biu/cache_ctrl_logic/n221 [8]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u579  (\biu/cache_ctrl_logic/n222 [9], \biu/cache_ctrl_logic/n220 [9], \biu/cache_ctrl_logic/n221 [9]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  not \biu/cache_ctrl_logic/u58  (\biu/cache_ctrl_logic/n38 , \biu/cache_ctrl_logic/l1d_pte [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(205)
  or \biu/cache_ctrl_logic/u580  (\biu/cache_ctrl_logic/n222 [10], \biu/cache_ctrl_logic/n220 [10], \biu/cache_ctrl_logic/n221 [10]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u581  (\biu/cache_ctrl_logic/n222 [11], \biu/cache_ctrl_logic/n220 [11], \biu/cache_ctrl_logic/n221 [11]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u582  (\biu/cache_ctrl_logic/n222 [12], \biu/cache_ctrl_logic/n220 [12], \biu/cache_ctrl_logic/n221 [12]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u583  (\biu/cache_ctrl_logic/n222 [13], \biu/cache_ctrl_logic/n220 [13], \biu/cache_ctrl_logic/n221 [13]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u584  (\biu/cache_ctrl_logic/n222 [14], \biu/cache_ctrl_logic/n220 [14], \biu/cache_ctrl_logic/n221 [14]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u585  (\biu/cache_ctrl_logic/n222 [15], \biu/cache_ctrl_logic/n220 [15], \biu/cache_ctrl_logic/n221 [15]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u586  (\biu/cache_ctrl_logic/n222 [16], \biu/cache_ctrl_logic/n220 [16], \biu/cache_ctrl_logic/n221 [16]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u587  (\biu/cache_ctrl_logic/n222 [17], \biu/cache_ctrl_logic/n220 [17], \biu/cache_ctrl_logic/n221 [17]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u588  (\biu/cache_ctrl_logic/n222 [18], \biu/cache_ctrl_logic/n220 [18], \biu/cache_ctrl_logic/n221 [18]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u589  (\biu/cache_ctrl_logic/n222 [19], \biu/cache_ctrl_logic/n220 [19], \biu/cache_ctrl_logic/n221 [19]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u59  (\biu/cache_ctrl_logic/n39 , \biu/cache_ctrl_logic/n37 , \biu/cache_ctrl_logic/n38 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(205)
  or \biu/cache_ctrl_logic/u590  (\biu/cache_ctrl_logic/n222 [20], \biu/cache_ctrl_logic/n220 [20], \biu/cache_ctrl_logic/n221 [20]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u591  (\biu/cache_ctrl_logic/n222 [21], \biu/cache_ctrl_logic/n220 [21], \biu/cache_ctrl_logic/n221 [21]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u592  (\biu/cache_ctrl_logic/n222 [22], \biu/cache_ctrl_logic/n220 [22], \biu/cache_ctrl_logic/n221 [22]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u593  (\biu/cache_ctrl_logic/n222 [23], \biu/cache_ctrl_logic/n220 [23], \biu/cache_ctrl_logic/n221 [23]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u594  (\biu/cache_ctrl_logic/n222 [24], \biu/cache_ctrl_logic/n220 [24], \biu/cache_ctrl_logic/n221 [24]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u595  (\biu/cache_ctrl_logic/n222 [25], \biu/cache_ctrl_logic/n220 [25], \biu/cache_ctrl_logic/n221 [25]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u596  (\biu/cache_ctrl_logic/n222 [26], \biu/cache_ctrl_logic/n220 [26], \biu/cache_ctrl_logic/n221 [26]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u597  (\biu/cache_ctrl_logic/n222 [27], \biu/cache_ctrl_logic/n220 [27], \biu/cache_ctrl_logic/n221 [27]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u598  (\biu/cache_ctrl_logic/n222 [28], \biu/cache_ctrl_logic/n220 [28], \biu/cache_ctrl_logic/n221 [28]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u599  (\biu/cache_ctrl_logic/n222 [29], \biu/cache_ctrl_logic/n220 [29], \biu/cache_ctrl_logic/n221 [29]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  and \biu/cache_ctrl_logic/u6  (\biu/cache_ctrl_logic/pte_l1i_upd , \biu/cache_ctrl_logic/l1i_write_through , \biu/cache_ctrl_logic/n0 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(180)
  and \biu/cache_ctrl_logic/u60  (\biu/cache_ctrl_logic/n40 , \biu/cache_ctrl_logic/n20 , \biu/cache_ctrl_logic/n39 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(205)
  or \biu/cache_ctrl_logic/u600  (\biu/cache_ctrl_logic/n222 [30], \biu/cache_ctrl_logic/n220 [30], \biu/cache_ctrl_logic/n221 [30]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u601  (\biu/cache_ctrl_logic/n222 [31], \biu/cache_ctrl_logic/n220 [31], \biu/cache_ctrl_logic/n221 [31]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u602  (\biu/cache_ctrl_logic/n222 [32], \biu/cache_ctrl_logic/n220 [32], \biu/cache_ctrl_logic/n221 [32]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u603  (\biu/cache_ctrl_logic/n222 [33], \biu/cache_ctrl_logic/n220 [33], \biu/cache_ctrl_logic/n221 [33]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u604  (\biu/cache_ctrl_logic/n222 [34], \biu/cache_ctrl_logic/n220 [34], \biu/cache_ctrl_logic/n221 [34]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u605  (\biu/cache_ctrl_logic/n222 [35], \biu/cache_ctrl_logic/n220 [35], \biu/cache_ctrl_logic/n221 [35]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u606  (\biu/cache_ctrl_logic/n222 [36], \biu/cache_ctrl_logic/n220 [36], \biu/cache_ctrl_logic/n221 [36]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u607  (\biu/cache_ctrl_logic/n222 [37], \biu/cache_ctrl_logic/n220 [37], \biu/cache_ctrl_logic/n221 [37]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u608  (\biu/cache_ctrl_logic/n222 [38], \biu/cache_ctrl_logic/n220 [38], \biu/cache_ctrl_logic/n221 [38]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u609  (\biu/cache_ctrl_logic/n222 [39], \biu/cache_ctrl_logic/n220 [39], \biu/cache_ctrl_logic/n221 [39]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u61  (\biu/cache_ctrl_logic/n232 [5], \biu/cache_ctrl_logic/n230 [5], \biu/cache_ctrl_logic/n231 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u610  (\biu/cache_ctrl_logic/n222 [40], \biu/cache_ctrl_logic/n220 [40], \biu/cache_ctrl_logic/n221 [40]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u611  (\biu/cache_ctrl_logic/n222 [41], \biu/cache_ctrl_logic/n220 [41], \biu/cache_ctrl_logic/n221 [41]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u612  (\biu/cache_ctrl_logic/n222 [42], \biu/cache_ctrl_logic/n220 [42], \biu/cache_ctrl_logic/n221 [42]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u613  (\biu/cache_ctrl_logic/n222 [43], \biu/cache_ctrl_logic/n220 [43], \biu/cache_ctrl_logic/n221 [43]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u614  (\biu/cache_ctrl_logic/n222 [44], \biu/cache_ctrl_logic/n220 [44], \biu/cache_ctrl_logic/n221 [44]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u615  (\biu/cache_ctrl_logic/n222 [45], \biu/cache_ctrl_logic/n220 [45], \biu/cache_ctrl_logic/n221 [45]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u616  (\biu/cache_ctrl_logic/n222 [46], \biu/cache_ctrl_logic/n220 [46], \biu/cache_ctrl_logic/n221 [46]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u617  (\biu/cache_ctrl_logic/n222 [47], \biu/cache_ctrl_logic/n220 [47], \biu/cache_ctrl_logic/n221 [47]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u618  (\biu/cache_ctrl_logic/n222 [48], \biu/cache_ctrl_logic/n220 [48], \biu/cache_ctrl_logic/n221 [48]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u619  (\biu/cache_ctrl_logic/n222 [49], \biu/cache_ctrl_logic/n220 [49], \biu/cache_ctrl_logic/n221 [49]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u62  (\biu/cache_ctrl_logic/n232 [4], \biu/cache_ctrl_logic/n230 [4], \biu/cache_ctrl_logic/n231 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u620  (\biu/cache_ctrl_logic/n222 [50], \biu/cache_ctrl_logic/n220 [50], \biu/cache_ctrl_logic/n221 [50]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u621  (\biu/cache_ctrl_logic/n222 [51], \biu/cache_ctrl_logic/n220 [51], \biu/cache_ctrl_logic/n221 [51]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u622  (\biu/cache_ctrl_logic/n222 [52], \biu/cache_ctrl_logic/n220 [52], \biu/cache_ctrl_logic/n221 [52]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u623  (\biu/cache_ctrl_logic/n222 [53], \biu/cache_ctrl_logic/n220 [53], \biu/cache_ctrl_logic/n221 [53]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u624  (\biu/cache_ctrl_logic/n222 [54], \biu/cache_ctrl_logic/n220 [54], \biu/cache_ctrl_logic/n221 [54]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u625  (\biu/cache_ctrl_logic/n222 [55], \biu/cache_ctrl_logic/n220 [55], \biu/cache_ctrl_logic/n221 [55]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u626  (\biu/cache_ctrl_logic/n222 [56], \biu/cache_ctrl_logic/n220 [56], \biu/cache_ctrl_logic/n221 [56]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u627  (\biu/cache_ctrl_logic/n222 [57], \biu/cache_ctrl_logic/n220 [57], \biu/cache_ctrl_logic/n221 [57]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u628  (\biu/cache_ctrl_logic/n222 [58], \biu/cache_ctrl_logic/n220 [58], \biu/cache_ctrl_logic/n221 [58]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u629  (\biu/cache_ctrl_logic/n222 [59], \biu/cache_ctrl_logic/n220 [59], \biu/cache_ctrl_logic/n221 [59]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u63  (\biu/cache_ctrl_logic/n41 , \biu/cache_ctrl_logic/l1i_pte [1], \biu/cache_ctrl_logic/n32 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(205)
  or \biu/cache_ctrl_logic/u630  (\biu/cache_ctrl_logic/n222 [60], \biu/cache_ctrl_logic/n220 [60], \biu/cache_ctrl_logic/n221 [60]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u631  (\biu/cache_ctrl_logic/n222 [61], \biu/cache_ctrl_logic/n220 [61], \biu/cache_ctrl_logic/n221 [61]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u632  (\biu/cache_ctrl_logic/n222 [62], \biu/cache_ctrl_logic/n220 [62], \biu/cache_ctrl_logic/n221 [62]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u633  (\biu/cache_ctrl_logic/n222 [63], \biu/cache_ctrl_logic/n220 [63], \biu/cache_ctrl_logic/n221 [63]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(509)
  or \biu/cache_ctrl_logic/u634  (\biu/cache_ctrl_logic/n220 [1], \biu/cache_ctrl_logic/n218 [1], \biu/cache_ctrl_logic/n219 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u635  (\biu/cache_ctrl_logic/n220 [2], \biu/cache_ctrl_logic/n218 [2], \biu/cache_ctrl_logic/n219 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u636  (\biu/cache_ctrl_logic/n220 [3], \biu/cache_ctrl_logic/n218 [3], \biu/cache_ctrl_logic/n219 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u637  (\biu/cache_ctrl_logic/n220 [4], \biu/cache_ctrl_logic/n218 [4], \biu/cache_ctrl_logic/n219 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u638  (\biu/cache_ctrl_logic/n220 [5], \biu/cache_ctrl_logic/n218 [5], \biu/cache_ctrl_logic/n219 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u639  (\biu/cache_ctrl_logic/n220 [6], \biu/cache_ctrl_logic/n218 [6], \biu/cache_ctrl_logic/n219 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  and \biu/cache_ctrl_logic/u64  (\biu/cache_ctrl_logic/n42 , read, \biu/cache_ctrl_logic/n41 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(205)
  or \biu/cache_ctrl_logic/u640  (\biu/cache_ctrl_logic/n220 [7], \biu/cache_ctrl_logic/n218 [7], \biu/cache_ctrl_logic/n219 [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u641  (\biu/cache_ctrl_logic/n220 [8], \biu/cache_ctrl_logic/n218 [8], \biu/cache_ctrl_logic/n219 [8]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u642  (\biu/cache_ctrl_logic/n220 [9], \biu/cache_ctrl_logic/n218 [9], \biu/cache_ctrl_logic/n219 [9]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u643  (\biu/cache_ctrl_logic/n220 [10], \biu/cache_ctrl_logic/n218 [10], \biu/cache_ctrl_logic/n219 [10]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u644  (\biu/cache_ctrl_logic/n220 [11], \biu/cache_ctrl_logic/n218 [11], \biu/cache_ctrl_logic/n219 [11]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u645  (\biu/cache_ctrl_logic/n220 [12], \biu/cache_ctrl_logic/n218 [12], \biu/cache_ctrl_logic/n219 [12]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u646  (\biu/cache_ctrl_logic/n220 [13], \biu/cache_ctrl_logic/n218 [13], \biu/cache_ctrl_logic/n219 [13]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u647  (\biu/cache_ctrl_logic/n220 [14], \biu/cache_ctrl_logic/n218 [14], \biu/cache_ctrl_logic/n219 [14]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u648  (\biu/cache_ctrl_logic/n220 [15], \biu/cache_ctrl_logic/n218 [15], \biu/cache_ctrl_logic/n219 [15]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u649  (\biu/cache_ctrl_logic/n220 [16], \biu/cache_ctrl_logic/n218 [16], \biu/cache_ctrl_logic/n219 [16]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u65  (\biu/cache_ctrl_logic/n43 , \biu/cache_ctrl_logic/n31 , \biu/cache_ctrl_logic/n42 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(205)
  or \biu/cache_ctrl_logic/u650  (\biu/cache_ctrl_logic/n220 [17], \biu/cache_ctrl_logic/n218 [17], \biu/cache_ctrl_logic/n219 [17]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u651  (\biu/cache_ctrl_logic/n220 [18], \biu/cache_ctrl_logic/n218 [18], \biu/cache_ctrl_logic/n219 [18]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u652  (\biu/cache_ctrl_logic/n220 [19], \biu/cache_ctrl_logic/n218 [19], \biu/cache_ctrl_logic/n219 [19]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u653  (\biu/cache_ctrl_logic/n220 [20], \biu/cache_ctrl_logic/n218 [20], \biu/cache_ctrl_logic/n219 [20]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u654  (\biu/cache_ctrl_logic/n220 [21], \biu/cache_ctrl_logic/n218 [21], \biu/cache_ctrl_logic/n219 [21]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u655  (\biu/cache_ctrl_logic/n220 [22], \biu/cache_ctrl_logic/n218 [22], \biu/cache_ctrl_logic/n219 [22]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u656  (\biu/cache_ctrl_logic/n220 [23], \biu/cache_ctrl_logic/n218 [23], \biu/cache_ctrl_logic/n219 [23]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u657  (\biu/cache_ctrl_logic/n220 [24], \biu/cache_ctrl_logic/n218 [24], \biu/cache_ctrl_logic/n219 [24]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u658  (\biu/cache_ctrl_logic/n220 [25], \biu/cache_ctrl_logic/n218 [25], \biu/cache_ctrl_logic/n219 [25]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u659  (\biu/cache_ctrl_logic/n220 [26], \biu/cache_ctrl_logic/n218 [26], \biu/cache_ctrl_logic/n219 [26]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  and \biu/cache_ctrl_logic/u66  (\biu/cache_ctrl_logic/n44 , \biu/cache_ctrl_logic/n40 , \biu/cache_ctrl_logic/n43 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(205)
  or \biu/cache_ctrl_logic/u660  (\biu/cache_ctrl_logic/n220 [27], \biu/cache_ctrl_logic/n218 [27], \biu/cache_ctrl_logic/n219 [27]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u661  (\biu/cache_ctrl_logic/n220 [28], \biu/cache_ctrl_logic/n218 [28], \biu/cache_ctrl_logic/n219 [28]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u662  (\biu/cache_ctrl_logic/n220 [29], \biu/cache_ctrl_logic/n218 [29], \biu/cache_ctrl_logic/n219 [29]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u663  (\biu/cache_ctrl_logic/n220 [30], \biu/cache_ctrl_logic/n218 [30], \biu/cache_ctrl_logic/n219 [30]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u664  (\biu/cache_ctrl_logic/n220 [31], \biu/cache_ctrl_logic/n218 [31], \biu/cache_ctrl_logic/n219 [31]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u665  (\biu/cache_ctrl_logic/n220 [32], \biu/cache_ctrl_logic/n218 [32], \biu/cache_ctrl_logic/n219 [32]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u666  (\biu/cache_ctrl_logic/n220 [33], \biu/cache_ctrl_logic/n218 [33], \biu/cache_ctrl_logic/n219 [33]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u667  (\biu/cache_ctrl_logic/n220 [34], \biu/cache_ctrl_logic/n218 [34], \biu/cache_ctrl_logic/n219 [34]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u668  (\biu/cache_ctrl_logic/n220 [35], \biu/cache_ctrl_logic/n218 [35], \biu/cache_ctrl_logic/n219 [35]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u669  (\biu/cache_ctrl_logic/n220 [36], \biu/cache_ctrl_logic/n218 [36], \biu/cache_ctrl_logic/n219 [36]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u67  (\biu/cache_ctrl_logic/n45 , \biu/cache_ctrl_logic/n36 , \biu/cache_ctrl_logic/n44 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(205)
  or \biu/cache_ctrl_logic/u670  (\biu/cache_ctrl_logic/n220 [37], \biu/cache_ctrl_logic/n218 [37], \biu/cache_ctrl_logic/n219 [37]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u671  (\biu/cache_ctrl_logic/n220 [38], \biu/cache_ctrl_logic/n218 [38], \biu/cache_ctrl_logic/n219 [38]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u672  (\biu/cache_ctrl_logic/n220 [39], \biu/cache_ctrl_logic/n218 [39], \biu/cache_ctrl_logic/n219 [39]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u673  (\biu/cache_ctrl_logic/n220 [40], \biu/cache_ctrl_logic/n218 [40], \biu/cache_ctrl_logic/n219 [40]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u674  (\biu/cache_ctrl_logic/n220 [41], \biu/cache_ctrl_logic/n218 [41], \biu/cache_ctrl_logic/n219 [41]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u675  (\biu/cache_ctrl_logic/n220 [42], \biu/cache_ctrl_logic/n218 [42], \biu/cache_ctrl_logic/n219 [42]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u676  (\biu/cache_ctrl_logic/n220 [43], \biu/cache_ctrl_logic/n218 [43], \biu/cache_ctrl_logic/n219 [43]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u677  (\biu/cache_ctrl_logic/n220 [44], \biu/cache_ctrl_logic/n218 [44], \biu/cache_ctrl_logic/n219 [44]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u678  (\biu/cache_ctrl_logic/n220 [45], \biu/cache_ctrl_logic/n218 [45], \biu/cache_ctrl_logic/n219 [45]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u679  (\biu/cache_ctrl_logic/n220 [46], \biu/cache_ctrl_logic/n218 [46], \biu/cache_ctrl_logic/n219 [46]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u68  (\biu/cache_ctrl_logic/n232 [3], \biu/cache_ctrl_logic/n230 [3], \biu/cache_ctrl_logic/n231 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u680  (\biu/cache_ctrl_logic/n220 [47], \biu/cache_ctrl_logic/n218 [47], \biu/cache_ctrl_logic/n219 [47]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u681  (\biu/cache_ctrl_logic/n220 [48], \biu/cache_ctrl_logic/n218 [48], \biu/cache_ctrl_logic/n219 [48]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u682  (\biu/cache_ctrl_logic/n220 [49], \biu/cache_ctrl_logic/n218 [49], \biu/cache_ctrl_logic/n219 [49]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u683  (\biu/cache_ctrl_logic/n220 [50], \biu/cache_ctrl_logic/n218 [50], \biu/cache_ctrl_logic/n219 [50]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u684  (\biu/cache_ctrl_logic/n220 [51], \biu/cache_ctrl_logic/n218 [51], \biu/cache_ctrl_logic/n219 [51]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u685  (\biu/cache_ctrl_logic/n220 [52], \biu/cache_ctrl_logic/n218 [52], \biu/cache_ctrl_logic/n219 [52]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u686  (\biu/cache_ctrl_logic/n220 [53], \biu/cache_ctrl_logic/n218 [53], \biu/cache_ctrl_logic/n219 [53]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u687  (\biu/cache_ctrl_logic/n220 [54], \biu/cache_ctrl_logic/n218 [54], \biu/cache_ctrl_logic/n219 [54]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u688  (\biu/cache_ctrl_logic/n220 [55], \biu/cache_ctrl_logic/n218 [55], \biu/cache_ctrl_logic/n219 [55]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u689  (\biu/cache_ctrl_logic/n220 [56], \biu/cache_ctrl_logic/n218 [56], \biu/cache_ctrl_logic/n219 [56]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u69  (\biu/cache_ctrl_logic/n46 , \biu/cache_ctrl_logic/n45 , \biu/cache_ctrl_logic/n27 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(206)
  or \biu/cache_ctrl_logic/u690  (\biu/cache_ctrl_logic/n220 [57], \biu/cache_ctrl_logic/n218 [57], \biu/cache_ctrl_logic/n219 [57]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u691  (\biu/cache_ctrl_logic/n220 [58], \biu/cache_ctrl_logic/n218 [58], \biu/cache_ctrl_logic/n219 [58]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u692  (\biu/cache_ctrl_logic/n220 [59], \biu/cache_ctrl_logic/n218 [59], \biu/cache_ctrl_logic/n219 [59]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u693  (\biu/cache_ctrl_logic/n220 [60], \biu/cache_ctrl_logic/n218 [60], \biu/cache_ctrl_logic/n219 [60]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u694  (\biu/cache_ctrl_logic/n220 [61], \biu/cache_ctrl_logic/n218 [61], \biu/cache_ctrl_logic/n219 [61]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u695  (\biu/cache_ctrl_logic/n220 [62], \biu/cache_ctrl_logic/n218 [62], \biu/cache_ctrl_logic/n219 [62]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u696  (\biu/cache_ctrl_logic/n220 [63], \biu/cache_ctrl_logic/n218 [63], \biu/cache_ctrl_logic/n219 [63]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(508)
  or \biu/cache_ctrl_logic/u697  (\biu/cache_ctrl_logic/n218 [1], \biu/cache_ctrl_logic/n216 [1], \biu/cache_ctrl_logic/n217 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u698  (\biu/cache_ctrl_logic/n218 [2], \biu/cache_ctrl_logic/n216 [2], \biu/cache_ctrl_logic/n217 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u699  (\biu/cache_ctrl_logic/n218 [3], \biu/cache_ctrl_logic/n216 [3], \biu/cache_ctrl_logic/n217 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  and \biu/cache_ctrl_logic/u7  (\biu/cache_ctrl_logic/l1d_write_through , \biu/cache_ctrl_logic/ex_l1d_chkok , write);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(181)
  or \biu/cache_ctrl_logic/u70  (\biu/cache_ctrl_logic/n47 , \biu/cache_ctrl_logic/n46 , \biu/bus_unit/mmu/n31 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(206)
  or \biu/cache_ctrl_logic/u700  (\biu/cache_ctrl_logic/n218 [4], \biu/cache_ctrl_logic/n216 [4], \biu/cache_ctrl_logic/n217 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u701  (\biu/cache_ctrl_logic/n218 [5], \biu/cache_ctrl_logic/n216 [5], \biu/cache_ctrl_logic/n217 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u702  (\biu/cache_ctrl_logic/n218 [6], \biu/cache_ctrl_logic/n216 [6], \biu/cache_ctrl_logic/n217 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u703  (\biu/cache_ctrl_logic/n218 [7], \biu/cache_ctrl_logic/n216 [7], \biu/cache_ctrl_logic/n217 [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u704  (\biu/cache_ctrl_logic/n218 [8], \biu/cache_ctrl_logic/n216 [8], \biu/cache_ctrl_logic/n217 [8]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u705  (\biu/cache_ctrl_logic/n218 [9], \biu/cache_ctrl_logic/n216 [9], \biu/cache_ctrl_logic/n217 [9]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u706  (\biu/cache_ctrl_logic/n218 [10], \biu/cache_ctrl_logic/n216 [10], \biu/cache_ctrl_logic/n217 [10]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u707  (\biu/cache_ctrl_logic/n218 [11], \biu/cache_ctrl_logic/n216 [11], \biu/cache_ctrl_logic/n217 [11]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u708  (\biu/cache_ctrl_logic/n218 [12], \biu/cache_ctrl_logic/n216 [12], \biu/cache_ctrl_logic/n217 [12]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u709  (\biu/cache_ctrl_logic/n218 [13], \biu/cache_ctrl_logic/n216 [13], \biu/cache_ctrl_logic/n217 [13]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  and \biu/cache_ctrl_logic/u71  (\biu/cache_ctrl_logic/ex_l1d_chkok , \biu/cache_ctrl_logic/ex_l1d_hit , \biu/cache_ctrl_logic/n47 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(206)
  or \biu/cache_ctrl_logic/u710  (\biu/cache_ctrl_logic/n218 [14], \biu/cache_ctrl_logic/n216 [14], \biu/cache_ctrl_logic/n217 [14]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u711  (\biu/cache_ctrl_logic/n218 [15], \biu/cache_ctrl_logic/n216 [15], \biu/cache_ctrl_logic/n217 [15]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u712  (\biu/cache_ctrl_logic/n218 [16], \biu/cache_ctrl_logic/n216 [16], \biu/cache_ctrl_logic/n217 [16]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u713  (\biu/cache_ctrl_logic/n218 [17], \biu/cache_ctrl_logic/n216 [17], \biu/cache_ctrl_logic/n217 [17]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u714  (\biu/cache_ctrl_logic/n218 [18], \biu/cache_ctrl_logic/n216 [18], \biu/cache_ctrl_logic/n217 [18]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u715  (\biu/cache_ctrl_logic/n218 [19], \biu/cache_ctrl_logic/n216 [19], \biu/cache_ctrl_logic/n217 [19]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u716  (\biu/cache_ctrl_logic/n218 [20], \biu/cache_ctrl_logic/n216 [20], \biu/cache_ctrl_logic/n217 [20]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u717  (\biu/cache_ctrl_logic/n218 [21], \biu/cache_ctrl_logic/n216 [21], \biu/cache_ctrl_logic/n217 [21]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u718  (\biu/cache_ctrl_logic/n218 [22], \biu/cache_ctrl_logic/n216 [22], \biu/cache_ctrl_logic/n217 [22]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u719  (\biu/cache_ctrl_logic/n218 [23], \biu/cache_ctrl_logic/n216 [23], \biu/cache_ctrl_logic/n217 [23]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  and \biu/cache_ctrl_logic/u72  (\biu/cache_ctrl_logic/n49 , \biu/cache_ctrl_logic/n48 , \biu/cache_ctrl_logic/l1i_pte [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(207)
  or \biu/cache_ctrl_logic/u720  (\biu/cache_ctrl_logic/n218 [24], \biu/cache_ctrl_logic/n216 [24], \biu/cache_ctrl_logic/n217 [24]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u721  (\biu/cache_ctrl_logic/n218 [25], \biu/cache_ctrl_logic/n216 [25], \biu/cache_ctrl_logic/n217 [25]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u722  (\biu/cache_ctrl_logic/n218 [26], \biu/cache_ctrl_logic/n216 [26], \biu/cache_ctrl_logic/n217 [26]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u723  (\biu/cache_ctrl_logic/n218 [27], \biu/cache_ctrl_logic/n216 [27], \biu/cache_ctrl_logic/n217 [27]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u724  (\biu/cache_ctrl_logic/n218 [28], \biu/cache_ctrl_logic/n216 [28], \biu/cache_ctrl_logic/n217 [28]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u725  (\biu/cache_ctrl_logic/n218 [29], \biu/cache_ctrl_logic/n216 [29], \biu/cache_ctrl_logic/n217 [29]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u726  (\biu/cache_ctrl_logic/n218 [30], \biu/cache_ctrl_logic/n216 [30], \biu/cache_ctrl_logic/n217 [30]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u727  (\biu/cache_ctrl_logic/n218 [31], \biu/cache_ctrl_logic/n216 [31], \biu/cache_ctrl_logic/n217 [31]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u728  (\biu/cache_ctrl_logic/n218 [32], \biu/cache_ctrl_logic/n216 [32], \biu/cache_ctrl_logic/n217 [32]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u729  (\biu/cache_ctrl_logic/n218 [33], \biu/cache_ctrl_logic/n216 [33], \biu/cache_ctrl_logic/n217 [33]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u73  (\biu/cache_ctrl_logic/n51 , \biu/cache_ctrl_logic/n49 , \biu/cache_ctrl_logic/n50 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(208)
  or \biu/cache_ctrl_logic/u730  (\biu/cache_ctrl_logic/n218 [34], \biu/cache_ctrl_logic/n216 [34], \biu/cache_ctrl_logic/n217 [34]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u731  (\biu/cache_ctrl_logic/n218 [35], \biu/cache_ctrl_logic/n216 [35], \biu/cache_ctrl_logic/n217 [35]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u732  (\biu/cache_ctrl_logic/n218 [36], \biu/cache_ctrl_logic/n216 [36], \biu/cache_ctrl_logic/n217 [36]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u733  (\biu/cache_ctrl_logic/n218 [37], \biu/cache_ctrl_logic/n216 [37], \biu/cache_ctrl_logic/n217 [37]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u734  (\biu/cache_ctrl_logic/n218 [38], \biu/cache_ctrl_logic/n216 [38], \biu/cache_ctrl_logic/n217 [38]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u735  (\biu/cache_ctrl_logic/n218 [39], \biu/cache_ctrl_logic/n216 [39], \biu/cache_ctrl_logic/n217 [39]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u736  (\biu/cache_ctrl_logic/n218 [40], \biu/cache_ctrl_logic/n216 [40], \biu/cache_ctrl_logic/n217 [40]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u737  (\biu/cache_ctrl_logic/n218 [41], \biu/cache_ctrl_logic/n216 [41], \biu/cache_ctrl_logic/n217 [41]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u738  (\biu/cache_ctrl_logic/n218 [42], \biu/cache_ctrl_logic/n216 [42], \biu/cache_ctrl_logic/n217 [42]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u739  (\biu/cache_ctrl_logic/n218 [43], \biu/cache_ctrl_logic/n216 [43], \biu/cache_ctrl_logic/n217 [43]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u74  (\biu/cache_ctrl_logic/n53 , \biu/cache_ctrl_logic/n51 , \biu/cache_ctrl_logic/n52 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(209)
  or \biu/cache_ctrl_logic/u740  (\biu/cache_ctrl_logic/n218 [44], \biu/cache_ctrl_logic/n216 [44], \biu/cache_ctrl_logic/n217 [44]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u741  (\biu/cache_ctrl_logic/n218 [45], \biu/cache_ctrl_logic/n216 [45], \biu/cache_ctrl_logic/n217 [45]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u742  (\biu/cache_ctrl_logic/n218 [46], \biu/cache_ctrl_logic/n216 [46], \biu/cache_ctrl_logic/n217 [46]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u743  (\biu/cache_ctrl_logic/n218 [47], \biu/cache_ctrl_logic/n216 [47], \biu/cache_ctrl_logic/n217 [47]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u744  (\biu/cache_ctrl_logic/n218 [48], \biu/cache_ctrl_logic/n216 [48], \biu/cache_ctrl_logic/n217 [48]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u745  (\biu/cache_ctrl_logic/n218 [49], \biu/cache_ctrl_logic/n216 [49], \biu/cache_ctrl_logic/n217 [49]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u746  (\biu/cache_ctrl_logic/n218 [50], \biu/cache_ctrl_logic/n216 [50], \biu/cache_ctrl_logic/n217 [50]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u747  (\biu/cache_ctrl_logic/n218 [51], \biu/cache_ctrl_logic/n216 [51], \biu/cache_ctrl_logic/n217 [51]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u748  (\biu/cache_ctrl_logic/n218 [52], \biu/cache_ctrl_logic/n216 [52], \biu/cache_ctrl_logic/n217 [52]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u749  (\biu/cache_ctrl_logic/n218 [53], \biu/cache_ctrl_logic/n216 [53], \biu/cache_ctrl_logic/n217 [53]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u75  (\biu/cache_ctrl_logic/n54 , \biu/cache_ctrl_logic/n53 , \biu/bus_unit/mmu/n31 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(209)
  or \biu/cache_ctrl_logic/u750  (\biu/cache_ctrl_logic/n218 [54], \biu/cache_ctrl_logic/n216 [54], \biu/cache_ctrl_logic/n217 [54]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u751  (\biu/cache_ctrl_logic/n218 [55], \biu/cache_ctrl_logic/n216 [55], \biu/cache_ctrl_logic/n217 [55]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u752  (\biu/cache_ctrl_logic/n218 [56], \biu/cache_ctrl_logic/n216 [56], \biu/cache_ctrl_logic/n217 [56]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u753  (\biu/cache_ctrl_logic/n218 [57], \biu/cache_ctrl_logic/n216 [57], \biu/cache_ctrl_logic/n217 [57]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u754  (\biu/cache_ctrl_logic/n218 [58], \biu/cache_ctrl_logic/n216 [58], \biu/cache_ctrl_logic/n217 [58]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u755  (\biu/cache_ctrl_logic/n218 [59], \biu/cache_ctrl_logic/n216 [59], \biu/cache_ctrl_logic/n217 [59]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u756  (\biu/cache_ctrl_logic/n218 [60], \biu/cache_ctrl_logic/n216 [60], \biu/cache_ctrl_logic/n217 [60]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u757  (\biu/cache_ctrl_logic/n218 [61], \biu/cache_ctrl_logic/n216 [61], \biu/cache_ctrl_logic/n217 [61]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u758  (\biu/cache_ctrl_logic/n218 [62], \biu/cache_ctrl_logic/n216 [62], \biu/cache_ctrl_logic/n217 [62]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  or \biu/cache_ctrl_logic/u759  (\biu/cache_ctrl_logic/n218 [63], \biu/cache_ctrl_logic/n216 [63], \biu/cache_ctrl_logic/n217 [63]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(507)
  and \biu/cache_ctrl_logic/u76  (\biu/cache_ctrl_logic/if_l1i_chkok , \biu/cache_ctrl_logic/if_l1i_hit , \biu/cache_ctrl_logic/n54 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(209)
  or \biu/cache_ctrl_logic/u760  (\biu/cache_ctrl_logic/n216 [1], \biu/cache_ctrl_logic/n214 [1], \biu/cache_ctrl_logic/n215 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u761  (\biu/cache_ctrl_logic/n216 [2], \biu/cache_ctrl_logic/n214 [2], \biu/cache_ctrl_logic/n215 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u762  (\biu/cache_ctrl_logic/n216 [3], \biu/cache_ctrl_logic/n214 [3], \biu/cache_ctrl_logic/n215 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u763  (\biu/cache_ctrl_logic/n216 [4], \biu/cache_ctrl_logic/n214 [4], \biu/cache_ctrl_logic/n215 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u764  (\biu/cache_ctrl_logic/n216 [5], \biu/cache_ctrl_logic/n214 [5], \biu/cache_ctrl_logic/n215 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u765  (\biu/cache_ctrl_logic/n216 [6], \biu/cache_ctrl_logic/n214 [6], \biu/cache_ctrl_logic/n215 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u766  (\biu/cache_ctrl_logic/n216 [7], \biu/cache_ctrl_logic/n214 [7], \biu/cache_ctrl_logic/n215 [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u767  (\biu/cache_ctrl_logic/n216 [8], \biu/cache_ctrl_logic/n214 [8], \biu/cache_ctrl_logic/n215 [8]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u768  (\biu/cache_ctrl_logic/n216 [9], \biu/cache_ctrl_logic/n214 [9], \biu/cache_ctrl_logic/n215 [9]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u769  (\biu/cache_ctrl_logic/n216 [10], \biu/cache_ctrl_logic/n214 [10], \biu/cache_ctrl_logic/n215 [10]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  and \biu/cache_ctrl_logic/u77  (\biu/cache_ctrl_logic/n56 , \biu/cache_ctrl_logic/n55 , cache_flush_biu);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(218)
  or \biu/cache_ctrl_logic/u770  (\biu/cache_ctrl_logic/n216 [11], \biu/cache_ctrl_logic/n214 [11], \biu/cache_ctrl_logic/n215 [11]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u771  (\biu/cache_ctrl_logic/n216 [12], \biu/cache_ctrl_logic/n214 [12], \biu/cache_ctrl_logic/n215 [12]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u772  (\biu/cache_ctrl_logic/n216 [13], \biu/cache_ctrl_logic/n214 [13], \biu/cache_ctrl_logic/n215 [13]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u773  (\biu/cache_ctrl_logic/n216 [14], \biu/cache_ctrl_logic/n214 [14], \biu/cache_ctrl_logic/n215 [14]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u774  (\biu/cache_ctrl_logic/n216 [15], \biu/cache_ctrl_logic/n214 [15], \biu/cache_ctrl_logic/n215 [15]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u775  (\biu/cache_ctrl_logic/n216 [16], \biu/cache_ctrl_logic/n214 [16], \biu/cache_ctrl_logic/n215 [16]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u776  (\biu/cache_ctrl_logic/n216 [17], \biu/cache_ctrl_logic/n214 [17], \biu/cache_ctrl_logic/n215 [17]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u777  (\biu/cache_ctrl_logic/n216 [18], \biu/cache_ctrl_logic/n214 [18], \biu/cache_ctrl_logic/n215 [18]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u778  (\biu/cache_ctrl_logic/n216 [19], \biu/cache_ctrl_logic/n214 [19], \biu/cache_ctrl_logic/n215 [19]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u779  (\biu/cache_ctrl_logic/n216 [20], \biu/cache_ctrl_logic/n214 [20], \biu/cache_ctrl_logic/n215 [20]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u78  (\biu/cache_ctrl_logic/n232 [2], \biu/cache_ctrl_logic/n230 [2], \biu/cache_ctrl_logic/n231 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u780  (\biu/cache_ctrl_logic/n216 [21], \biu/cache_ctrl_logic/n214 [21], \biu/cache_ctrl_logic/n215 [21]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u781  (\biu/cache_ctrl_logic/n216 [22], \biu/cache_ctrl_logic/n214 [22], \biu/cache_ctrl_logic/n215 [22]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u782  (\biu/cache_ctrl_logic/n216 [23], \biu/cache_ctrl_logic/n214 [23], \biu/cache_ctrl_logic/n215 [23]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u783  (\biu/cache_ctrl_logic/n216 [24], \biu/cache_ctrl_logic/n214 [24], \biu/cache_ctrl_logic/n215 [24]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u784  (\biu/cache_ctrl_logic/n216 [25], \biu/cache_ctrl_logic/n214 [25], \biu/cache_ctrl_logic/n215 [25]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u785  (\biu/cache_ctrl_logic/n216 [26], \biu/cache_ctrl_logic/n214 [26], \biu/cache_ctrl_logic/n215 [26]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u786  (\biu/cache_ctrl_logic/n216 [27], \biu/cache_ctrl_logic/n214 [27], \biu/cache_ctrl_logic/n215 [27]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u787  (\biu/cache_ctrl_logic/n216 [28], \biu/cache_ctrl_logic/n214 [28], \biu/cache_ctrl_logic/n215 [28]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u788  (\biu/cache_ctrl_logic/n216 [29], \biu/cache_ctrl_logic/n214 [29], \biu/cache_ctrl_logic/n215 [29]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u789  (\biu/cache_ctrl_logic/n216 [30], \biu/cache_ctrl_logic/n214 [30], \biu/cache_ctrl_logic/n215 [30]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  and \biu/cache_ctrl_logic/u79  (\biu/cache_ctrl_logic/n57 , \biu/cache_ctrl_logic/n55 , \biu/cache_ctrl_logic/l1d_miss );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(222)
  or \biu/cache_ctrl_logic/u790  (\biu/cache_ctrl_logic/n216 [31], \biu/cache_ctrl_logic/n214 [31], \biu/cache_ctrl_logic/n215 [31]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u791  (\biu/cache_ctrl_logic/n216 [32], \biu/cache_ctrl_logic/n214 [32], \biu/cache_ctrl_logic/n215 [32]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u792  (\biu/cache_ctrl_logic/n216 [33], \biu/cache_ctrl_logic/n214 [33], \biu/cache_ctrl_logic/n215 [33]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u793  (\biu/cache_ctrl_logic/n216 [34], \biu/cache_ctrl_logic/n214 [34], \biu/cache_ctrl_logic/n215 [34]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u794  (\biu/cache_ctrl_logic/n216 [35], \biu/cache_ctrl_logic/n214 [35], \biu/cache_ctrl_logic/n215 [35]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u795  (\biu/cache_ctrl_logic/n216 [36], \biu/cache_ctrl_logic/n214 [36], \biu/cache_ctrl_logic/n215 [36]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u796  (\biu/cache_ctrl_logic/n216 [37], \biu/cache_ctrl_logic/n214 [37], \biu/cache_ctrl_logic/n215 [37]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u797  (\biu/cache_ctrl_logic/n216 [38], \biu/cache_ctrl_logic/n214 [38], \biu/cache_ctrl_logic/n215 [38]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u798  (\biu/cache_ctrl_logic/n216 [39], \biu/cache_ctrl_logic/n214 [39], \biu/cache_ctrl_logic/n215 [39]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u799  (\biu/cache_ctrl_logic/n216 [40], \biu/cache_ctrl_logic/n214 [40], \biu/cache_ctrl_logic/n215 [40]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  not \biu/cache_ctrl_logic/u8  (\biu/cache_ctrl_logic/n1 , \biu/cache_ctrl_logic/l1d_pte [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(181)
  and \biu/cache_ctrl_logic/u80  (\biu/cache_ctrl_logic/n58 , unpage, write);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(223)
  or \biu/cache_ctrl_logic/u800  (\biu/cache_ctrl_logic/n216 [41], \biu/cache_ctrl_logic/n214 [41], \biu/cache_ctrl_logic/n215 [41]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u801  (\biu/cache_ctrl_logic/n216 [42], \biu/cache_ctrl_logic/n214 [42], \biu/cache_ctrl_logic/n215 [42]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u802  (\biu/cache_ctrl_logic/n216 [43], \biu/cache_ctrl_logic/n214 [43], \biu/cache_ctrl_logic/n215 [43]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u803  (\biu/cache_ctrl_logic/n216 [44], \biu/cache_ctrl_logic/n214 [44], \biu/cache_ctrl_logic/n215 [44]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u804  (\biu/cache_ctrl_logic/n216 [45], \biu/cache_ctrl_logic/n214 [45], \biu/cache_ctrl_logic/n215 [45]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u805  (\biu/cache_ctrl_logic/n216 [46], \biu/cache_ctrl_logic/n214 [46], \biu/cache_ctrl_logic/n215 [46]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u806  (\biu/cache_ctrl_logic/n216 [47], \biu/cache_ctrl_logic/n214 [47], \biu/cache_ctrl_logic/n215 [47]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u807  (\biu/cache_ctrl_logic/n216 [48], \biu/cache_ctrl_logic/n214 [48], \biu/cache_ctrl_logic/n215 [48]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u808  (\biu/cache_ctrl_logic/n216 [49], \biu/cache_ctrl_logic/n214 [49], \biu/cache_ctrl_logic/n215 [49]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u809  (\biu/cache_ctrl_logic/n216 [50], \biu/cache_ctrl_logic/n214 [50], \biu/cache_ctrl_logic/n215 [50]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  and \biu/cache_ctrl_logic/u81  (\biu/cache_ctrl_logic/n59 , unpage, read);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(223)
  or \biu/cache_ctrl_logic/u810  (\biu/cache_ctrl_logic/n216 [51], \biu/cache_ctrl_logic/n214 [51], \biu/cache_ctrl_logic/n215 [51]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u811  (\biu/cache_ctrl_logic/n216 [52], \biu/cache_ctrl_logic/n214 [52], \biu/cache_ctrl_logic/n215 [52]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u812  (\biu/cache_ctrl_logic/n216 [53], \biu/cache_ctrl_logic/n214 [53], \biu/cache_ctrl_logic/n215 [53]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u813  (\biu/cache_ctrl_logic/n216 [54], \biu/cache_ctrl_logic/n214 [54], \biu/cache_ctrl_logic/n215 [54]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u814  (\biu/cache_ctrl_logic/n216 [55], \biu/cache_ctrl_logic/n214 [55], \biu/cache_ctrl_logic/n215 [55]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u815  (\biu/cache_ctrl_logic/n216 [56], \biu/cache_ctrl_logic/n214 [56], \biu/cache_ctrl_logic/n215 [56]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u816  (\biu/cache_ctrl_logic/n216 [57], \biu/cache_ctrl_logic/n214 [57], \biu/cache_ctrl_logic/n215 [57]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u817  (\biu/cache_ctrl_logic/n216 [58], \biu/cache_ctrl_logic/n214 [58], \biu/cache_ctrl_logic/n215 [58]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u818  (\biu/cache_ctrl_logic/n216 [59], \biu/cache_ctrl_logic/n214 [59], \biu/cache_ctrl_logic/n215 [59]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u819  (\biu/cache_ctrl_logic/n216 [60], \biu/cache_ctrl_logic/n214 [60], \biu/cache_ctrl_logic/n215 [60]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  not \biu/cache_ctrl_logic/u82  (\biu/cache_ctrl_logic/n70 [2], \biu/cache_ctrl_logic/n69 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(250)
  or \biu/cache_ctrl_logic/u820  (\biu/cache_ctrl_logic/n216 [61], \biu/cache_ctrl_logic/n214 [61], \biu/cache_ctrl_logic/n215 [61]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u821  (\biu/cache_ctrl_logic/n216 [62], \biu/cache_ctrl_logic/n214 [62], \biu/cache_ctrl_logic/n215 [62]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u822  (\biu/cache_ctrl_logic/n216 [63], \biu/cache_ctrl_logic/n214 [63], \biu/cache_ctrl_logic/n215 [63]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(506)
  or \biu/cache_ctrl_logic/u823  (\biu/cache_ctrl_logic/n214 [1], \biu/cache_ctrl_logic/n211 [1], \biu/cache_ctrl_logic/n213 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u824  (\biu/cache_ctrl_logic/n214 [2], \biu/cache_ctrl_logic/n211 [2], \biu/cache_ctrl_logic/n213 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u825  (\biu/cache_ctrl_logic/n214 [3], \biu/cache_ctrl_logic/n211 [3], \biu/cache_ctrl_logic/n213 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u826  (\biu/cache_ctrl_logic/n214 [4], \biu/cache_ctrl_logic/n211 [4], \biu/cache_ctrl_logic/n213 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u827  (\biu/cache_ctrl_logic/n214 [5], \biu/cache_ctrl_logic/n211 [5], \biu/cache_ctrl_logic/n213 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u828  (\biu/cache_ctrl_logic/n214 [6], \biu/cache_ctrl_logic/n211 [6], \biu/cache_ctrl_logic/n213 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u829  (\biu/cache_ctrl_logic/n214 [7], \biu/cache_ctrl_logic/n211 [7], \biu/cache_ctrl_logic/n213 [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u83  (\biu/cache_ctrl_logic/n232 [1], \biu/cache_ctrl_logic/n230 [1], \biu/cache_ctrl_logic/n231 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(519)
  or \biu/cache_ctrl_logic/u830  (\biu/cache_ctrl_logic/n214 [8], \biu/cache_ctrl_logic/n211 [8], \biu/cache_ctrl_logic/n213 [8]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u831  (\biu/cache_ctrl_logic/n214 [9], \biu/cache_ctrl_logic/n211 [9], \biu/cache_ctrl_logic/n213 [9]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u832  (\biu/cache_ctrl_logic/n214 [10], \biu/cache_ctrl_logic/n211 [10], \biu/cache_ctrl_logic/n213 [10]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u833  (\biu/cache_ctrl_logic/n214 [11], \biu/cache_ctrl_logic/n211 [11], \biu/cache_ctrl_logic/n213 [11]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u834  (\biu/cache_ctrl_logic/n214 [12], \biu/cache_ctrl_logic/n211 [12], \biu/cache_ctrl_logic/n213 [12]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u835  (\biu/cache_ctrl_logic/n214 [13], \biu/cache_ctrl_logic/n211 [13], \biu/cache_ctrl_logic/n213 [13]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u836  (\biu/cache_ctrl_logic/n214 [14], \biu/cache_ctrl_logic/n211 [14], \biu/cache_ctrl_logic/n213 [14]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u837  (\biu/cache_ctrl_logic/n214 [15], \biu/cache_ctrl_logic/n211 [15], \biu/cache_ctrl_logic/n213 [15]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u838  (\biu/cache_ctrl_logic/n214 [16], \biu/cache_ctrl_logic/n211 [16], \biu/cache_ctrl_logic/n213 [16]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u839  (\biu/cache_ctrl_logic/n214 [17], \biu/cache_ctrl_logic/n211 [17], \biu/cache_ctrl_logic/n213 [17]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  and \biu/cache_ctrl_logic/u84  (\biu/cache_ctrl_logic/n62 , \biu/cache_ctrl_logic/n55 , \biu/cache_ctrl_logic/l1i_miss );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(225)
  or \biu/cache_ctrl_logic/u840  (\biu/cache_ctrl_logic/n214 [18], \biu/cache_ctrl_logic/n211 [18], \biu/cache_ctrl_logic/n213 [18]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u841  (\biu/cache_ctrl_logic/n214 [19], \biu/cache_ctrl_logic/n211 [19], \biu/cache_ctrl_logic/n213 [19]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u842  (\biu/cache_ctrl_logic/n214 [20], \biu/cache_ctrl_logic/n211 [20], \biu/cache_ctrl_logic/n213 [20]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u843  (\biu/cache_ctrl_logic/n214 [21], \biu/cache_ctrl_logic/n211 [21], \biu/cache_ctrl_logic/n213 [21]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u844  (\biu/cache_ctrl_logic/n214 [22], \biu/cache_ctrl_logic/n211 [22], \biu/cache_ctrl_logic/n213 [22]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u845  (\biu/cache_ctrl_logic/n214 [23], \biu/cache_ctrl_logic/n211 [23], \biu/cache_ctrl_logic/n213 [23]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u846  (\biu/cache_ctrl_logic/n214 [24], \biu/cache_ctrl_logic/n211 [24], \biu/cache_ctrl_logic/n213 [24]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u847  (\biu/cache_ctrl_logic/n214 [25], \biu/cache_ctrl_logic/n211 [25], \biu/cache_ctrl_logic/n213 [25]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u848  (\biu/cache_ctrl_logic/n214 [26], \biu/cache_ctrl_logic/n211 [26], \biu/cache_ctrl_logic/n213 [26]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u849  (\biu/cache_ctrl_logic/n214 [27], \biu/cache_ctrl_logic/n211 [27], \biu/cache_ctrl_logic/n213 [27]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u85  (\biu/write_data [63], \biu/cache_ctrl_logic/n232 [63], \biu/cache_ctrl_logic/n233 [63]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u850  (\biu/cache_ctrl_logic/n214 [28], \biu/cache_ctrl_logic/n211 [28], \biu/cache_ctrl_logic/n213 [28]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u851  (\biu/cache_ctrl_logic/n214 [29], \biu/cache_ctrl_logic/n211 [29], \biu/cache_ctrl_logic/n213 [29]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u852  (\biu/cache_ctrl_logic/n214 [30], \biu/cache_ctrl_logic/n211 [30], \biu/cache_ctrl_logic/n213 [30]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u853  (\biu/cache_ctrl_logic/n214 [31], \biu/cache_ctrl_logic/n211 [31], \biu/cache_ctrl_logic/n213 [31]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u854  (\biu/cache_ctrl_logic/n214 [32], \biu/cache_ctrl_logic/n211 [32], \biu/cache_ctrl_logic/n213 [32]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u855  (\biu/cache_ctrl_logic/n214 [33], \biu/cache_ctrl_logic/n211 [33], \biu/cache_ctrl_logic/n213 [33]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u856  (\biu/cache_ctrl_logic/n214 [34], \biu/cache_ctrl_logic/n211 [34], \biu/cache_ctrl_logic/n213 [34]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u857  (\biu/cache_ctrl_logic/n214 [35], \biu/cache_ctrl_logic/n211 [35], \biu/cache_ctrl_logic/n213 [35]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u858  (\biu/cache_ctrl_logic/n214 [36], \biu/cache_ctrl_logic/n211 [36], \biu/cache_ctrl_logic/n213 [36]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u859  (\biu/cache_ctrl_logic/n214 [37], \biu/cache_ctrl_logic/n211 [37], \biu/cache_ctrl_logic/n213 [37]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  and \biu/cache_ctrl_logic/u86  (\biu/cache_ctrl_logic/n63 , \biu/cache_ctrl_logic/n55 , \biu/cache_ctrl_logic/pte_l1d_upd );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(228)
  or \biu/cache_ctrl_logic/u860  (\biu/cache_ctrl_logic/n214 [38], \biu/cache_ctrl_logic/n211 [38], \biu/cache_ctrl_logic/n213 [38]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u861  (\biu/cache_ctrl_logic/n214 [39], \biu/cache_ctrl_logic/n211 [39], \biu/cache_ctrl_logic/n213 [39]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u862  (\biu/cache_ctrl_logic/n214 [40], \biu/cache_ctrl_logic/n211 [40], \biu/cache_ctrl_logic/n213 [40]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u863  (\biu/cache_ctrl_logic/n214 [41], \biu/cache_ctrl_logic/n211 [41], \biu/cache_ctrl_logic/n213 [41]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u864  (\biu/cache_ctrl_logic/n214 [42], \biu/cache_ctrl_logic/n211 [42], \biu/cache_ctrl_logic/n213 [42]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u865  (\biu/cache_ctrl_logic/n214 [43], \biu/cache_ctrl_logic/n211 [43], \biu/cache_ctrl_logic/n213 [43]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u866  (\biu/cache_ctrl_logic/n214 [44], \biu/cache_ctrl_logic/n211 [44], \biu/cache_ctrl_logic/n213 [44]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u867  (\biu/cache_ctrl_logic/n214 [45], \biu/cache_ctrl_logic/n211 [45], \biu/cache_ctrl_logic/n213 [45]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u868  (\biu/cache_ctrl_logic/n214 [46], \biu/cache_ctrl_logic/n211 [46], \biu/cache_ctrl_logic/n213 [46]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u869  (\biu/cache_ctrl_logic/n214 [47], \biu/cache_ctrl_logic/n211 [47], \biu/cache_ctrl_logic/n213 [47]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u87  (\biu/write_data [62], \biu/cache_ctrl_logic/n232 [62], \biu/cache_ctrl_logic/n233 [62]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u870  (\biu/cache_ctrl_logic/n214 [48], \biu/cache_ctrl_logic/n211 [48], \biu/cache_ctrl_logic/n213 [48]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u871  (\biu/cache_ctrl_logic/n214 [49], \biu/cache_ctrl_logic/n211 [49], \biu/cache_ctrl_logic/n213 [49]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u872  (\biu/cache_ctrl_logic/n214 [50], \biu/cache_ctrl_logic/n211 [50], \biu/cache_ctrl_logic/n213 [50]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u873  (\biu/cache_ctrl_logic/n214 [51], \biu/cache_ctrl_logic/n211 [51], \biu/cache_ctrl_logic/n213 [51]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u874  (\biu/cache_ctrl_logic/n214 [52], \biu/cache_ctrl_logic/n211 [52], \biu/cache_ctrl_logic/n213 [52]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u875  (\biu/cache_ctrl_logic/n214 [53], \biu/cache_ctrl_logic/n211 [53], \biu/cache_ctrl_logic/n213 [53]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u876  (\biu/cache_ctrl_logic/n214 [54], \biu/cache_ctrl_logic/n211 [54], \biu/cache_ctrl_logic/n213 [54]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u877  (\biu/cache_ctrl_logic/n214 [55], \biu/cache_ctrl_logic/n211 [55], \biu/cache_ctrl_logic/n213 [55]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u878  (\biu/cache_ctrl_logic/n214 [56], \biu/cache_ctrl_logic/n211 [56], \biu/cache_ctrl_logic/n213 [56]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u879  (\biu/cache_ctrl_logic/n214 [57], \biu/cache_ctrl_logic/n211 [57], \biu/cache_ctrl_logic/n213 [57]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  and \biu/cache_ctrl_logic/u88  (\biu/cache_ctrl_logic/n64 , \biu/cache_ctrl_logic/n55 , \biu/cache_ctrl_logic/pte_l1i_upd );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(231)
  or \biu/cache_ctrl_logic/u880  (\biu/cache_ctrl_logic/n214 [58], \biu/cache_ctrl_logic/n211 [58], \biu/cache_ctrl_logic/n213 [58]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u881  (\biu/cache_ctrl_logic/n214 [59], \biu/cache_ctrl_logic/n211 [59], \biu/cache_ctrl_logic/n213 [59]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u882  (\biu/cache_ctrl_logic/n214 [60], \biu/cache_ctrl_logic/n211 [60], \biu/cache_ctrl_logic/n213 [60]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u883  (\biu/cache_ctrl_logic/n214 [61], \biu/cache_ctrl_logic/n211 [61], \biu/cache_ctrl_logic/n213 [61]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u884  (\biu/cache_ctrl_logic/n214 [62], \biu/cache_ctrl_logic/n211 [62], \biu/cache_ctrl_logic/n213 [62]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u885  (\biu/cache_ctrl_logic/n214 [63], \biu/cache_ctrl_logic/n211 [63], \biu/cache_ctrl_logic/n213 [63]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(505)
  or \biu/cache_ctrl_logic/u886  (\biu/cache_ctrl_logic/n211 [1], \biu/cache_ctrl_logic/n208 [1], \biu/cache_ctrl_logic/n210 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u887  (\biu/cache_ctrl_logic/n211 [2], \biu/cache_ctrl_logic/n208 [2], \biu/cache_ctrl_logic/n210 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u888  (\biu/cache_ctrl_logic/n211 [3], \biu/cache_ctrl_logic/n208 [3], \biu/cache_ctrl_logic/n210 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u889  (\biu/cache_ctrl_logic/n211 [4], \biu/cache_ctrl_logic/n208 [4], \biu/cache_ctrl_logic/n210 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u89  (\biu/write_data [61], \biu/cache_ctrl_logic/n232 [61], \biu/cache_ctrl_logic/n233 [61]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u890  (\biu/cache_ctrl_logic/n211 [5], \biu/cache_ctrl_logic/n208 [5], \biu/cache_ctrl_logic/n210 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u891  (\biu/cache_ctrl_logic/n211 [6], \biu/cache_ctrl_logic/n208 [6], \biu/cache_ctrl_logic/n210 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u892  (\biu/cache_ctrl_logic/n211 [7], \biu/cache_ctrl_logic/n208 [7], \biu/cache_ctrl_logic/n210 [7]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u893  (\biu/cache_ctrl_logic/n211 [8], \biu/cache_ctrl_logic/n208 [8], \biu/cache_ctrl_logic/n210 [8]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u894  (\biu/cache_ctrl_logic/n211 [9], \biu/cache_ctrl_logic/n208 [9], \biu/cache_ctrl_logic/n210 [9]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u895  (\biu/cache_ctrl_logic/n211 [10], \biu/cache_ctrl_logic/n208 [10], \biu/cache_ctrl_logic/n210 [10]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u896  (\biu/cache_ctrl_logic/n211 [11], \biu/cache_ctrl_logic/n208 [11], \biu/cache_ctrl_logic/n210 [11]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u897  (\biu/cache_ctrl_logic/n211 [12], \biu/cache_ctrl_logic/n208 [12], \biu/cache_ctrl_logic/n210 [12]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u898  (\biu/cache_ctrl_logic/n211 [13], \biu/cache_ctrl_logic/n208 [13], \biu/cache_ctrl_logic/n210 [13]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u899  (\biu/cache_ctrl_logic/n211 [14], \biu/cache_ctrl_logic/n208 [14], \biu/cache_ctrl_logic/n210 [14]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  and \biu/cache_ctrl_logic/u9  (\biu/cache_ctrl_logic/pte_l1d_upd , \biu/cache_ctrl_logic/l1d_write_through , \biu/cache_ctrl_logic/n1 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(181)
  and \biu/cache_ctrl_logic/u90  (\biu/cache_ctrl_logic/n65 , \biu/cache_ctrl_logic/n55 , \biu/cache_ctrl_logic/l1d_write_through );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(235)
  or \biu/cache_ctrl_logic/u900  (\biu/cache_ctrl_logic/n211 [15], \biu/cache_ctrl_logic/n208 [15], \biu/cache_ctrl_logic/n210 [15]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u901  (\biu/cache_ctrl_logic/n211 [16], \biu/cache_ctrl_logic/n208 [16], \biu/cache_ctrl_logic/n210 [16]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u902  (\biu/cache_ctrl_logic/n211 [17], \biu/cache_ctrl_logic/n208 [17], \biu/cache_ctrl_logic/n210 [17]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u903  (\biu/cache_ctrl_logic/n211 [18], \biu/cache_ctrl_logic/n208 [18], \biu/cache_ctrl_logic/n210 [18]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u904  (\biu/cache_ctrl_logic/n211 [19], \biu/cache_ctrl_logic/n208 [19], \biu/cache_ctrl_logic/n210 [19]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u905  (\biu/cache_ctrl_logic/n211 [20], \biu/cache_ctrl_logic/n208 [20], \biu/cache_ctrl_logic/n210 [20]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u906  (\biu/cache_ctrl_logic/n211 [21], \biu/cache_ctrl_logic/n208 [21], \biu/cache_ctrl_logic/n210 [21]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u907  (\biu/cache_ctrl_logic/n211 [22], \biu/cache_ctrl_logic/n208 [22], \biu/cache_ctrl_logic/n210 [22]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u908  (\biu/cache_ctrl_logic/n211 [23], \biu/cache_ctrl_logic/n208 [23], \biu/cache_ctrl_logic/n210 [23]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u909  (\biu/cache_ctrl_logic/n211 [24], \biu/cache_ctrl_logic/n208 [24], \biu/cache_ctrl_logic/n210 [24]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u91  (\biu/write_data [60], \biu/cache_ctrl_logic/n232 [60], \biu/cache_ctrl_logic/n233 [60]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u910  (\biu/cache_ctrl_logic/n211 [25], \biu/cache_ctrl_logic/n208 [25], \biu/cache_ctrl_logic/n210 [25]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u911  (\biu/cache_ctrl_logic/n211 [26], \biu/cache_ctrl_logic/n208 [26], \biu/cache_ctrl_logic/n210 [26]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u912  (\biu/cache_ctrl_logic/n211 [27], \biu/cache_ctrl_logic/n208 [27], \biu/cache_ctrl_logic/n210 [27]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u913  (\biu/cache_ctrl_logic/n211 [28], \biu/cache_ctrl_logic/n208 [28], \biu/cache_ctrl_logic/n210 [28]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u914  (\biu/cache_ctrl_logic/n211 [29], \biu/cache_ctrl_logic/n208 [29], \biu/cache_ctrl_logic/n210 [29]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u915  (\biu/cache_ctrl_logic/n211 [30], \biu/cache_ctrl_logic/n208 [30], \biu/cache_ctrl_logic/n210 [30]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u916  (\biu/cache_ctrl_logic/n211 [31], \biu/cache_ctrl_logic/n208 [31], \biu/cache_ctrl_logic/n210 [31]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u917  (\biu/cache_ctrl_logic/n211 [32], \biu/cache_ctrl_logic/n208 [32], \biu/cache_ctrl_logic/n210 [32]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u918  (\biu/cache_ctrl_logic/n211 [33], \biu/cache_ctrl_logic/n208 [33], \biu/cache_ctrl_logic/n210 [33]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u919  (\biu/cache_ctrl_logic/n211 [34], \biu/cache_ctrl_logic/n208 [34], \biu/cache_ctrl_logic/n210 [34]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  and \biu/cache_ctrl_logic/u92  (\biu/cache_ctrl_logic/n66 , \biu/cache_ctrl_logic/n55 , \biu/cache_ctrl_logic/l1i_write_through );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(238)
  or \biu/cache_ctrl_logic/u920  (\biu/cache_ctrl_logic/n211 [35], \biu/cache_ctrl_logic/n208 [35], \biu/cache_ctrl_logic/n210 [35]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u921  (\biu/cache_ctrl_logic/n211 [36], \biu/cache_ctrl_logic/n208 [36], \biu/cache_ctrl_logic/n210 [36]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u922  (\biu/cache_ctrl_logic/n211 [37], \biu/cache_ctrl_logic/n208 [37], \biu/cache_ctrl_logic/n210 [37]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u923  (\biu/cache_ctrl_logic/n211 [38], \biu/cache_ctrl_logic/n208 [38], \biu/cache_ctrl_logic/n210 [38]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u924  (\biu/cache_ctrl_logic/n211 [39], \biu/cache_ctrl_logic/n208 [39], \biu/cache_ctrl_logic/n210 [39]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u925  (\biu/cache_ctrl_logic/n211 [40], \biu/cache_ctrl_logic/n208 [40], \biu/cache_ctrl_logic/n210 [40]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u926  (\biu/cache_ctrl_logic/n211 [41], \biu/cache_ctrl_logic/n208 [41], \biu/cache_ctrl_logic/n210 [41]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u927  (\biu/cache_ctrl_logic/n211 [42], \biu/cache_ctrl_logic/n208 [42], \biu/cache_ctrl_logic/n210 [42]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u928  (\biu/cache_ctrl_logic/n211 [43], \biu/cache_ctrl_logic/n208 [43], \biu/cache_ctrl_logic/n210 [43]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u929  (\biu/cache_ctrl_logic/n211 [44], \biu/cache_ctrl_logic/n208 [44], \biu/cache_ctrl_logic/n210 [44]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  and \biu/cache_ctrl_logic/u93  (\biu/cache_ctrl_logic/n68 , \biu/trans_rdy , \biu/cacheable );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(250)
  or \biu/cache_ctrl_logic/u930  (\biu/cache_ctrl_logic/n211 [45], \biu/cache_ctrl_logic/n208 [45], \biu/cache_ctrl_logic/n210 [45]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u931  (\biu/cache_ctrl_logic/n211 [46], \biu/cache_ctrl_logic/n208 [46], \biu/cache_ctrl_logic/n210 [46]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u932  (\biu/cache_ctrl_logic/n211 [47], \biu/cache_ctrl_logic/n208 [47], \biu/cache_ctrl_logic/n210 [47]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u933  (\biu/cache_ctrl_logic/n211 [48], \biu/cache_ctrl_logic/n208 [48], \biu/cache_ctrl_logic/n210 [48]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u934  (\biu/cache_ctrl_logic/n211 [49], \biu/cache_ctrl_logic/n208 [49], \biu/cache_ctrl_logic/n210 [49]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u935  (\biu/cache_ctrl_logic/n211 [50], \biu/cache_ctrl_logic/n208 [50], \biu/cache_ctrl_logic/n210 [50]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u936  (\biu/cache_ctrl_logic/n211 [51], \biu/cache_ctrl_logic/n208 [51], \biu/cache_ctrl_logic/n210 [51]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u937  (\biu/cache_ctrl_logic/n211 [52], \biu/cache_ctrl_logic/n208 [52], \biu/cache_ctrl_logic/n210 [52]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u938  (\biu/cache_ctrl_logic/n211 [53], \biu/cache_ctrl_logic/n208 [53], \biu/cache_ctrl_logic/n210 [53]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u939  (\biu/cache_ctrl_logic/n211 [54], \biu/cache_ctrl_logic/n208 [54], \biu/cache_ctrl_logic/n210 [54]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u94  (\biu/cache_ctrl_logic/n69 , \biu/trans_rdy , \biu/bus_error );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(250)
  or \biu/cache_ctrl_logic/u940  (\biu/cache_ctrl_logic/n211 [55], \biu/cache_ctrl_logic/n208 [55], \biu/cache_ctrl_logic/n210 [55]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u941  (\biu/cache_ctrl_logic/n211 [56], \biu/cache_ctrl_logic/n208 [56], \biu/cache_ctrl_logic/n210 [56]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u942  (\biu/cache_ctrl_logic/n211 [57], \biu/cache_ctrl_logic/n208 [57], \biu/cache_ctrl_logic/n210 [57]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u943  (\biu/cache_ctrl_logic/n211 [58], \biu/cache_ctrl_logic/n208 [58], \biu/cache_ctrl_logic/n210 [58]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u944  (\biu/cache_ctrl_logic/n211 [59], \biu/cache_ctrl_logic/n208 [59], \biu/cache_ctrl_logic/n210 [59]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u945  (\biu/cache_ctrl_logic/n211 [60], \biu/cache_ctrl_logic/n208 [60], \biu/cache_ctrl_logic/n210 [60]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u946  (\biu/cache_ctrl_logic/n211 [61], \biu/cache_ctrl_logic/n208 [61], \biu/cache_ctrl_logic/n210 [61]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u947  (\biu/cache_ctrl_logic/n211 [62], \biu/cache_ctrl_logic/n208 [62], \biu/cache_ctrl_logic/n210 [62]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u948  (\biu/cache_ctrl_logic/n211 [63], \biu/cache_ctrl_logic/n208 [63], \biu/cache_ctrl_logic/n210 [63]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(504)
  or \biu/cache_ctrl_logic/u949  (\biu/cache_ctrl_logic/n186 [1], \biu/cache_ctrl_logic/n190 [0], \biu/cache_ctrl_logic/n185 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(472)
  not \biu/cache_ctrl_logic/u95  (\biu/cache_ctrl_logic/n73 [2], \biu/trans_rdy );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(254)
  or \biu/cache_ctrl_logic/u950  (\biu/cache_ctrl_logic/n186 [2], \biu/cache_ctrl_logic/n190 [1], \biu/cache_ctrl_logic/n185 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(472)
  or \biu/cache_ctrl_logic/u951  (\biu/cache_ctrl_logic/n186 [3], \biu/cache_ctrl_logic/n190 [2], \biu/cache_ctrl_logic/n185 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(472)
  or \biu/cache_ctrl_logic/u952  (\biu/cache_ctrl_logic/n186 [4], \biu/cache_ctrl_logic/n190 [3], \biu/cache_ctrl_logic/n185 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(472)
  or \biu/cache_ctrl_logic/u953  (\biu/cache_ctrl_logic/n186 [5], \biu/cache_ctrl_logic/n190 [4], \biu/cache_ctrl_logic/n185 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(472)
  or \biu/cache_ctrl_logic/u954  (\biu/cache_ctrl_logic/n190 [1], \biu/cache_ctrl_logic/n193 [0], \biu/cache_ctrl_logic/n189 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(471)
  or \biu/cache_ctrl_logic/u955  (\biu/cache_ctrl_logic/n190 [2], \biu/cache_ctrl_logic/n193 [1], \biu/cache_ctrl_logic/n189 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(471)
  or \biu/cache_ctrl_logic/u956  (\biu/cache_ctrl_logic/n190 [3], \biu/cache_ctrl_logic/n193 [2], \biu/cache_ctrl_logic/n189 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(471)
  or \biu/cache_ctrl_logic/u957  (\biu/cache_ctrl_logic/n190 [4], \biu/cache_ctrl_logic/n189 [6], \biu/cache_ctrl_logic/n189 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(471)
  or \biu/cache_ctrl_logic/u958  (\biu/cache_ctrl_logic/n193 [1], \biu/cache_ctrl_logic/n189 [6], \biu/cache_ctrl_logic/n189 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(466)
  or \biu/cache_ctrl_logic/u959  (\biu/cache_ctrl_logic/n193 [2], \biu/cache_ctrl_logic/n189 [6], \biu/cache_ctrl_logic/n189 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(466)
  not \biu/cache_ctrl_logic/u96  (\biu/cache_ctrl_logic/n80 [2], \biu/cache_ctrl_logic/n79 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  and \biu/cache_ctrl_logic/u960  (\biu/cache_ctrl_logic/n189 [1], \biu/cache_ctrl_logic/n187 , \biu/cache_ctrl_logic/n176 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(470)
  and \biu/cache_ctrl_logic/u961  (\biu/cache_ctrl_logic/n189 [2], \biu/cache_ctrl_logic/n191 , \biu/cache_ctrl_logic/n176 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(470)
  and \biu/cache_ctrl_logic/u962  (\biu/cache_ctrl_logic/n189 [4], \biu/cache_ctrl_logic/n194 , \biu/cache_ctrl_logic/n176 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(470)
  and \biu/cache_ctrl_logic/u963  (\biu/cache_ctrl_logic/n189 [5], \biu/cache_ctrl_logic/n172 , \biu/cache_ctrl_logic/n188 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(470)
  and \biu/cache_ctrl_logic/u964  (\biu/cache_ctrl_logic/n189 [6], \biu/cache_ctrl_logic/n172 , \biu/cache_ctrl_logic/n178 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(470)
  and \biu/cache_ctrl_logic/u965  (\biu/cache_ctrl_logic/n185 [1], \biu/cache_ctrl_logic/n187 , \biu/cache_ctrl_logic/n184 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(448)
  and \biu/cache_ctrl_logic/u966  (\biu/cache_ctrl_logic/n185 [2], \biu/cache_ctrl_logic/n191 , \biu/cache_ctrl_logic/n184 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(448)
  and \biu/cache_ctrl_logic/u967  (\biu/cache_ctrl_logic/n185 [3], \biu/cache_ctrl_logic/n194 , \biu/cache_ctrl_logic/n184 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(448)
  and \biu/cache_ctrl_logic/u968  (\biu/cache_ctrl_logic/n185 [4], \biu/cache_ctrl_logic/n195 , \biu/cache_ctrl_logic/n174 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(448)
  and \biu/cache_ctrl_logic/u969  (\biu/cache_ctrl_logic/n185 [5], \biu/cache_ctrl_logic/n196 , \biu/cache_ctrl_logic/n174 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(448)
  and \biu/cache_ctrl_logic/u97  (\biu/cache_ctrl_logic/n76 , \biu/page_fault , write);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  and \biu/cache_ctrl_logic/u974  (\biu/cache_ctrl_logic/n182 [1], \biu/cache_ctrl_logic/n187 , \biu/cache_ctrl_logic/n177 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(446)
  and \biu/cache_ctrl_logic/u975  (\biu/cache_ctrl_logic/n182 [2], \biu/cache_ctrl_logic/n191 , \biu/cache_ctrl_logic/n177 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(446)
  and \biu/cache_ctrl_logic/u976  (\biu/cache_ctrl_logic/n182 [3], \biu/cache_ctrl_logic/n194 , \biu/cache_ctrl_logic/n177 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(446)
  and \biu/cache_ctrl_logic/u977  (\biu/cache_ctrl_logic/n182 [4], \biu/cache_ctrl_logic/n195 , \biu/cache_ctrl_logic/n175 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(446)
  and \biu/cache_ctrl_logic/u978  (\biu/cache_ctrl_logic/n182 [5], \biu/cache_ctrl_logic/n196 , \biu/cache_ctrl_logic/n175 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(446)
  and \biu/cache_ctrl_logic/u979  (\biu/cache_ctrl_logic/n182 [6], \biu/cache_ctrl_logic/n197 , \biu/cache_ctrl_logic/n173 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(446)
  and \biu/cache_ctrl_logic/u98  (\biu/cache_ctrl_logic/n77 , \biu/page_fault , read);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(259)
  and \biu/cache_ctrl_logic/u980  (\biu/cache_ctrl_logic/n182 [7], \biu/cache_ctrl_logic/n172 , \biu/cache_ctrl_logic/n181 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(446)
  or \biu/cache_ctrl_logic/u983  (\biu/cache_ctrl_logic/n181 [6], \biu/cache_ctrl_logic/n184 [3], \biu/cache_ctrl_logic/n178 );  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(446)
  or \biu/cache_ctrl_logic/u985  (\biu/cache_ctrl_logic/ex_bsel [2], \biu/cache_ctrl_logic/n186 [0], \biu/cache_ctrl_logic/n182 [1]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(473)
  or \biu/cache_ctrl_logic/u986  (\biu/cache_ctrl_logic/ex_bsel [3], \biu/cache_ctrl_logic/n186 [1], \biu/cache_ctrl_logic/n182 [2]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(473)
  or \biu/cache_ctrl_logic/u987  (\biu/cache_ctrl_logic/ex_bsel [4], \biu/cache_ctrl_logic/n186 [2], \biu/cache_ctrl_logic/n182 [3]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(473)
  or \biu/cache_ctrl_logic/u988  (\biu/cache_ctrl_logic/ex_bsel [5], \biu/cache_ctrl_logic/n186 [3], \biu/cache_ctrl_logic/n182 [4]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(473)
  or \biu/cache_ctrl_logic/u989  (\biu/cache_ctrl_logic/ex_bsel [6], \biu/cache_ctrl_logic/n186 [4], \biu/cache_ctrl_logic/n182 [5]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(473)
  or \biu/cache_ctrl_logic/u99  (\biu/write_data [59], \biu/cache_ctrl_logic/n232 [59], \biu/cache_ctrl_logic/n233 [59]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(520)
  or \biu/cache_ctrl_logic/u990  (\biu/cache_ctrl_logic/ex_bsel [7], \biu/cache_ctrl_logic/n186 [5], \biu/cache_ctrl_logic/n182 [6]);  // ../../RTL/CPU/BIU/cache_ctrl_logic.v(473)
  not \biu/ex_data_sel[1]_inv  (\biu/ex_data_sel[1]_neg , \biu/ex_data_sel [1]);
  binary_mux_s1_w1 \biu/mux0_b0  (
    .i0(addr_if[3]),
    .i1(addr_ex[3]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n0 [0]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux0_b1  (
    .i0(addr_if[4]),
    .i1(addr_ex[4]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n0 [1]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux0_b2  (
    .i0(addr_if[5]),
    .i1(addr_ex[5]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n0 [2]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux0_b3  (
    .i0(addr_if[6]),
    .i1(addr_ex[6]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n0 [3]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux0_b4  (
    .i0(addr_if[7]),
    .i1(addr_ex[7]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n0 [4]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux0_b5  (
    .i0(addr_if[8]),
    .i1(addr_ex[8]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n0 [5]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux0_b6  (
    .i0(addr_if[9]),
    .i1(addr_ex[9]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n0 [6]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux0_b7  (
    .i0(addr_if[10]),
    .i1(addr_ex[10]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n0 [7]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux0_b8  (
    .i0(addr_if[11]),
    .i1(addr_ex[11]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n0 [8]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux1_b0  (
    .i0(\biu/n0 [0]),
    .i1(\biu/cache_counter [0]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_addr [0]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux1_b1  (
    .i0(\biu/n0 [1]),
    .i1(\biu/cache_counter [1]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_addr [1]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux1_b2  (
    .i0(\biu/n0 [2]),
    .i1(\biu/cache_counter [2]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_addr [2]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux1_b3  (
    .i0(\biu/n0 [3]),
    .i1(\biu/cache_counter [3]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_addr [3]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux1_b4  (
    .i0(\biu/n0 [4]),
    .i1(\biu/cache_counter [4]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_addr [4]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux1_b5  (
    .i0(\biu/n0 [5]),
    .i1(\biu/cache_counter [5]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_addr [5]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux1_b6  (
    .i0(\biu/n0 [6]),
    .i1(\biu/cache_counter [6]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_addr [6]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux1_b7  (
    .i0(\biu/n0 [7]),
    .i1(\biu/cache_counter [7]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_addr [7]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux1_b8  (
    .i0(\biu/n0 [8]),
    .i1(\biu/cache_counter [8]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_addr [8]));  // ../../RTL/CPU/BIU/biu.v(131)
  binary_mux_s1_w1 \biu/mux2_b0  (
    .i0(addr_ex[0]),
    .i1(\biu/cache_counter [0]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1d_addr [0]));  // ../../RTL/CPU/BIU/biu.v(133)
  binary_mux_s1_w1 \biu/mux2_b1  (
    .i0(addr_ex[1]),
    .i1(\biu/cache_counter [1]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1d_addr [1]));  // ../../RTL/CPU/BIU/biu.v(133)
  binary_mux_s1_w1 \biu/mux2_b2  (
    .i0(addr_ex[2]),
    .i1(\biu/cache_counter [2]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1d_addr [2]));  // ../../RTL/CPU/BIU/biu.v(133)
  binary_mux_s1_w1 \biu/mux2_b3  (
    .i0(addr_ex[3]),
    .i1(\biu/cache_counter [3]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1d_addr [3]));  // ../../RTL/CPU/BIU/biu.v(133)
  binary_mux_s1_w1 \biu/mux2_b4  (
    .i0(addr_ex[4]),
    .i1(\biu/cache_counter [4]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1d_addr [4]));  // ../../RTL/CPU/BIU/biu.v(133)
  binary_mux_s1_w1 \biu/mux2_b5  (
    .i0(addr_ex[5]),
    .i1(\biu/cache_counter [5]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1d_addr [5]));  // ../../RTL/CPU/BIU/biu.v(133)
  binary_mux_s1_w1 \biu/mux2_b6  (
    .i0(addr_ex[6]),
    .i1(\biu/cache_counter [6]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1d_addr [6]));  // ../../RTL/CPU/BIU/biu.v(133)
  binary_mux_s1_w1 \biu/mux2_b7  (
    .i0(addr_ex[7]),
    .i1(\biu/cache_counter [7]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1d_addr [7]));  // ../../RTL/CPU/BIU/biu.v(133)
  binary_mux_s1_w1 \biu/mux2_b8  (
    .i0(addr_ex[8]),
    .i1(\biu/cache_counter [8]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1d_addr [8]));  // ../../RTL/CPU/BIU/biu.v(133)
  binary_mux_s1_w1 \biu/mux3_b0  (
    .i0(\exu/lsu/n1 [0]),
    .i1(uncache_data[0]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [0]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b1  (
    .i0(\exu/lsu/n1 [1]),
    .i1(uncache_data[1]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [1]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b10  (
    .i0(\exu/lsu/n4 [10]),
    .i1(uncache_data[10]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [10]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b11  (
    .i0(\exu/lsu/n4 [11]),
    .i1(uncache_data[11]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [11]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b12  (
    .i0(\exu/lsu/n4 [12]),
    .i1(uncache_data[12]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [12]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b13  (
    .i0(\exu/lsu/n4 [13]),
    .i1(uncache_data[13]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [13]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b14  (
    .i0(\exu/lsu/n4 [14]),
    .i1(uncache_data[14]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [14]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b15  (
    .i0(\exu/lsu/n4 [15]),
    .i1(uncache_data[15]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [15]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b16  (
    .i0(\exu/lsu/n7 [16]),
    .i1(uncache_data[16]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [16]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b17  (
    .i0(\exu/lsu/n7 [17]),
    .i1(uncache_data[17]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [17]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b18  (
    .i0(\exu/lsu/n7 [18]),
    .i1(uncache_data[18]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [18]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b19  (
    .i0(\exu/lsu/n7 [19]),
    .i1(uncache_data[19]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [19]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b2  (
    .i0(\exu/lsu/n1 [2]),
    .i1(uncache_data[2]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [2]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b20  (
    .i0(\exu/lsu/n7 [20]),
    .i1(uncache_data[20]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [20]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b21  (
    .i0(\exu/lsu/n7 [21]),
    .i1(uncache_data[21]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [21]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b22  (
    .i0(\exu/lsu/n7 [22]),
    .i1(uncache_data[22]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [22]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b23  (
    .i0(\exu/lsu/n7 [23]),
    .i1(uncache_data[23]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [23]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b24  (
    .i0(\exu/lsu/n10 [24]),
    .i1(uncache_data[24]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [24]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b25  (
    .i0(\exu/lsu/n10 [25]),
    .i1(uncache_data[25]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [25]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b26  (
    .i0(\exu/lsu/n10 [26]),
    .i1(uncache_data[26]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [26]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b27  (
    .i0(\exu/lsu/n10 [27]),
    .i1(uncache_data[27]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [27]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b28  (
    .i0(\exu/lsu/n10 [28]),
    .i1(uncache_data[28]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [28]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b29  (
    .i0(\exu/lsu/n10 [29]),
    .i1(uncache_data[29]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [29]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b3  (
    .i0(\exu/lsu/n1 [3]),
    .i1(uncache_data[3]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [3]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b30  (
    .i0(\exu/lsu/n10 [30]),
    .i1(uncache_data[30]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [30]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b31  (
    .i0(\exu/lsu/n10 [31]),
    .i1(uncache_data[31]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [31]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b32  (
    .i0(\exu/lsu/n10 [32]),
    .i1(uncache_data[32]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [32]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b33  (
    .i0(\exu/lsu/n10 [33]),
    .i1(uncache_data[33]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [33]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b34  (
    .i0(\exu/lsu/n10 [34]),
    .i1(uncache_data[34]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [34]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b35  (
    .i0(\exu/lsu/n10 [35]),
    .i1(uncache_data[35]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [35]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b36  (
    .i0(\exu/lsu/n10 [36]),
    .i1(uncache_data[36]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [36]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b37  (
    .i0(\exu/lsu/n10 [37]),
    .i1(uncache_data[37]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [37]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b38  (
    .i0(\exu/lsu/n10 [38]),
    .i1(uncache_data[38]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [38]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b39  (
    .i0(\exu/lsu/n10 [39]),
    .i1(uncache_data[39]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [39]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b4  (
    .i0(\exu/lsu/n1 [4]),
    .i1(uncache_data[4]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [4]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b40  (
    .i0(\exu/lsu/n10 [40]),
    .i1(uncache_data[40]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [40]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b41  (
    .i0(\exu/lsu/n10 [41]),
    .i1(uncache_data[41]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [41]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b42  (
    .i0(\exu/lsu/n10 [42]),
    .i1(uncache_data[42]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [42]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b43  (
    .i0(\exu/lsu/n10 [43]),
    .i1(uncache_data[43]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [43]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b44  (
    .i0(\exu/lsu/n10 [44]),
    .i1(uncache_data[44]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [44]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b45  (
    .i0(\exu/lsu/n10 [45]),
    .i1(uncache_data[45]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [45]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b46  (
    .i0(\exu/lsu/n10 [46]),
    .i1(uncache_data[46]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [46]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b47  (
    .i0(\exu/lsu/n10 [47]),
    .i1(uncache_data[47]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [47]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b48  (
    .i0(\exu/lsu/n10 [48]),
    .i1(uncache_data[48]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [48]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b49  (
    .i0(\exu/lsu/n10 [49]),
    .i1(uncache_data[49]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [49]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b5  (
    .i0(\exu/lsu/n1 [5]),
    .i1(uncache_data[5]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [5]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b50  (
    .i0(\exu/lsu/n10 [50]),
    .i1(uncache_data[50]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [50]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b51  (
    .i0(\exu/lsu/n10 [51]),
    .i1(uncache_data[51]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [51]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b52  (
    .i0(\exu/lsu/n10 [52]),
    .i1(uncache_data[52]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [52]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b53  (
    .i0(\exu/lsu/n10 [53]),
    .i1(uncache_data[53]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [53]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b54  (
    .i0(\exu/lsu/n10 [54]),
    .i1(uncache_data[54]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [54]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b55  (
    .i0(\exu/lsu/n10 [55]),
    .i1(uncache_data[55]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [55]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b56  (
    .i0(\exu/lsu/n10 [56]),
    .i1(uncache_data[56]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [56]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b57  (
    .i0(\exu/lsu/n10 [57]),
    .i1(uncache_data[57]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [57]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b58  (
    .i0(\exu/lsu/n10 [58]),
    .i1(uncache_data[58]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [58]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b59  (
    .i0(\exu/lsu/n10 [59]),
    .i1(uncache_data[59]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [59]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b6  (
    .i0(\exu/lsu/n1 [6]),
    .i1(uncache_data[6]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [6]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b60  (
    .i0(\exu/lsu/n10 [60]),
    .i1(uncache_data[60]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [60]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b61  (
    .i0(\exu/lsu/n10 [61]),
    .i1(uncache_data[61]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [61]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b62  (
    .i0(\exu/lsu/n10 [62]),
    .i1(uncache_data[62]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [62]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b63  (
    .i0(\exu/lsu/n10 [63]),
    .i1(uncache_data[63]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [63]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b7  (
    .i0(\exu/lsu/n1 [7]),
    .i1(uncache_data[7]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [7]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b8  (
    .i0(\exu/lsu/n4 [8]),
    .i1(uncache_data[8]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [8]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux3_b9  (
    .i0(\exu/lsu/n4 [9]),
    .i1(uncache_data[9]),
    .sel(\biu/cache_addr_sel ),
    .o(\biu/l1i_in [9]));  // ../../RTL/CPU/BIU/biu.v(135)
  binary_mux_s1_w1 \biu/mux4_b0  (
    .i0(\biu/l1d_out [0]),
    .i1(ins_read[0]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [0]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b1  (
    .i0(\biu/l1d_out [1]),
    .i1(ins_read[1]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [1]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b10  (
    .i0(\biu/l1d_out [10]),
    .i1(ins_read[10]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [10]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b11  (
    .i0(\biu/l1d_out [11]),
    .i1(ins_read[11]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [11]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b12  (
    .i0(\biu/l1d_out [12]),
    .i1(ins_read[12]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [12]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b13  (
    .i0(\biu/l1d_out [13]),
    .i1(ins_read[13]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [13]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b14  (
    .i0(\biu/l1d_out [14]),
    .i1(ins_read[14]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [14]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b15  (
    .i0(\biu/l1d_out [15]),
    .i1(ins_read[15]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [15]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b16  (
    .i0(\biu/l1d_out [16]),
    .i1(ins_read[16]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [16]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b17  (
    .i0(\biu/l1d_out [17]),
    .i1(ins_read[17]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [17]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b18  (
    .i0(\biu/l1d_out [18]),
    .i1(ins_read[18]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [18]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b19  (
    .i0(\biu/l1d_out [19]),
    .i1(ins_read[19]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [19]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b2  (
    .i0(\biu/l1d_out [2]),
    .i1(ins_read[2]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [2]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b20  (
    .i0(\biu/l1d_out [20]),
    .i1(ins_read[20]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [20]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b21  (
    .i0(\biu/l1d_out [21]),
    .i1(ins_read[21]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [21]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b22  (
    .i0(\biu/l1d_out [22]),
    .i1(ins_read[22]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [22]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b23  (
    .i0(\biu/l1d_out [23]),
    .i1(ins_read[23]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [23]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b24  (
    .i0(\biu/l1d_out [24]),
    .i1(ins_read[24]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [24]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b25  (
    .i0(\biu/l1d_out [25]),
    .i1(ins_read[25]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [25]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b26  (
    .i0(\biu/l1d_out [26]),
    .i1(ins_read[26]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [26]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b27  (
    .i0(\biu/l1d_out [27]),
    .i1(ins_read[27]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [27]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b28  (
    .i0(\biu/l1d_out [28]),
    .i1(ins_read[28]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [28]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b29  (
    .i0(\biu/l1d_out [29]),
    .i1(ins_read[29]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [29]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b3  (
    .i0(\biu/l1d_out [3]),
    .i1(ins_read[3]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [3]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b30  (
    .i0(\biu/l1d_out [30]),
    .i1(ins_read[30]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [30]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b31  (
    .i0(\biu/l1d_out [31]),
    .i1(ins_read[31]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [31]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b32  (
    .i0(\biu/l1d_out [32]),
    .i1(ins_read[32]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [32]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b33  (
    .i0(\biu/l1d_out [33]),
    .i1(ins_read[33]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [33]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b34  (
    .i0(\biu/l1d_out [34]),
    .i1(ins_read[34]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [34]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b35  (
    .i0(\biu/l1d_out [35]),
    .i1(ins_read[35]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [35]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b36  (
    .i0(\biu/l1d_out [36]),
    .i1(ins_read[36]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [36]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b37  (
    .i0(\biu/l1d_out [37]),
    .i1(ins_read[37]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [37]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b38  (
    .i0(\biu/l1d_out [38]),
    .i1(ins_read[38]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [38]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b39  (
    .i0(\biu/l1d_out [39]),
    .i1(ins_read[39]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [39]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b4  (
    .i0(\biu/l1d_out [4]),
    .i1(ins_read[4]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [4]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b40  (
    .i0(\biu/l1d_out [40]),
    .i1(ins_read[40]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [40]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b41  (
    .i0(\biu/l1d_out [41]),
    .i1(ins_read[41]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [41]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b42  (
    .i0(\biu/l1d_out [42]),
    .i1(ins_read[42]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [42]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b43  (
    .i0(\biu/l1d_out [43]),
    .i1(ins_read[43]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [43]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b44  (
    .i0(\biu/l1d_out [44]),
    .i1(ins_read[44]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [44]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b45  (
    .i0(\biu/l1d_out [45]),
    .i1(ins_read[45]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [45]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b46  (
    .i0(\biu/l1d_out [46]),
    .i1(ins_read[46]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [46]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b47  (
    .i0(\biu/l1d_out [47]),
    .i1(ins_read[47]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [47]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b48  (
    .i0(\biu/l1d_out [48]),
    .i1(ins_read[48]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [48]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b49  (
    .i0(\biu/l1d_out [49]),
    .i1(ins_read[49]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [49]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b5  (
    .i0(\biu/l1d_out [5]),
    .i1(ins_read[5]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [5]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b50  (
    .i0(\biu/l1d_out [50]),
    .i1(ins_read[50]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [50]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b51  (
    .i0(\biu/l1d_out [51]),
    .i1(ins_read[51]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [51]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b52  (
    .i0(\biu/l1d_out [52]),
    .i1(ins_read[52]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [52]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b53  (
    .i0(\biu/l1d_out [53]),
    .i1(ins_read[53]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [53]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b54  (
    .i0(\biu/l1d_out [54]),
    .i1(ins_read[54]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [54]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b55  (
    .i0(\biu/l1d_out [55]),
    .i1(ins_read[55]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [55]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b56  (
    .i0(\biu/l1d_out [56]),
    .i1(ins_read[56]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [56]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b57  (
    .i0(\biu/l1d_out [57]),
    .i1(ins_read[57]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [57]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b58  (
    .i0(\biu/l1d_out [58]),
    .i1(ins_read[58]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [58]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b59  (
    .i0(\biu/l1d_out [59]),
    .i1(ins_read[59]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [59]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b6  (
    .i0(\biu/l1d_out [6]),
    .i1(ins_read[6]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [6]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b60  (
    .i0(\biu/l1d_out [60]),
    .i1(ins_read[60]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [60]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b61  (
    .i0(\biu/l1d_out [61]),
    .i1(ins_read[61]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [61]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b62  (
    .i0(\biu/l1d_out [62]),
    .i1(ins_read[62]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [62]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b63  (
    .i0(\biu/l1d_out [63]),
    .i1(ins_read[63]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [63]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b7  (
    .i0(\biu/l1d_out [7]),
    .i1(ins_read[7]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [7]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b8  (
    .i0(\biu/l1d_out [8]),
    .i1(ins_read[8]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [8]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux4_b9  (
    .i0(\biu/l1d_out [9]),
    .i1(ins_read[9]),
    .sel(\biu/ex_data_sel [0]),
    .o(\biu/n1 [9]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b0  (
    .i0(\biu/n1 [0]),
    .i1(uncache_data[0]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[0]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b1  (
    .i0(\biu/n1 [1]),
    .i1(uncache_data[1]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[1]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b10  (
    .i0(\biu/n1 [10]),
    .i1(uncache_data[10]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[10]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b11  (
    .i0(\biu/n1 [11]),
    .i1(uncache_data[11]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[11]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b12  (
    .i0(\biu/n1 [12]),
    .i1(uncache_data[12]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[12]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b13  (
    .i0(\biu/n1 [13]),
    .i1(uncache_data[13]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[13]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b14  (
    .i0(\biu/n1 [14]),
    .i1(uncache_data[14]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[14]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b15  (
    .i0(\biu/n1 [15]),
    .i1(uncache_data[15]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[15]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b16  (
    .i0(\biu/n1 [16]),
    .i1(uncache_data[16]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[16]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b17  (
    .i0(\biu/n1 [17]),
    .i1(uncache_data[17]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[17]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b18  (
    .i0(\biu/n1 [18]),
    .i1(uncache_data[18]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[18]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b19  (
    .i0(\biu/n1 [19]),
    .i1(uncache_data[19]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[19]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b2  (
    .i0(\biu/n1 [2]),
    .i1(uncache_data[2]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[2]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b20  (
    .i0(\biu/n1 [20]),
    .i1(uncache_data[20]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[20]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b21  (
    .i0(\biu/n1 [21]),
    .i1(uncache_data[21]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[21]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b22  (
    .i0(\biu/n1 [22]),
    .i1(uncache_data[22]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[22]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b23  (
    .i0(\biu/n1 [23]),
    .i1(uncache_data[23]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[23]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b24  (
    .i0(\biu/n1 [24]),
    .i1(uncache_data[24]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[24]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b25  (
    .i0(\biu/n1 [25]),
    .i1(uncache_data[25]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[25]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b26  (
    .i0(\biu/n1 [26]),
    .i1(uncache_data[26]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[26]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b27  (
    .i0(\biu/n1 [27]),
    .i1(uncache_data[27]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[27]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b28  (
    .i0(\biu/n1 [28]),
    .i1(uncache_data[28]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[28]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b29  (
    .i0(\biu/n1 [29]),
    .i1(uncache_data[29]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[29]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b3  (
    .i0(\biu/n1 [3]),
    .i1(uncache_data[3]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[3]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b30  (
    .i0(\biu/n1 [30]),
    .i1(uncache_data[30]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[30]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b31  (
    .i0(\biu/n1 [31]),
    .i1(uncache_data[31]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[31]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b32  (
    .i0(\biu/n1 [32]),
    .i1(uncache_data[32]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[32]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b33  (
    .i0(\biu/n1 [33]),
    .i1(uncache_data[33]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[33]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b34  (
    .i0(\biu/n1 [34]),
    .i1(uncache_data[34]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[34]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b35  (
    .i0(\biu/n1 [35]),
    .i1(uncache_data[35]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[35]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b36  (
    .i0(\biu/n1 [36]),
    .i1(uncache_data[36]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[36]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b37  (
    .i0(\biu/n1 [37]),
    .i1(uncache_data[37]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[37]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b38  (
    .i0(\biu/n1 [38]),
    .i1(uncache_data[38]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[38]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b39  (
    .i0(\biu/n1 [39]),
    .i1(uncache_data[39]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[39]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b4  (
    .i0(\biu/n1 [4]),
    .i1(uncache_data[4]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[4]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b40  (
    .i0(\biu/n1 [40]),
    .i1(uncache_data[40]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[40]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b41  (
    .i0(\biu/n1 [41]),
    .i1(uncache_data[41]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[41]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b42  (
    .i0(\biu/n1 [42]),
    .i1(uncache_data[42]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[42]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b43  (
    .i0(\biu/n1 [43]),
    .i1(uncache_data[43]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[43]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b44  (
    .i0(\biu/n1 [44]),
    .i1(uncache_data[44]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[44]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b45  (
    .i0(\biu/n1 [45]),
    .i1(uncache_data[45]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[45]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b46  (
    .i0(\biu/n1 [46]),
    .i1(uncache_data[46]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[46]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b47  (
    .i0(\biu/n1 [47]),
    .i1(uncache_data[47]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[47]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b48  (
    .i0(\biu/n1 [48]),
    .i1(uncache_data[48]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[48]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b49  (
    .i0(\biu/n1 [49]),
    .i1(uncache_data[49]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[49]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b5  (
    .i0(\biu/n1 [5]),
    .i1(uncache_data[5]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[5]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b50  (
    .i0(\biu/n1 [50]),
    .i1(uncache_data[50]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[50]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b51  (
    .i0(\biu/n1 [51]),
    .i1(uncache_data[51]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[51]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b52  (
    .i0(\biu/n1 [52]),
    .i1(uncache_data[52]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[52]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b53  (
    .i0(\biu/n1 [53]),
    .i1(uncache_data[53]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[53]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b54  (
    .i0(\biu/n1 [54]),
    .i1(uncache_data[54]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[54]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b55  (
    .i0(\biu/n1 [55]),
    .i1(uncache_data[55]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[55]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b56  (
    .i0(\biu/n1 [56]),
    .i1(uncache_data[56]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[56]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b57  (
    .i0(\biu/n1 [57]),
    .i1(uncache_data[57]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[57]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b58  (
    .i0(\biu/n1 [58]),
    .i1(uncache_data[58]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[58]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b59  (
    .i0(\biu/n1 [59]),
    .i1(uncache_data[59]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[59]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b6  (
    .i0(\biu/n1 [6]),
    .i1(uncache_data[6]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[6]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b60  (
    .i0(\biu/n1 [60]),
    .i1(uncache_data[60]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[60]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b61  (
    .i0(\biu/n1 [61]),
    .i1(uncache_data[61]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[61]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b62  (
    .i0(\biu/n1 [62]),
    .i1(uncache_data[62]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[62]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b63  (
    .i0(\biu/n1 [63]),
    .i1(uncache_data[63]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[63]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b7  (
    .i0(\biu/n1 [7]),
    .i1(uncache_data[7]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[7]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b8  (
    .i0(\biu/n1 [8]),
    .i1(uncache_data[8]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[8]));  // ../../RTL/CPU/BIU/biu.v(139)
  binary_mux_s1_w1 \biu/mux5_b9  (
    .i0(\biu/n1 [9]),
    .i1(uncache_data[9]),
    .sel(\biu/ex_data_sel [1]),
    .o(data_read[9]));  // ../../RTL/CPU/BIU/biu.v(139)
  not \biu/opc[1]_inv  (\biu/opc[1]_neg , \biu/opc [1]);
  not \biu/pa_cov_inv  (\biu/pa_cov_neg , \biu/pa_cov );
  not \biu/page_fault_inv  (\biu/page_fault_neg , \biu/page_fault );
  not \biu/wr_inv  (\biu/wr_neg , \biu/wr );
  add_pu60_pu60_o61 \cu_ru/add0_2  (
    .i0(\cu_ru/tvec [63:4]),
    .i1({56'b00000000000000000000000000000000000000000000000000000000,\cu_ru/trap_cause [3:0]}),
    .o({\cu_ru/add0_2_co ,\cu_ru/n43 [59:0]}));  // ../../RTL/CPU/CU&RU/cu_ru.v(357)
  EG_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(64),
    .DATA_WIDTH_W(64))
    \cu_ru/al_ram_gpr  (
    .di(data_rd),
    .raddr(\cu_ru/n46 ),
    .waddr(\cu_ru/n52 ),
    .wclk(clk),
    .we(\cu_ru/n53 ),
    .do(\cu_ru/n47 ));
  EG_LOGIC_DRAM #(
    .ADDR_WIDTH_R(5),
    .ADDR_WIDTH_W(5),
    .DATA_DEPTH_R(32),
    .DATA_DEPTH_W(32),
    .DATA_WIDTH_R(64),
    .DATA_WIDTH_W(64))
    \cu_ru/al_ram_gpr_al_u0  (
    .di(data_rd),
    .raddr(\cu_ru/n49 ),
    .waddr(\cu_ru/n52 ),
    .wclk(clk),
    .we(\cu_ru/n53 ),
    .do(\cu_ru/n50 ));
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b0  (
    .clk(clk),
    .d(data_csr[0]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[0]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b1  (
    .clk(clk),
    .d(data_csr[1]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[1]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b10  (
    .clk(clk),
    .d(data_csr[10]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[10]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b11  (
    .clk(clk),
    .d(data_csr[11]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[11]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b12  (
    .clk(clk),
    .d(data_csr[12]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[12]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b13  (
    .clk(clk),
    .d(data_csr[13]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[13]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b14  (
    .clk(clk),
    .d(data_csr[14]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[14]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b15  (
    .clk(clk),
    .d(data_csr[15]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[15]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b16  (
    .clk(clk),
    .d(data_csr[16]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[16]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b17  (
    .clk(clk),
    .d(data_csr[17]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[17]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b18  (
    .clk(clk),
    .d(data_csr[18]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[18]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b19  (
    .clk(clk),
    .d(data_csr[19]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[19]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b2  (
    .clk(clk),
    .d(data_csr[2]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[2]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b20  (
    .clk(clk),
    .d(data_csr[20]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[20]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b21  (
    .clk(clk),
    .d(data_csr[21]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[21]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b22  (
    .clk(clk),
    .d(data_csr[22]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[22]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b23  (
    .clk(clk),
    .d(data_csr[23]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[23]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b24  (
    .clk(clk),
    .d(data_csr[24]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[24]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b25  (
    .clk(clk),
    .d(data_csr[25]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[25]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b26  (
    .clk(clk),
    .d(data_csr[26]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[26]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b27  (
    .clk(clk),
    .d(data_csr[27]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[27]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b28  (
    .clk(clk),
    .d(data_csr[28]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[28]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b29  (
    .clk(clk),
    .d(data_csr[29]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[29]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b3  (
    .clk(clk),
    .d(data_csr[3]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[3]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b30  (
    .clk(clk),
    .d(data_csr[30]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[30]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b31  (
    .clk(clk),
    .d(data_csr[31]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[31]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b32  (
    .clk(clk),
    .d(data_csr[32]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[32]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b33  (
    .clk(clk),
    .d(data_csr[33]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[33]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b34  (
    .clk(clk),
    .d(data_csr[34]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[34]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b35  (
    .clk(clk),
    .d(data_csr[35]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[35]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b36  (
    .clk(clk),
    .d(data_csr[36]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[36]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b37  (
    .clk(clk),
    .d(data_csr[37]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[37]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b38  (
    .clk(clk),
    .d(data_csr[38]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[38]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b39  (
    .clk(clk),
    .d(data_csr[39]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[39]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b4  (
    .clk(clk),
    .d(data_csr[4]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[4]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b40  (
    .clk(clk),
    .d(data_csr[40]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[40]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b41  (
    .clk(clk),
    .d(data_csr[41]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[41]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b42  (
    .clk(clk),
    .d(data_csr[42]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[42]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b43  (
    .clk(clk),
    .d(data_csr[43]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[43]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b5  (
    .clk(clk),
    .d(data_csr[5]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[5]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b6  (
    .clk(clk),
    .d(data_csr[6]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[6]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b7  (
    .clk(clk),
    .d(data_csr[7]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[7]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b8  (
    .clk(clk),
    .d(data_csr[8]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[8]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg0_b9  (
    .clk(clk),
    .d(data_csr[9]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[9]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg1_b0  (
    .clk(clk),
    .d(data_csr[60]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[60]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg1_b1  (
    .clk(clk),
    .d(data_csr[61]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[61]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg1_b2  (
    .clk(clk),
    .d(data_csr[62]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[62]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  reg_sr_as_w1 \cu_ru/csr_satp/reg1_b3  (
    .clk(clk),
    .d(data_csr[63]),
    .en(\cu_ru/csr_satp/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(satp[63]));  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(25)
  and \cu_ru/csr_satp/u4  (\cu_ru/csr_satp/n0 , \cu_ru/srw_satp_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/csr_satp.v(21)
  eq_w12 \cu_ru/eq0  (
    .i0(csr_index),
    .i1(12'b000100000000),
    .o(\cu_ru/n0 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(264)
  eq_w12 \cu_ru/eq1  (
    .i0(csr_index),
    .i1(12'b000100000100),
    .o(\cu_ru/n1 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(265)
  eq_w12 \cu_ru/eq10  (
    .i0(csr_index),
    .i1(12'b001100000010),
    .o(\cu_ru/n10 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(280)
  eq_w12 \cu_ru/eq11  (
    .i0(csr_index),
    .i1(12'b001100000011),
    .o(\cu_ru/n11 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(281)
  eq_w12 \cu_ru/eq12  (
    .i0(csr_index),
    .i1(12'b001100000100),
    .o(\cu_ru/n12 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(282)
  eq_w12 \cu_ru/eq13  (
    .i0(csr_index),
    .i1(12'b001100000101),
    .o(\cu_ru/n13 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(283)
  eq_w12 \cu_ru/eq14  (
    .i0(csr_index),
    .i1(12'b001101000000),
    .o(\cu_ru/n14 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(285)
  eq_w12 \cu_ru/eq15  (
    .i0(csr_index),
    .i1(12'b001101000001),
    .o(\cu_ru/n15 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(286)
  eq_w12 \cu_ru/eq16  (
    .i0(csr_index),
    .i1(12'b001101000010),
    .o(\cu_ru/n16 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(287)
  eq_w12 \cu_ru/eq17  (
    .i0(csr_index),
    .i1(12'b001101000011),
    .o(\cu_ru/n17 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(288)
  eq_w12 \cu_ru/eq18  (
    .i0(csr_index),
    .i1(12'b001101000100),
    .o(\cu_ru/n18 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(289)
  eq_w12 \cu_ru/eq19  (
    .i0(csr_index),
    .i1(12'b101100000000),
    .o(\cu_ru/n19 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(293)
  eq_w12 \cu_ru/eq2  (
    .i0(csr_index),
    .i1(12'b000100000101),
    .o(\cu_ru/n2 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(266)
  eq_w12 \cu_ru/eq20  (
    .i0(csr_index),
    .i1(12'b001100100000),
    .o(\cu_ru/n20 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(297)
  eq_w12 \cu_ru/eq21  (
    .i0(id_ins[31:20]),
    .i1(12'b110000000000),
    .o(\cu_ru/read_cycle_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(300)
  eq_w12 \cu_ru/eq22  (
    .i0(id_ins[31:20]),
    .i1(12'b110000000001),
    .o(\cu_ru/read_time_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(301)
  eq_w12 \cu_ru/eq23  (
    .i0(id_ins[31:20]),
    .i1(12'b110000000010),
    .o(\cu_ru/read_instret_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(302)
  eq_w12 \cu_ru/eq24  (
    .i0(id_ins[31:20]),
    .i1(12'b000100000000),
    .o(\cu_ru/read_sstatus_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(305)
  eq_w12 \cu_ru/eq25  (
    .i0(id_ins[31:20]),
    .i1(12'b000100000100),
    .o(\cu_ru/read_sie_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(306)
  eq_w12 \cu_ru/eq26  (
    .i0(id_ins[31:20]),
    .i1(12'b000100000101),
    .o(\cu_ru/read_stvec_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(307)
  eq_w12 \cu_ru/eq27  (
    .i0(id_ins[31:20]),
    .i1(12'b000101000000),
    .o(\cu_ru/read_sscratch_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(309)
  eq_w12 \cu_ru/eq28  (
    .i0(id_ins[31:20]),
    .i1(12'b000101000001),
    .o(\cu_ru/read_sepc_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(310)
  eq_w12 \cu_ru/eq29  (
    .i0(id_ins[31:20]),
    .i1(12'b000101000010),
    .o(\cu_ru/read_scause_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(311)
  eq_w12 \cu_ru/eq3  (
    .i0(csr_index),
    .i1(12'b000101000000),
    .o(\cu_ru/n3 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(268)
  eq_w12 \cu_ru/eq30  (
    .i0(id_ins[31:20]),
    .i1(12'b000101000011),
    .o(\cu_ru/read_stval_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(312)
  eq_w12 \cu_ru/eq31  (
    .i0(id_ins[31:20]),
    .i1(12'b000101000100),
    .o(\cu_ru/read_sip_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(313)
  eq_w12 \cu_ru/eq32  (
    .i0(id_ins[31:20]),
    .i1(12'b000110000000),
    .o(\cu_ru/read_satp_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(314)
  eq_w12 \cu_ru/eq33  (
    .i0(id_ins[31:20]),
    .i1(12'b111100010001),
    .o(\cu_ru/read_mvendorid_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(315)
  eq_w12 \cu_ru/eq34  (
    .i0(id_ins[31:20]),
    .i1(12'b111100010010),
    .o(\cu_ru/read_marchid_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(316)
  eq_w12 \cu_ru/eq35  (
    .i0(id_ins[31:20]),
    .i1(12'b111100010011),
    .o(\cu_ru/read_mimp_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(317)
  eq_w12 \cu_ru/eq37  (
    .i0(id_ins[31:20]),
    .i1(12'b001100000000),
    .o(\cu_ru/read_mstatus_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(319)
  eq_w12 \cu_ru/eq39  (
    .i0(id_ins[31:20]),
    .i1(12'b001100000010),
    .o(\cu_ru/read_medeleg_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(321)
  eq_w12 \cu_ru/eq4  (
    .i0(csr_index),
    .i1(12'b000101000001),
    .o(\cu_ru/n4 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(269)
  eq_w12 \cu_ru/eq40  (
    .i0(id_ins[31:20]),
    .i1(12'b001100000011),
    .o(\cu_ru/read_mideleg_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(322)
  eq_w12 \cu_ru/eq41  (
    .i0(id_ins[31:20]),
    .i1(12'b001100000100),
    .o(\cu_ru/read_mie_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(323)
  eq_w12 \cu_ru/eq42  (
    .i0(id_ins[31:20]),
    .i1(12'b001100000101),
    .o(\cu_ru/read_mtvec_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(324)
  eq_w12 \cu_ru/eq43  (
    .i0(id_ins[31:20]),
    .i1(12'b001101000000),
    .o(\cu_ru/read_mscratch_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(326)
  eq_w12 \cu_ru/eq44  (
    .i0(id_ins[31:20]),
    .i1(12'b001101000001),
    .o(\cu_ru/read_mepc_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(327)
  eq_w12 \cu_ru/eq45  (
    .i0(id_ins[31:20]),
    .i1(12'b001101000010),
    .o(\cu_ru/read_mcause_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(328)
  eq_w12 \cu_ru/eq46  (
    .i0(id_ins[31:20]),
    .i1(12'b001101000011),
    .o(\cu_ru/read_mtval_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(329)
  eq_w12 \cu_ru/eq47  (
    .i0(id_ins[31:20]),
    .i1(12'b001101000100),
    .o(\cu_ru/read_mip_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(330)
  eq_w12 \cu_ru/eq48  (
    .i0(id_ins[31:20]),
    .i1(12'b101100000000),
    .o(\cu_ru/read_mcycle_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(334)
  eq_w12 \cu_ru/eq49  (
    .i0(id_ins[31:20]),
    .i1(12'b101100000010),
    .o(\cu_ru/read_minstret_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(335)
  eq_w12 \cu_ru/eq5  (
    .i0(csr_index),
    .i1(12'b000101000010),
    .o(\cu_ru/n5 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(270)
  eq_w12 \cu_ru/eq50  (
    .i0(id_ins[31:20]),
    .i1(12'b001100100000),
    .o(\cu_ru/read_mcounterinhibit_sel ));  // ../../RTL/CPU/CU&RU/cu_ru.v(338)
  eq_w5 \cu_ru/eq51  (
    .i0(id_rs1_index),
    .i1(5'b00000),
    .o(\cu_ru/n45 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  eq_w5 \cu_ru/eq52  (
    .i0(id_rs2_index),
    .i1(5'b00000),
    .o(\cu_ru/n48 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  eq_w12 \cu_ru/eq6  (
    .i0(csr_index),
    .i1(12'b000101000011),
    .o(\cu_ru/n6 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(271)
  eq_w12 \cu_ru/eq7  (
    .i0(csr_index),
    .i1(12'b000101000100),
    .o(\cu_ru/n7 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(272)
  eq_w12 \cu_ru/eq8  (
    .i0(csr_index),
    .i1(12'b000110000000),
    .o(\cu_ru/n8 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(273)
  eq_w12 \cu_ru/eq9  (
    .i0(csr_index),
    .i1(12'b001100000000),
    .o(\cu_ru/n9 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(278)
  not \cu_ru/exception_inv  (\cu_ru/exception_neg , \cu_ru/exception );
  add_pu64_pu64_o64 \cu_ru/m_cycle_event/add0  (
    .i0(\cu_ru/mcycle ),
    .i1(64'b0000000000000000000000000000000000000000000000000000000000000001),
    .o(\cu_ru/m_cycle_event/n2 ));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  add_pu64_pu64_o64 \cu_ru/m_cycle_event/add1  (
    .i0(\cu_ru/minstret ),
    .i1(64'b0000000000000000000000000000000000000000000000000000000000000001),
    .o(\cu_ru/m_cycle_event/n4 ));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(38)
  reg_sr_as_w1 \cu_ru/m_cycle_event/cy_reg  (
    .clk(clk),
    .d(data_csr[0]),
    .en(\cu_ru/m_cycle_event/n13 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcountinhibit ));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(51)
  reg_sr_as_w1 \cu_ru/m_cycle_event/ir_reg  (
    .clk(clk),
    .d(data_csr[2]),
    .en(\cu_ru/m_cycle_event/n13 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_cycle_event/mcountinhibit[2] ));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(51)
  not \cu_ru/m_cycle_event/mcountinhibit[2]_inv  (\cu_ru/m_cycle_event/mcountinhibit[2]_neg , \cu_ru/m_cycle_event/mcountinhibit[2] );
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b0  (
    .i0(\cu_ru/m_cycle_event/n2 [0]),
    .i1(\cu_ru/mcycle [0]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b1  (
    .i0(\cu_ru/m_cycle_event/n2 [1]),
    .i1(\cu_ru/mcycle [1]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b10  (
    .i0(\cu_ru/m_cycle_event/n2 [10]),
    .i1(\cu_ru/mcycle [10]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b11  (
    .i0(\cu_ru/m_cycle_event/n2 [11]),
    .i1(\cu_ru/mcycle [11]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b12  (
    .i0(\cu_ru/m_cycle_event/n2 [12]),
    .i1(\cu_ru/mcycle [12]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b13  (
    .i0(\cu_ru/m_cycle_event/n2 [13]),
    .i1(\cu_ru/mcycle [13]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b14  (
    .i0(\cu_ru/m_cycle_event/n2 [14]),
    .i1(\cu_ru/mcycle [14]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b15  (
    .i0(\cu_ru/m_cycle_event/n2 [15]),
    .i1(\cu_ru/mcycle [15]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b16  (
    .i0(\cu_ru/m_cycle_event/n2 [16]),
    .i1(\cu_ru/mcycle [16]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b17  (
    .i0(\cu_ru/m_cycle_event/n2 [17]),
    .i1(\cu_ru/mcycle [17]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b18  (
    .i0(\cu_ru/m_cycle_event/n2 [18]),
    .i1(\cu_ru/mcycle [18]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b19  (
    .i0(\cu_ru/m_cycle_event/n2 [19]),
    .i1(\cu_ru/mcycle [19]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b2  (
    .i0(\cu_ru/m_cycle_event/n2 [2]),
    .i1(\cu_ru/mcycle [2]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b20  (
    .i0(\cu_ru/m_cycle_event/n2 [20]),
    .i1(\cu_ru/mcycle [20]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b21  (
    .i0(\cu_ru/m_cycle_event/n2 [21]),
    .i1(\cu_ru/mcycle [21]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b22  (
    .i0(\cu_ru/m_cycle_event/n2 [22]),
    .i1(\cu_ru/mcycle [22]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b23  (
    .i0(\cu_ru/m_cycle_event/n2 [23]),
    .i1(\cu_ru/mcycle [23]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b24  (
    .i0(\cu_ru/m_cycle_event/n2 [24]),
    .i1(\cu_ru/mcycle [24]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b25  (
    .i0(\cu_ru/m_cycle_event/n2 [25]),
    .i1(\cu_ru/mcycle [25]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b26  (
    .i0(\cu_ru/m_cycle_event/n2 [26]),
    .i1(\cu_ru/mcycle [26]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b27  (
    .i0(\cu_ru/m_cycle_event/n2 [27]),
    .i1(\cu_ru/mcycle [27]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b28  (
    .i0(\cu_ru/m_cycle_event/n2 [28]),
    .i1(\cu_ru/mcycle [28]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b29  (
    .i0(\cu_ru/m_cycle_event/n2 [29]),
    .i1(\cu_ru/mcycle [29]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b3  (
    .i0(\cu_ru/m_cycle_event/n2 [3]),
    .i1(\cu_ru/mcycle [3]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b30  (
    .i0(\cu_ru/m_cycle_event/n2 [30]),
    .i1(\cu_ru/mcycle [30]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b31  (
    .i0(\cu_ru/m_cycle_event/n2 [31]),
    .i1(\cu_ru/mcycle [31]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b32  (
    .i0(\cu_ru/m_cycle_event/n2 [32]),
    .i1(\cu_ru/mcycle [32]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b33  (
    .i0(\cu_ru/m_cycle_event/n2 [33]),
    .i1(\cu_ru/mcycle [33]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b34  (
    .i0(\cu_ru/m_cycle_event/n2 [34]),
    .i1(\cu_ru/mcycle [34]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b35  (
    .i0(\cu_ru/m_cycle_event/n2 [35]),
    .i1(\cu_ru/mcycle [35]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b36  (
    .i0(\cu_ru/m_cycle_event/n2 [36]),
    .i1(\cu_ru/mcycle [36]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b37  (
    .i0(\cu_ru/m_cycle_event/n2 [37]),
    .i1(\cu_ru/mcycle [37]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b38  (
    .i0(\cu_ru/m_cycle_event/n2 [38]),
    .i1(\cu_ru/mcycle [38]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b39  (
    .i0(\cu_ru/m_cycle_event/n2 [39]),
    .i1(\cu_ru/mcycle [39]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b4  (
    .i0(\cu_ru/m_cycle_event/n2 [4]),
    .i1(\cu_ru/mcycle [4]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b40  (
    .i0(\cu_ru/m_cycle_event/n2 [40]),
    .i1(\cu_ru/mcycle [40]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b41  (
    .i0(\cu_ru/m_cycle_event/n2 [41]),
    .i1(\cu_ru/mcycle [41]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b42  (
    .i0(\cu_ru/m_cycle_event/n2 [42]),
    .i1(\cu_ru/mcycle [42]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b43  (
    .i0(\cu_ru/m_cycle_event/n2 [43]),
    .i1(\cu_ru/mcycle [43]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b44  (
    .i0(\cu_ru/m_cycle_event/n2 [44]),
    .i1(\cu_ru/mcycle [44]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b45  (
    .i0(\cu_ru/m_cycle_event/n2 [45]),
    .i1(\cu_ru/mcycle [45]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b46  (
    .i0(\cu_ru/m_cycle_event/n2 [46]),
    .i1(\cu_ru/mcycle [46]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b47  (
    .i0(\cu_ru/m_cycle_event/n2 [47]),
    .i1(\cu_ru/mcycle [47]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b48  (
    .i0(\cu_ru/m_cycle_event/n2 [48]),
    .i1(\cu_ru/mcycle [48]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b49  (
    .i0(\cu_ru/m_cycle_event/n2 [49]),
    .i1(\cu_ru/mcycle [49]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b5  (
    .i0(\cu_ru/m_cycle_event/n2 [5]),
    .i1(\cu_ru/mcycle [5]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b50  (
    .i0(\cu_ru/m_cycle_event/n2 [50]),
    .i1(\cu_ru/mcycle [50]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b51  (
    .i0(\cu_ru/m_cycle_event/n2 [51]),
    .i1(\cu_ru/mcycle [51]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b52  (
    .i0(\cu_ru/m_cycle_event/n2 [52]),
    .i1(\cu_ru/mcycle [52]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b53  (
    .i0(\cu_ru/m_cycle_event/n2 [53]),
    .i1(\cu_ru/mcycle [53]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b54  (
    .i0(\cu_ru/m_cycle_event/n2 [54]),
    .i1(\cu_ru/mcycle [54]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b55  (
    .i0(\cu_ru/m_cycle_event/n2 [55]),
    .i1(\cu_ru/mcycle [55]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b56  (
    .i0(\cu_ru/m_cycle_event/n2 [56]),
    .i1(\cu_ru/mcycle [56]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b57  (
    .i0(\cu_ru/m_cycle_event/n2 [57]),
    .i1(\cu_ru/mcycle [57]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b58  (
    .i0(\cu_ru/m_cycle_event/n2 [58]),
    .i1(\cu_ru/mcycle [58]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b59  (
    .i0(\cu_ru/m_cycle_event/n2 [59]),
    .i1(\cu_ru/mcycle [59]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b6  (
    .i0(\cu_ru/m_cycle_event/n2 [6]),
    .i1(\cu_ru/mcycle [6]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b60  (
    .i0(\cu_ru/m_cycle_event/n2 [60]),
    .i1(\cu_ru/mcycle [60]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b61  (
    .i0(\cu_ru/m_cycle_event/n2 [61]),
    .i1(\cu_ru/mcycle [61]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b62  (
    .i0(\cu_ru/m_cycle_event/n2 [62]),
    .i1(\cu_ru/mcycle [62]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b63  (
    .i0(\cu_ru/m_cycle_event/n2 [63]),
    .i1(\cu_ru/mcycle [63]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b7  (
    .i0(\cu_ru/m_cycle_event/n2 [7]),
    .i1(\cu_ru/mcycle [7]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b8  (
    .i0(\cu_ru/m_cycle_event/n2 [8]),
    .i1(\cu_ru/mcycle [8]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux0_b9  (
    .i0(\cu_ru/m_cycle_event/n2 [9]),
    .i1(\cu_ru/mcycle [9]),
    .sel(\cu_ru/mcountinhibit ),
    .o(\cu_ru/m_cycle_event/n3 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(37)
  and \cu_ru/m_cycle_event/mux2_b0_sel_is_2  (\cu_ru/m_cycle_event/mux2_b0_sel_is_2_o , \cu_ru/m_cycle_event/mcountinhibit[2]_neg , wb_valid);
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b0  (
    .i0(\cu_ru/m_cycle_event/n3 [0]),
    .i1(data_csr[0]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b1  (
    .i0(\cu_ru/m_cycle_event/n3 [1]),
    .i1(data_csr[1]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b10  (
    .i0(\cu_ru/m_cycle_event/n3 [10]),
    .i1(data_csr[10]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b11  (
    .i0(\cu_ru/m_cycle_event/n3 [11]),
    .i1(data_csr[11]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b12  (
    .i0(\cu_ru/m_cycle_event/n3 [12]),
    .i1(data_csr[12]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b13  (
    .i0(\cu_ru/m_cycle_event/n3 [13]),
    .i1(data_csr[13]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b14  (
    .i0(\cu_ru/m_cycle_event/n3 [14]),
    .i1(data_csr[14]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b15  (
    .i0(\cu_ru/m_cycle_event/n3 [15]),
    .i1(data_csr[15]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b16  (
    .i0(\cu_ru/m_cycle_event/n3 [16]),
    .i1(data_csr[16]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b17  (
    .i0(\cu_ru/m_cycle_event/n3 [17]),
    .i1(data_csr[17]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b18  (
    .i0(\cu_ru/m_cycle_event/n3 [18]),
    .i1(data_csr[18]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b19  (
    .i0(\cu_ru/m_cycle_event/n3 [19]),
    .i1(data_csr[19]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b2  (
    .i0(\cu_ru/m_cycle_event/n3 [2]),
    .i1(data_csr[2]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b20  (
    .i0(\cu_ru/m_cycle_event/n3 [20]),
    .i1(data_csr[20]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b21  (
    .i0(\cu_ru/m_cycle_event/n3 [21]),
    .i1(data_csr[21]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b22  (
    .i0(\cu_ru/m_cycle_event/n3 [22]),
    .i1(data_csr[22]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b23  (
    .i0(\cu_ru/m_cycle_event/n3 [23]),
    .i1(data_csr[23]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b24  (
    .i0(\cu_ru/m_cycle_event/n3 [24]),
    .i1(data_csr[24]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b25  (
    .i0(\cu_ru/m_cycle_event/n3 [25]),
    .i1(data_csr[25]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b26  (
    .i0(\cu_ru/m_cycle_event/n3 [26]),
    .i1(data_csr[26]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b27  (
    .i0(\cu_ru/m_cycle_event/n3 [27]),
    .i1(data_csr[27]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b28  (
    .i0(\cu_ru/m_cycle_event/n3 [28]),
    .i1(data_csr[28]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b29  (
    .i0(\cu_ru/m_cycle_event/n3 [29]),
    .i1(data_csr[29]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b3  (
    .i0(\cu_ru/m_cycle_event/n3 [3]),
    .i1(data_csr[3]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b30  (
    .i0(\cu_ru/m_cycle_event/n3 [30]),
    .i1(data_csr[30]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b31  (
    .i0(\cu_ru/m_cycle_event/n3 [31]),
    .i1(data_csr[31]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b32  (
    .i0(\cu_ru/m_cycle_event/n3 [32]),
    .i1(data_csr[32]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b33  (
    .i0(\cu_ru/m_cycle_event/n3 [33]),
    .i1(data_csr[33]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b34  (
    .i0(\cu_ru/m_cycle_event/n3 [34]),
    .i1(data_csr[34]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b35  (
    .i0(\cu_ru/m_cycle_event/n3 [35]),
    .i1(data_csr[35]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b36  (
    .i0(\cu_ru/m_cycle_event/n3 [36]),
    .i1(data_csr[36]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b37  (
    .i0(\cu_ru/m_cycle_event/n3 [37]),
    .i1(data_csr[37]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b38  (
    .i0(\cu_ru/m_cycle_event/n3 [38]),
    .i1(data_csr[38]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b39  (
    .i0(\cu_ru/m_cycle_event/n3 [39]),
    .i1(data_csr[39]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b4  (
    .i0(\cu_ru/m_cycle_event/n3 [4]),
    .i1(data_csr[4]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b40  (
    .i0(\cu_ru/m_cycle_event/n3 [40]),
    .i1(data_csr[40]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b41  (
    .i0(\cu_ru/m_cycle_event/n3 [41]),
    .i1(data_csr[41]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b42  (
    .i0(\cu_ru/m_cycle_event/n3 [42]),
    .i1(data_csr[42]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b43  (
    .i0(\cu_ru/m_cycle_event/n3 [43]),
    .i1(data_csr[43]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b44  (
    .i0(\cu_ru/m_cycle_event/n3 [44]),
    .i1(data_csr[44]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b45  (
    .i0(\cu_ru/m_cycle_event/n3 [45]),
    .i1(data_csr[45]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b46  (
    .i0(\cu_ru/m_cycle_event/n3 [46]),
    .i1(data_csr[46]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b47  (
    .i0(\cu_ru/m_cycle_event/n3 [47]),
    .i1(data_csr[47]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b48  (
    .i0(\cu_ru/m_cycle_event/n3 [48]),
    .i1(data_csr[48]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b49  (
    .i0(\cu_ru/m_cycle_event/n3 [49]),
    .i1(data_csr[49]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b5  (
    .i0(\cu_ru/m_cycle_event/n3 [5]),
    .i1(data_csr[5]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b50  (
    .i0(\cu_ru/m_cycle_event/n3 [50]),
    .i1(data_csr[50]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b51  (
    .i0(\cu_ru/m_cycle_event/n3 [51]),
    .i1(data_csr[51]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b52  (
    .i0(\cu_ru/m_cycle_event/n3 [52]),
    .i1(data_csr[52]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b53  (
    .i0(\cu_ru/m_cycle_event/n3 [53]),
    .i1(data_csr[53]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b54  (
    .i0(\cu_ru/m_cycle_event/n3 [54]),
    .i1(data_csr[54]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b55  (
    .i0(\cu_ru/m_cycle_event/n3 [55]),
    .i1(data_csr[55]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b56  (
    .i0(\cu_ru/m_cycle_event/n3 [56]),
    .i1(data_csr[56]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b57  (
    .i0(\cu_ru/m_cycle_event/n3 [57]),
    .i1(data_csr[57]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b58  (
    .i0(\cu_ru/m_cycle_event/n3 [58]),
    .i1(data_csr[58]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b59  (
    .i0(\cu_ru/m_cycle_event/n3 [59]),
    .i1(data_csr[59]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b6  (
    .i0(\cu_ru/m_cycle_event/n3 [6]),
    .i1(data_csr[6]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b60  (
    .i0(\cu_ru/m_cycle_event/n3 [60]),
    .i1(data_csr[60]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b61  (
    .i0(\cu_ru/m_cycle_event/n3 [61]),
    .i1(data_csr[61]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b62  (
    .i0(\cu_ru/m_cycle_event/n3 [62]),
    .i1(data_csr[62]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b63  (
    .i0(\cu_ru/m_cycle_event/n3 [63]),
    .i1(data_csr[63]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b7  (
    .i0(\cu_ru/m_cycle_event/n3 [7]),
    .i1(data_csr[7]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b8  (
    .i0(\cu_ru/m_cycle_event/n3 [8]),
    .i1(data_csr[8]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  binary_mux_s1_w1 \cu_ru/m_cycle_event/mux5_b9  (
    .i0(\cu_ru/m_cycle_event/n3 [9]),
    .i1(data_csr[9]),
    .sel(\cu_ru/m_cycle_event/n0 ),
    .o(\cu_ru/m_cycle_event/n9 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(39)
  and \cu_ru/m_cycle_event/mux6_b0_sel_is_2  (\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o , \cu_ru/m_cycle_event/n0_neg , \cu_ru/m_cycle_event/mux2_b0_sel_is_2_o );
  not \cu_ru/m_cycle_event/n0_inv  (\cu_ru/m_cycle_event/n0_neg , \cu_ru/m_cycle_event/n0 );
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b0  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [0]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [0]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b1  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [1]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [1]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b10  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [10]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [10]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b11  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [11]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [11]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b12  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [12]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [12]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b13  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [13]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [13]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b14  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [14]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [14]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b15  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [15]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [15]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b16  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [16]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [16]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b17  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [17]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [17]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b18  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [18]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [18]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b19  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [19]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [19]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b2  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [2]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [2]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b20  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [20]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [20]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b21  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [21]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [21]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b22  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [22]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [22]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b23  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [23]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [23]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b24  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [24]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [24]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b25  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [25]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [25]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b26  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [26]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [26]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b27  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [27]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [27]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b28  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [28]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [28]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b29  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [29]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [29]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b3  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [3]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [3]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b30  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [30]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [30]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b31  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [31]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [31]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b32  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [32]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [32]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b33  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [33]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [33]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b34  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [34]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [34]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b35  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [35]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [35]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b36  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [36]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [36]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b37  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [37]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [37]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b38  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [38]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [38]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b39  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [39]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [39]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b4  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [4]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [4]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b40  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [40]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [40]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b41  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [41]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [41]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b42  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [42]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [42]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b43  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [43]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [43]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b44  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [44]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [44]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b45  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [45]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [45]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b46  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [46]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [46]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b47  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [47]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [47]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b48  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [48]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [48]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b49  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [49]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [49]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b5  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [5]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [5]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b50  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [50]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [50]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b51  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [51]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [51]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b52  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [52]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [52]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b53  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [53]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [53]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b54  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [54]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [54]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b55  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [55]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [55]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b56  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [56]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [56]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b57  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [57]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [57]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b58  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [58]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [58]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b59  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [59]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [59]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b6  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [6]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [6]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b60  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [60]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [60]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b61  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [61]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [61]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b62  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [62]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [62]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b63  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [63]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [63]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b7  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [7]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [7]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b8  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [8]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [8]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg0_b9  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n4 [9]),
    .en(\cu_ru/m_cycle_event/mux6_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/minstret [9]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b0  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [0]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b1  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [1]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b10  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [10]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b11  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [11]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b12  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [12]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b13  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [13]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b14  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [14]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b15  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [15]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b16  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [16]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b17  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [17]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b18  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [18]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b19  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [19]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b2  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [2]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b20  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [20]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b21  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [21]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b22  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [22]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b23  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [23]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b24  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [24]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b25  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [25]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b26  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [26]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b27  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [27]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b28  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [28]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b29  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [29]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b3  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [3]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b30  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [30]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b31  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [31]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b32  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [32]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b33  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [33]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b34  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [34]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b35  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [35]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b36  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [36]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b37  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [37]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b38  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [38]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b39  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [39]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b4  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [4]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b40  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [40]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b41  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [41]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b42  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [42]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b43  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [43]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b44  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [44]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b45  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [45]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b46  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [46]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b47  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [47]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b48  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [48]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b49  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [49]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b5  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [5]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b50  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [50]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b51  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [51]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b52  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [52]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b53  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [53]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b54  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [54]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b55  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [55]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b56  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [56]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b57  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [57]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b58  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [58]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b59  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [59]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b6  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [6]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b60  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [60]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b61  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [61]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b62  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [62]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b63  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [63]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b7  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [7]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b8  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [8]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  reg_sr_as_w1 \cu_ru/m_cycle_event/reg1_b9  (
    .clk(clk),
    .d(\cu_ru/m_cycle_event/n9 [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcycle [9]));  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(40)
  and \cu_ru/m_cycle_event/u4  (\cu_ru/m_cycle_event/n0 , \cu_ru/mrw_mcycle_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(30)
  and \cu_ru/m_cycle_event/u8  (\cu_ru/m_cycle_event/n13 , \cu_ru/mrw_mcounterinhibit_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_cycle_event.v(47)
  AL_MUX \cu_ru/m_s_cause/mux2_b0  (
    .i0(\cu_ru/scause [0]),
    .i1(data_csr[0]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [0]));
  and \cu_ru/m_s_cause/mux2_b0_sel_is_2  (\cu_ru/m_s_cause/mux2_b0_sel_is_2_o , \cu_ru/m_s_cause/n0_neg , \cu_ru/m_s_cause/n1 );
  AL_MUX \cu_ru/m_s_cause/mux2_b1  (
    .i0(\cu_ru/scause [1]),
    .i1(data_csr[1]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [1]));
  AL_MUX \cu_ru/m_s_cause/mux2_b10  (
    .i0(\cu_ru/scause [10]),
    .i1(data_csr[10]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [10]));
  AL_MUX \cu_ru/m_s_cause/mux2_b11  (
    .i0(\cu_ru/scause [11]),
    .i1(data_csr[11]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [11]));
  AL_MUX \cu_ru/m_s_cause/mux2_b12  (
    .i0(\cu_ru/scause [12]),
    .i1(data_csr[12]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [12]));
  AL_MUX \cu_ru/m_s_cause/mux2_b13  (
    .i0(\cu_ru/scause [13]),
    .i1(data_csr[13]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [13]));
  AL_MUX \cu_ru/m_s_cause/mux2_b14  (
    .i0(\cu_ru/scause [14]),
    .i1(data_csr[14]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [14]));
  AL_MUX \cu_ru/m_s_cause/mux2_b15  (
    .i0(\cu_ru/scause [15]),
    .i1(data_csr[15]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [15]));
  AL_MUX \cu_ru/m_s_cause/mux2_b16  (
    .i0(\cu_ru/scause [16]),
    .i1(data_csr[16]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [16]));
  AL_MUX \cu_ru/m_s_cause/mux2_b17  (
    .i0(\cu_ru/scause [17]),
    .i1(data_csr[17]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [17]));
  AL_MUX \cu_ru/m_s_cause/mux2_b18  (
    .i0(\cu_ru/scause [18]),
    .i1(data_csr[18]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [18]));
  AL_MUX \cu_ru/m_s_cause/mux2_b19  (
    .i0(\cu_ru/scause [19]),
    .i1(data_csr[19]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [19]));
  AL_MUX \cu_ru/m_s_cause/mux2_b2  (
    .i0(\cu_ru/scause [2]),
    .i1(data_csr[2]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [2]));
  AL_MUX \cu_ru/m_s_cause/mux2_b20  (
    .i0(\cu_ru/scause [20]),
    .i1(data_csr[20]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [20]));
  AL_MUX \cu_ru/m_s_cause/mux2_b21  (
    .i0(\cu_ru/scause [21]),
    .i1(data_csr[21]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [21]));
  AL_MUX \cu_ru/m_s_cause/mux2_b22  (
    .i0(\cu_ru/scause [22]),
    .i1(data_csr[22]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [22]));
  AL_MUX \cu_ru/m_s_cause/mux2_b23  (
    .i0(\cu_ru/scause [23]),
    .i1(data_csr[23]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [23]));
  AL_MUX \cu_ru/m_s_cause/mux2_b24  (
    .i0(\cu_ru/scause [24]),
    .i1(data_csr[24]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [24]));
  AL_MUX \cu_ru/m_s_cause/mux2_b25  (
    .i0(\cu_ru/scause [25]),
    .i1(data_csr[25]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [25]));
  AL_MUX \cu_ru/m_s_cause/mux2_b26  (
    .i0(\cu_ru/scause [26]),
    .i1(data_csr[26]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [26]));
  AL_MUX \cu_ru/m_s_cause/mux2_b27  (
    .i0(\cu_ru/scause [27]),
    .i1(data_csr[27]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [27]));
  AL_MUX \cu_ru/m_s_cause/mux2_b28  (
    .i0(\cu_ru/scause [28]),
    .i1(data_csr[28]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [28]));
  AL_MUX \cu_ru/m_s_cause/mux2_b29  (
    .i0(\cu_ru/scause [29]),
    .i1(data_csr[29]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [29]));
  AL_MUX \cu_ru/m_s_cause/mux2_b3  (
    .i0(\cu_ru/scause [3]),
    .i1(data_csr[3]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [3]));
  AL_MUX \cu_ru/m_s_cause/mux2_b30  (
    .i0(\cu_ru/scause [30]),
    .i1(data_csr[30]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [30]));
  AL_MUX \cu_ru/m_s_cause/mux2_b31  (
    .i0(\cu_ru/scause [31]),
    .i1(data_csr[31]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [31]));
  AL_MUX \cu_ru/m_s_cause/mux2_b32  (
    .i0(\cu_ru/scause [32]),
    .i1(data_csr[32]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [32]));
  AL_MUX \cu_ru/m_s_cause/mux2_b33  (
    .i0(\cu_ru/scause [33]),
    .i1(data_csr[33]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [33]));
  AL_MUX \cu_ru/m_s_cause/mux2_b34  (
    .i0(\cu_ru/scause [34]),
    .i1(data_csr[34]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [34]));
  AL_MUX \cu_ru/m_s_cause/mux2_b35  (
    .i0(\cu_ru/scause [35]),
    .i1(data_csr[35]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [35]));
  AL_MUX \cu_ru/m_s_cause/mux2_b36  (
    .i0(\cu_ru/scause [36]),
    .i1(data_csr[36]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [36]));
  AL_MUX \cu_ru/m_s_cause/mux2_b37  (
    .i0(\cu_ru/scause [37]),
    .i1(data_csr[37]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [37]));
  AL_MUX \cu_ru/m_s_cause/mux2_b38  (
    .i0(\cu_ru/scause [38]),
    .i1(data_csr[38]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [38]));
  AL_MUX \cu_ru/m_s_cause/mux2_b39  (
    .i0(\cu_ru/scause [39]),
    .i1(data_csr[39]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [39]));
  AL_MUX \cu_ru/m_s_cause/mux2_b4  (
    .i0(\cu_ru/scause [4]),
    .i1(data_csr[4]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [4]));
  AL_MUX \cu_ru/m_s_cause/mux2_b40  (
    .i0(\cu_ru/scause [40]),
    .i1(data_csr[40]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [40]));
  AL_MUX \cu_ru/m_s_cause/mux2_b41  (
    .i0(\cu_ru/scause [41]),
    .i1(data_csr[41]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [41]));
  AL_MUX \cu_ru/m_s_cause/mux2_b42  (
    .i0(\cu_ru/scause [42]),
    .i1(data_csr[42]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [42]));
  AL_MUX \cu_ru/m_s_cause/mux2_b43  (
    .i0(\cu_ru/scause [43]),
    .i1(data_csr[43]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [43]));
  AL_MUX \cu_ru/m_s_cause/mux2_b44  (
    .i0(\cu_ru/scause [44]),
    .i1(data_csr[44]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [44]));
  AL_MUX \cu_ru/m_s_cause/mux2_b45  (
    .i0(\cu_ru/scause [45]),
    .i1(data_csr[45]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [45]));
  AL_MUX \cu_ru/m_s_cause/mux2_b46  (
    .i0(\cu_ru/scause [46]),
    .i1(data_csr[46]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [46]));
  AL_MUX \cu_ru/m_s_cause/mux2_b47  (
    .i0(\cu_ru/scause [47]),
    .i1(data_csr[47]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [47]));
  AL_MUX \cu_ru/m_s_cause/mux2_b48  (
    .i0(\cu_ru/scause [48]),
    .i1(data_csr[48]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [48]));
  AL_MUX \cu_ru/m_s_cause/mux2_b49  (
    .i0(\cu_ru/scause [49]),
    .i1(data_csr[49]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [49]));
  AL_MUX \cu_ru/m_s_cause/mux2_b5  (
    .i0(\cu_ru/scause [5]),
    .i1(data_csr[5]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [5]));
  AL_MUX \cu_ru/m_s_cause/mux2_b50  (
    .i0(\cu_ru/scause [50]),
    .i1(data_csr[50]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [50]));
  AL_MUX \cu_ru/m_s_cause/mux2_b51  (
    .i0(\cu_ru/scause [51]),
    .i1(data_csr[51]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [51]));
  AL_MUX \cu_ru/m_s_cause/mux2_b52  (
    .i0(\cu_ru/scause [52]),
    .i1(data_csr[52]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [52]));
  AL_MUX \cu_ru/m_s_cause/mux2_b53  (
    .i0(\cu_ru/scause [53]),
    .i1(data_csr[53]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [53]));
  AL_MUX \cu_ru/m_s_cause/mux2_b54  (
    .i0(\cu_ru/scause [54]),
    .i1(data_csr[54]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [54]));
  AL_MUX \cu_ru/m_s_cause/mux2_b55  (
    .i0(\cu_ru/scause [55]),
    .i1(data_csr[55]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [55]));
  AL_MUX \cu_ru/m_s_cause/mux2_b56  (
    .i0(\cu_ru/scause [56]),
    .i1(data_csr[56]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [56]));
  AL_MUX \cu_ru/m_s_cause/mux2_b57  (
    .i0(\cu_ru/scause [57]),
    .i1(data_csr[57]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [57]));
  AL_MUX \cu_ru/m_s_cause/mux2_b58  (
    .i0(\cu_ru/scause [58]),
    .i1(data_csr[58]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [58]));
  AL_MUX \cu_ru/m_s_cause/mux2_b59  (
    .i0(\cu_ru/scause [59]),
    .i1(data_csr[59]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [59]));
  AL_MUX \cu_ru/m_s_cause/mux2_b6  (
    .i0(\cu_ru/scause [6]),
    .i1(data_csr[6]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [6]));
  AL_MUX \cu_ru/m_s_cause/mux2_b60  (
    .i0(\cu_ru/scause [60]),
    .i1(data_csr[60]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [60]));
  AL_MUX \cu_ru/m_s_cause/mux2_b61  (
    .i0(\cu_ru/scause [61]),
    .i1(data_csr[61]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [61]));
  AL_MUX \cu_ru/m_s_cause/mux2_b62  (
    .i0(\cu_ru/scause [62]),
    .i1(data_csr[62]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [62]));
  AL_MUX \cu_ru/m_s_cause/mux2_b63  (
    .i0(\cu_ru/scause [63]),
    .i1(data_csr[63]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [63]));
  AL_MUX \cu_ru/m_s_cause/mux2_b7  (
    .i0(\cu_ru/scause [7]),
    .i1(data_csr[7]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [7]));
  AL_MUX \cu_ru/m_s_cause/mux2_b8  (
    .i0(\cu_ru/scause [8]),
    .i1(data_csr[8]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [8]));
  AL_MUX \cu_ru/m_s_cause/mux2_b9  (
    .i0(\cu_ru/scause [9]),
    .i1(data_csr[9]),
    .sel(\cu_ru/m_s_cause/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n4 [9]));
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b0  (
    .i0(\cu_ru/m_s_cause/n4 [0]),
    .i1(\cu_ru/trap_cause [0]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b1  (
    .i0(\cu_ru/m_s_cause/n4 [1]),
    .i1(\cu_ru/trap_cause [1]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b10  (
    .i0(\cu_ru/m_s_cause/n4 [10]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b11  (
    .i0(\cu_ru/m_s_cause/n4 [11]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b12  (
    .i0(\cu_ru/m_s_cause/n4 [12]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b13  (
    .i0(\cu_ru/m_s_cause/n4 [13]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b14  (
    .i0(\cu_ru/m_s_cause/n4 [14]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b15  (
    .i0(\cu_ru/m_s_cause/n4 [15]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b16  (
    .i0(\cu_ru/m_s_cause/n4 [16]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b17  (
    .i0(\cu_ru/m_s_cause/n4 [17]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b18  (
    .i0(\cu_ru/m_s_cause/n4 [18]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b19  (
    .i0(\cu_ru/m_s_cause/n4 [19]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b2  (
    .i0(\cu_ru/m_s_cause/n4 [2]),
    .i1(\cu_ru/trap_cause [2]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b20  (
    .i0(\cu_ru/m_s_cause/n4 [20]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b21  (
    .i0(\cu_ru/m_s_cause/n4 [21]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b22  (
    .i0(\cu_ru/m_s_cause/n4 [22]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b23  (
    .i0(\cu_ru/m_s_cause/n4 [23]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b24  (
    .i0(\cu_ru/m_s_cause/n4 [24]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b25  (
    .i0(\cu_ru/m_s_cause/n4 [25]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b26  (
    .i0(\cu_ru/m_s_cause/n4 [26]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b27  (
    .i0(\cu_ru/m_s_cause/n4 [27]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b28  (
    .i0(\cu_ru/m_s_cause/n4 [28]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b29  (
    .i0(\cu_ru/m_s_cause/n4 [29]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b3  (
    .i0(\cu_ru/m_s_cause/n4 [3]),
    .i1(\cu_ru/trap_cause [3]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b30  (
    .i0(\cu_ru/m_s_cause/n4 [30]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b31  (
    .i0(\cu_ru/m_s_cause/n4 [31]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b32  (
    .i0(\cu_ru/m_s_cause/n4 [32]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b33  (
    .i0(\cu_ru/m_s_cause/n4 [33]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b34  (
    .i0(\cu_ru/m_s_cause/n4 [34]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b35  (
    .i0(\cu_ru/m_s_cause/n4 [35]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b36  (
    .i0(\cu_ru/m_s_cause/n4 [36]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b37  (
    .i0(\cu_ru/m_s_cause/n4 [37]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b38  (
    .i0(\cu_ru/m_s_cause/n4 [38]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b39  (
    .i0(\cu_ru/m_s_cause/n4 [39]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b4  (
    .i0(\cu_ru/m_s_cause/n4 [4]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b40  (
    .i0(\cu_ru/m_s_cause/n4 [40]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b41  (
    .i0(\cu_ru/m_s_cause/n4 [41]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b42  (
    .i0(\cu_ru/m_s_cause/n4 [42]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b43  (
    .i0(\cu_ru/m_s_cause/n4 [43]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b44  (
    .i0(\cu_ru/m_s_cause/n4 [44]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b45  (
    .i0(\cu_ru/m_s_cause/n4 [45]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b46  (
    .i0(\cu_ru/m_s_cause/n4 [46]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b47  (
    .i0(\cu_ru/m_s_cause/n4 [47]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b48  (
    .i0(\cu_ru/m_s_cause/n4 [48]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b49  (
    .i0(\cu_ru/m_s_cause/n4 [49]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b5  (
    .i0(\cu_ru/m_s_cause/n4 [5]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b50  (
    .i0(\cu_ru/m_s_cause/n4 [50]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b51  (
    .i0(\cu_ru/m_s_cause/n4 [51]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b52  (
    .i0(\cu_ru/m_s_cause/n4 [52]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b53  (
    .i0(\cu_ru/m_s_cause/n4 [53]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b54  (
    .i0(\cu_ru/m_s_cause/n4 [54]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b55  (
    .i0(\cu_ru/m_s_cause/n4 [55]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b56  (
    .i0(\cu_ru/m_s_cause/n4 [56]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b57  (
    .i0(\cu_ru/m_s_cause/n4 [57]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b58  (
    .i0(\cu_ru/m_s_cause/n4 [58]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b59  (
    .i0(\cu_ru/m_s_cause/n4 [59]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b6  (
    .i0(\cu_ru/m_s_cause/n4 [6]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b60  (
    .i0(\cu_ru/m_s_cause/n4 [60]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b61  (
    .i0(\cu_ru/m_s_cause/n4 [61]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b62  (
    .i0(\cu_ru/m_s_cause/n4 [62]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b63  (
    .i0(\cu_ru/m_s_cause/n4 [63]),
    .i1(\cu_ru/trap_cause [63]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b7  (
    .i0(\cu_ru/m_s_cause/n4 [7]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b8  (
    .i0(\cu_ru/m_s_cause/n4 [8]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux3_b9  (
    .i0(\cu_ru/m_s_cause/n4 [9]),
    .i1(1'b0),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_cause/n5 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  AL_MUX \cu_ru/m_s_cause/mux4_b0  (
    .i0(\cu_ru/mcause [0]),
    .i1(data_csr[0]),
    .sel(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n6 [0]));
  and \cu_ru/m_s_cause/mux4_b0_sel_is_2  (\cu_ru/m_s_cause/mux4_b0_sel_is_2_o , \cu_ru/trap_target_s_neg , \cu_ru/m_s_cause/n0 );
  AL_MUX \cu_ru/m_s_cause/mux4_b1  (
    .i0(\cu_ru/mcause [1]),
    .i1(data_csr[1]),
    .sel(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n6 [1]));
  AL_MUX \cu_ru/m_s_cause/mux4_b2  (
    .i0(\cu_ru/mcause [2]),
    .i1(data_csr[2]),
    .sel(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n6 [2]));
  AL_MUX \cu_ru/m_s_cause/mux4_b3  (
    .i0(\cu_ru/mcause [3]),
    .i1(data_csr[3]),
    .sel(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n6 [3]));
  AL_MUX \cu_ru/m_s_cause/mux4_b63  (
    .i0(\cu_ru/mcause [63]),
    .i1(data_csr[63]),
    .sel(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_cause/n6 [63]));
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux5_b0  (
    .i0(\cu_ru/m_s_cause/n6 [0]),
    .i1(\cu_ru/trap_cause [0]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_cause/n7 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux5_b1  (
    .i0(\cu_ru/m_s_cause/n6 [1]),
    .i1(\cu_ru/trap_cause [1]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_cause/n7 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux5_b2  (
    .i0(\cu_ru/m_s_cause/n6 [2]),
    .i1(\cu_ru/trap_cause [2]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_cause/n7 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux5_b3  (
    .i0(\cu_ru/m_s_cause/n6 [3]),
    .i1(\cu_ru/trap_cause [3]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_cause/n7 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  binary_mux_s1_w1 \cu_ru/m_s_cause/mux5_b63  (
    .i0(\cu_ru/m_s_cause/n6 [63]),
    .i1(\cu_ru/trap_cause [63]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_cause/n7 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(35)
  and \cu_ru/m_s_cause/mux7_b10_sel_is_0  (\cu_ru/m_s_cause/mux7_b10_sel_is_0_o , rst_neg, \cu_ru/trap_target_m_neg );
  not \cu_ru/m_s_cause/n0_inv  (\cu_ru/m_s_cause/n0_neg , \cu_ru/m_s_cause/n0 );
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b0  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [0]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b1  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [1]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b10  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [10]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b11  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [11]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b12  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [12]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b13  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [13]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b14  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [14]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b15  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [15]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b16  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [16]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b17  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [17]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b18  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [18]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b19  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [19]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b2  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [2]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b20  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [20]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b21  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [21]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b22  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [22]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b23  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [23]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b24  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [24]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b25  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [25]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b26  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [26]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b27  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [27]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b28  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [28]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b29  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [29]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b3  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [3]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b30  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [30]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b31  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [31]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b32  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [32]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b33  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [33]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b34  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [34]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b35  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [35]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b36  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [36]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b37  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [37]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b38  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [38]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b39  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [39]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b4  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [4]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b40  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [40]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b41  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [41]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b42  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [42]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b43  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [43]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b44  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [44]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b45  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [45]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b46  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [46]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b47  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [47]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b48  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [48]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b49  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [49]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b5  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [5]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b50  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [50]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b51  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [51]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b52  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [52]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b53  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [53]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b54  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [54]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b55  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [55]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b56  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [56]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b57  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [57]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b58  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [58]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b59  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [59]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b6  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [6]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b60  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [60]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b61  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [61]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b62  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [62]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b63  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [63]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b7  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [7]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b8  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [8]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg0_b9  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n5 [9]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/scause [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b0  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n7 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcause [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b1  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n7 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcause [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b10  (
    .clk(clk),
    .d(data_csr[10]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b11  (
    .clk(clk),
    .d(data_csr[11]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b12  (
    .clk(clk),
    .d(data_csr[12]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b13  (
    .clk(clk),
    .d(data_csr[13]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b14  (
    .clk(clk),
    .d(data_csr[14]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b15  (
    .clk(clk),
    .d(data_csr[15]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b16  (
    .clk(clk),
    .d(data_csr[16]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b17  (
    .clk(clk),
    .d(data_csr[17]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b18  (
    .clk(clk),
    .d(data_csr[18]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b19  (
    .clk(clk),
    .d(data_csr[19]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b2  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n7 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcause [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b20  (
    .clk(clk),
    .d(data_csr[20]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b21  (
    .clk(clk),
    .d(data_csr[21]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b22  (
    .clk(clk),
    .d(data_csr[22]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b23  (
    .clk(clk),
    .d(data_csr[23]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b24  (
    .clk(clk),
    .d(data_csr[24]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b25  (
    .clk(clk),
    .d(data_csr[25]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b26  (
    .clk(clk),
    .d(data_csr[26]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b27  (
    .clk(clk),
    .d(data_csr[27]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b28  (
    .clk(clk),
    .d(data_csr[28]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b29  (
    .clk(clk),
    .d(data_csr[29]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b3  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n7 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcause [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b30  (
    .clk(clk),
    .d(data_csr[30]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b31  (
    .clk(clk),
    .d(data_csr[31]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b32  (
    .clk(clk),
    .d(data_csr[32]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b33  (
    .clk(clk),
    .d(data_csr[33]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b34  (
    .clk(clk),
    .d(data_csr[34]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b35  (
    .clk(clk),
    .d(data_csr[35]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b36  (
    .clk(clk),
    .d(data_csr[36]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b37  (
    .clk(clk),
    .d(data_csr[37]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b38  (
    .clk(clk),
    .d(data_csr[38]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b39  (
    .clk(clk),
    .d(data_csr[39]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b4  (
    .clk(clk),
    .d(data_csr[4]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b40  (
    .clk(clk),
    .d(data_csr[40]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b41  (
    .clk(clk),
    .d(data_csr[41]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b42  (
    .clk(clk),
    .d(data_csr[42]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b43  (
    .clk(clk),
    .d(data_csr[43]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b44  (
    .clk(clk),
    .d(data_csr[44]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b45  (
    .clk(clk),
    .d(data_csr[45]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b46  (
    .clk(clk),
    .d(data_csr[46]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b47  (
    .clk(clk),
    .d(data_csr[47]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b48  (
    .clk(clk),
    .d(data_csr[48]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b49  (
    .clk(clk),
    .d(data_csr[49]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b5  (
    .clk(clk),
    .d(data_csr[5]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b50  (
    .clk(clk),
    .d(data_csr[50]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b51  (
    .clk(clk),
    .d(data_csr[51]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b52  (
    .clk(clk),
    .d(data_csr[52]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b53  (
    .clk(clk),
    .d(data_csr[53]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b54  (
    .clk(clk),
    .d(data_csr[54]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b55  (
    .clk(clk),
    .d(data_csr[55]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b56  (
    .clk(clk),
    .d(data_csr[56]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b57  (
    .clk(clk),
    .d(data_csr[57]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b58  (
    .clk(clk),
    .d(data_csr[58]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b59  (
    .clk(clk),
    .d(data_csr[59]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b6  (
    .clk(clk),
    .d(data_csr[6]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b60  (
    .clk(clk),
    .d(data_csr[60]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b61  (
    .clk(clk),
    .d(data_csr[61]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b62  (
    .clk(clk),
    .d(data_csr[62]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b63  (
    .clk(clk),
    .d(\cu_ru/m_s_cause/n7 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mcause [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b7  (
    .clk(clk),
    .d(data_csr[7]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b8  (
    .clk(clk),
    .d(data_csr[8]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  reg_sr_as_w1 \cu_ru/m_s_cause/reg1_b9  (
    .clk(clk),
    .d(data_csr[9]),
    .en(\cu_ru/m_s_cause/mux4_b0_sel_is_2_o ),
    .reset(~\cu_ru/m_s_cause/mux7_b10_sel_is_0_o ),
    .set(1'b0),
    .q(\cu_ru/mcause [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(36)
  and \cu_ru/m_s_cause/u1  (\cu_ru/m_s_cause/n0 , \cu_ru/mrw_mcause_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(30)
  and \cu_ru/m_s_cause/u2  (\cu_ru/m_s_cause/n1 , \cu_ru/srw_scause_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_cause.v(33)
  add_pu62_pu62_o62 \cu_ru/m_s_epc/add0  (
    .i0(wb_ins_pc[63:2]),
    .i1(62'b00000000000000000000000000000000000000000000000000000000000001),
    .o(\cu_ru/m_s_epc/n0 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b10  (
    .i0(\cu_ru/m_s_epc/n0 [8]),
    .i1(new_pc[10]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b11  (
    .i0(\cu_ru/m_s_epc/n0 [9]),
    .i1(new_pc[11]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b12  (
    .i0(\cu_ru/m_s_epc/n0 [10]),
    .i1(new_pc[12]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b13  (
    .i0(\cu_ru/m_s_epc/n0 [11]),
    .i1(new_pc[13]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b14  (
    .i0(\cu_ru/m_s_epc/n0 [12]),
    .i1(new_pc[14]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b15  (
    .i0(\cu_ru/m_s_epc/n0 [13]),
    .i1(new_pc[15]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b16  (
    .i0(\cu_ru/m_s_epc/n0 [14]),
    .i1(new_pc[16]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b17  (
    .i0(\cu_ru/m_s_epc/n0 [15]),
    .i1(new_pc[17]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b18  (
    .i0(\cu_ru/m_s_epc/n0 [16]),
    .i1(new_pc[18]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b19  (
    .i0(\cu_ru/m_s_epc/n0 [17]),
    .i1(new_pc[19]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b2  (
    .i0(\cu_ru/m_s_epc/n0 [0]),
    .i1(new_pc[2]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b20  (
    .i0(\cu_ru/m_s_epc/n0 [18]),
    .i1(new_pc[20]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b21  (
    .i0(\cu_ru/m_s_epc/n0 [19]),
    .i1(new_pc[21]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b22  (
    .i0(\cu_ru/m_s_epc/n0 [20]),
    .i1(new_pc[22]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b23  (
    .i0(\cu_ru/m_s_epc/n0 [21]),
    .i1(new_pc[23]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b24  (
    .i0(\cu_ru/m_s_epc/n0 [22]),
    .i1(new_pc[24]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b25  (
    .i0(\cu_ru/m_s_epc/n0 [23]),
    .i1(new_pc[25]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b26  (
    .i0(\cu_ru/m_s_epc/n0 [24]),
    .i1(new_pc[26]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b27  (
    .i0(\cu_ru/m_s_epc/n0 [25]),
    .i1(new_pc[27]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b28  (
    .i0(\cu_ru/m_s_epc/n0 [26]),
    .i1(new_pc[28]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b29  (
    .i0(\cu_ru/m_s_epc/n0 [27]),
    .i1(new_pc[29]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b3  (
    .i0(\cu_ru/m_s_epc/n0 [1]),
    .i1(new_pc[3]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b30  (
    .i0(\cu_ru/m_s_epc/n0 [28]),
    .i1(new_pc[30]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b31  (
    .i0(\cu_ru/m_s_epc/n0 [29]),
    .i1(new_pc[31]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b32  (
    .i0(\cu_ru/m_s_epc/n0 [30]),
    .i1(new_pc[32]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b33  (
    .i0(\cu_ru/m_s_epc/n0 [31]),
    .i1(new_pc[33]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b34  (
    .i0(\cu_ru/m_s_epc/n0 [32]),
    .i1(new_pc[34]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b35  (
    .i0(\cu_ru/m_s_epc/n0 [33]),
    .i1(new_pc[35]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b36  (
    .i0(\cu_ru/m_s_epc/n0 [34]),
    .i1(new_pc[36]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b37  (
    .i0(\cu_ru/m_s_epc/n0 [35]),
    .i1(new_pc[37]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b38  (
    .i0(\cu_ru/m_s_epc/n0 [36]),
    .i1(new_pc[38]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b39  (
    .i0(\cu_ru/m_s_epc/n0 [37]),
    .i1(new_pc[39]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b4  (
    .i0(\cu_ru/m_s_epc/n0 [2]),
    .i1(new_pc[4]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b40  (
    .i0(\cu_ru/m_s_epc/n0 [38]),
    .i1(new_pc[40]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b41  (
    .i0(\cu_ru/m_s_epc/n0 [39]),
    .i1(new_pc[41]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b42  (
    .i0(\cu_ru/m_s_epc/n0 [40]),
    .i1(new_pc[42]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b43  (
    .i0(\cu_ru/m_s_epc/n0 [41]),
    .i1(new_pc[43]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b44  (
    .i0(\cu_ru/m_s_epc/n0 [42]),
    .i1(new_pc[44]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b45  (
    .i0(\cu_ru/m_s_epc/n0 [43]),
    .i1(new_pc[45]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b46  (
    .i0(\cu_ru/m_s_epc/n0 [44]),
    .i1(new_pc[46]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b47  (
    .i0(\cu_ru/m_s_epc/n0 [45]),
    .i1(new_pc[47]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b48  (
    .i0(\cu_ru/m_s_epc/n0 [46]),
    .i1(new_pc[48]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b49  (
    .i0(\cu_ru/m_s_epc/n0 [47]),
    .i1(new_pc[49]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b5  (
    .i0(\cu_ru/m_s_epc/n0 [3]),
    .i1(new_pc[5]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b50  (
    .i0(\cu_ru/m_s_epc/n0 [48]),
    .i1(new_pc[50]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b51  (
    .i0(\cu_ru/m_s_epc/n0 [49]),
    .i1(new_pc[51]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b52  (
    .i0(\cu_ru/m_s_epc/n0 [50]),
    .i1(new_pc[52]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b53  (
    .i0(\cu_ru/m_s_epc/n0 [51]),
    .i1(new_pc[53]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b54  (
    .i0(\cu_ru/m_s_epc/n0 [52]),
    .i1(new_pc[54]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b55  (
    .i0(\cu_ru/m_s_epc/n0 [53]),
    .i1(new_pc[55]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b56  (
    .i0(\cu_ru/m_s_epc/n0 [54]),
    .i1(new_pc[56]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b57  (
    .i0(\cu_ru/m_s_epc/n0 [55]),
    .i1(new_pc[57]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b58  (
    .i0(\cu_ru/m_s_epc/n0 [56]),
    .i1(new_pc[58]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b59  (
    .i0(\cu_ru/m_s_epc/n0 [57]),
    .i1(new_pc[59]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b6  (
    .i0(\cu_ru/m_s_epc/n0 [4]),
    .i1(new_pc[6]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b60  (
    .i0(\cu_ru/m_s_epc/n0 [58]),
    .i1(new_pc[60]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b61  (
    .i0(\cu_ru/m_s_epc/n0 [59]),
    .i1(new_pc[61]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b62  (
    .i0(\cu_ru/m_s_epc/n0 [60]),
    .i1(new_pc[62]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b63  (
    .i0(\cu_ru/m_s_epc/n0 [61]),
    .i1(new_pc[63]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b7  (
    .i0(\cu_ru/m_s_epc/n0 [5]),
    .i1(new_pc[7]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b8  (
    .i0(\cu_ru/m_s_epc/n0 [6]),
    .i1(new_pc[8]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux0_b9  (
    .i0(\cu_ru/m_s_epc/n0 [7]),
    .i1(new_pc[9]),
    .sel(pc_jmp),
    .o(\cu_ru/m_s_epc/n1 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  AL_MUX \cu_ru/m_s_epc/mux1_b0  (
    .i0(wb_ins_pc[0]),
    .i1(new_pc[0]),
    .sel(\cu_ru/m_s_epc/mux1_b0_sel_is_3_o ),
    .o(\cu_ru/m_s_epc/n2 [0]));
  and \cu_ru/m_s_epc/mux1_b0_sel_is_3  (\cu_ru/m_s_epc/mux1_b0_sel_is_3_o , \cu_ru/next_pc , pc_jmp);
  AL_MUX \cu_ru/m_s_epc/mux1_b1  (
    .i0(wb_ins_pc[1]),
    .i1(new_pc[1]),
    .sel(\cu_ru/m_s_epc/mux1_b0_sel_is_3_o ),
    .o(\cu_ru/m_s_epc/n2 [1]));
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b10  (
    .i0(wb_ins_pc[10]),
    .i1(\cu_ru/m_s_epc/n1 [10]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b11  (
    .i0(wb_ins_pc[11]),
    .i1(\cu_ru/m_s_epc/n1 [11]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b12  (
    .i0(wb_ins_pc[12]),
    .i1(\cu_ru/m_s_epc/n1 [12]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b13  (
    .i0(wb_ins_pc[13]),
    .i1(\cu_ru/m_s_epc/n1 [13]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b14  (
    .i0(wb_ins_pc[14]),
    .i1(\cu_ru/m_s_epc/n1 [14]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b15  (
    .i0(wb_ins_pc[15]),
    .i1(\cu_ru/m_s_epc/n1 [15]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b16  (
    .i0(wb_ins_pc[16]),
    .i1(\cu_ru/m_s_epc/n1 [16]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b17  (
    .i0(wb_ins_pc[17]),
    .i1(\cu_ru/m_s_epc/n1 [17]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b18  (
    .i0(wb_ins_pc[18]),
    .i1(\cu_ru/m_s_epc/n1 [18]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b19  (
    .i0(wb_ins_pc[19]),
    .i1(\cu_ru/m_s_epc/n1 [19]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b2  (
    .i0(wb_ins_pc[2]),
    .i1(\cu_ru/m_s_epc/n1 [2]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b20  (
    .i0(wb_ins_pc[20]),
    .i1(\cu_ru/m_s_epc/n1 [20]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b21  (
    .i0(wb_ins_pc[21]),
    .i1(\cu_ru/m_s_epc/n1 [21]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b22  (
    .i0(wb_ins_pc[22]),
    .i1(\cu_ru/m_s_epc/n1 [22]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b23  (
    .i0(wb_ins_pc[23]),
    .i1(\cu_ru/m_s_epc/n1 [23]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b24  (
    .i0(wb_ins_pc[24]),
    .i1(\cu_ru/m_s_epc/n1 [24]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b25  (
    .i0(wb_ins_pc[25]),
    .i1(\cu_ru/m_s_epc/n1 [25]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b26  (
    .i0(wb_ins_pc[26]),
    .i1(\cu_ru/m_s_epc/n1 [26]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b27  (
    .i0(wb_ins_pc[27]),
    .i1(\cu_ru/m_s_epc/n1 [27]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b28  (
    .i0(wb_ins_pc[28]),
    .i1(\cu_ru/m_s_epc/n1 [28]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b29  (
    .i0(wb_ins_pc[29]),
    .i1(\cu_ru/m_s_epc/n1 [29]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b3  (
    .i0(wb_ins_pc[3]),
    .i1(\cu_ru/m_s_epc/n1 [3]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b30  (
    .i0(wb_ins_pc[30]),
    .i1(\cu_ru/m_s_epc/n1 [30]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b31  (
    .i0(wb_ins_pc[31]),
    .i1(\cu_ru/m_s_epc/n1 [31]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b32  (
    .i0(wb_ins_pc[32]),
    .i1(\cu_ru/m_s_epc/n1 [32]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b33  (
    .i0(wb_ins_pc[33]),
    .i1(\cu_ru/m_s_epc/n1 [33]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b34  (
    .i0(wb_ins_pc[34]),
    .i1(\cu_ru/m_s_epc/n1 [34]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b35  (
    .i0(wb_ins_pc[35]),
    .i1(\cu_ru/m_s_epc/n1 [35]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b36  (
    .i0(wb_ins_pc[36]),
    .i1(\cu_ru/m_s_epc/n1 [36]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b37  (
    .i0(wb_ins_pc[37]),
    .i1(\cu_ru/m_s_epc/n1 [37]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b38  (
    .i0(wb_ins_pc[38]),
    .i1(\cu_ru/m_s_epc/n1 [38]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b39  (
    .i0(wb_ins_pc[39]),
    .i1(\cu_ru/m_s_epc/n1 [39]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b4  (
    .i0(wb_ins_pc[4]),
    .i1(\cu_ru/m_s_epc/n1 [4]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b40  (
    .i0(wb_ins_pc[40]),
    .i1(\cu_ru/m_s_epc/n1 [40]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b41  (
    .i0(wb_ins_pc[41]),
    .i1(\cu_ru/m_s_epc/n1 [41]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b42  (
    .i0(wb_ins_pc[42]),
    .i1(\cu_ru/m_s_epc/n1 [42]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b43  (
    .i0(wb_ins_pc[43]),
    .i1(\cu_ru/m_s_epc/n1 [43]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b44  (
    .i0(wb_ins_pc[44]),
    .i1(\cu_ru/m_s_epc/n1 [44]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b45  (
    .i0(wb_ins_pc[45]),
    .i1(\cu_ru/m_s_epc/n1 [45]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b46  (
    .i0(wb_ins_pc[46]),
    .i1(\cu_ru/m_s_epc/n1 [46]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b47  (
    .i0(wb_ins_pc[47]),
    .i1(\cu_ru/m_s_epc/n1 [47]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b48  (
    .i0(wb_ins_pc[48]),
    .i1(\cu_ru/m_s_epc/n1 [48]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b49  (
    .i0(wb_ins_pc[49]),
    .i1(\cu_ru/m_s_epc/n1 [49]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b5  (
    .i0(wb_ins_pc[5]),
    .i1(\cu_ru/m_s_epc/n1 [5]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b50  (
    .i0(wb_ins_pc[50]),
    .i1(\cu_ru/m_s_epc/n1 [50]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b51  (
    .i0(wb_ins_pc[51]),
    .i1(\cu_ru/m_s_epc/n1 [51]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b52  (
    .i0(wb_ins_pc[52]),
    .i1(\cu_ru/m_s_epc/n1 [52]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b53  (
    .i0(wb_ins_pc[53]),
    .i1(\cu_ru/m_s_epc/n1 [53]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b54  (
    .i0(wb_ins_pc[54]),
    .i1(\cu_ru/m_s_epc/n1 [54]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b55  (
    .i0(wb_ins_pc[55]),
    .i1(\cu_ru/m_s_epc/n1 [55]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b56  (
    .i0(wb_ins_pc[56]),
    .i1(\cu_ru/m_s_epc/n1 [56]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b57  (
    .i0(wb_ins_pc[57]),
    .i1(\cu_ru/m_s_epc/n1 [57]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b58  (
    .i0(wb_ins_pc[58]),
    .i1(\cu_ru/m_s_epc/n1 [58]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b59  (
    .i0(wb_ins_pc[59]),
    .i1(\cu_ru/m_s_epc/n1 [59]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b6  (
    .i0(wb_ins_pc[6]),
    .i1(\cu_ru/m_s_epc/n1 [6]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b60  (
    .i0(wb_ins_pc[60]),
    .i1(\cu_ru/m_s_epc/n1 [60]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b61  (
    .i0(wb_ins_pc[61]),
    .i1(\cu_ru/m_s_epc/n1 [61]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b62  (
    .i0(wb_ins_pc[62]),
    .i1(\cu_ru/m_s_epc/n1 [62]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b63  (
    .i0(wb_ins_pc[63]),
    .i1(\cu_ru/m_s_epc/n1 [63]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b7  (
    .i0(wb_ins_pc[7]),
    .i1(\cu_ru/m_s_epc/n1 [7]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b8  (
    .i0(wb_ins_pc[8]),
    .i1(\cu_ru/m_s_epc/n1 [8]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux1_b9  (
    .i0(wb_ins_pc[9]),
    .i1(\cu_ru/m_s_epc/n1 [9]),
    .sel(\cu_ru/next_pc ),
    .o(\cu_ru/m_s_epc/n2 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(30)
  AL_MUX \cu_ru/m_s_epc/mux4_b0  (
    .i0(\cu_ru/sepc [0]),
    .i1(data_csr[0]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [0]));
  and \cu_ru/m_s_epc/mux4_b0_sel_is_2  (\cu_ru/m_s_epc/mux4_b0_sel_is_2_o , \cu_ru/m_s_epc/n3_neg , \cu_ru/m_s_epc/n4 );
  AL_MUX \cu_ru/m_s_epc/mux4_b1  (
    .i0(\cu_ru/sepc [1]),
    .i1(data_csr[1]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [1]));
  AL_MUX \cu_ru/m_s_epc/mux4_b10  (
    .i0(\cu_ru/sepc [10]),
    .i1(data_csr[10]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [10]));
  AL_MUX \cu_ru/m_s_epc/mux4_b11  (
    .i0(\cu_ru/sepc [11]),
    .i1(data_csr[11]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [11]));
  AL_MUX \cu_ru/m_s_epc/mux4_b12  (
    .i0(\cu_ru/sepc [12]),
    .i1(data_csr[12]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [12]));
  AL_MUX \cu_ru/m_s_epc/mux4_b13  (
    .i0(\cu_ru/sepc [13]),
    .i1(data_csr[13]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [13]));
  AL_MUX \cu_ru/m_s_epc/mux4_b14  (
    .i0(\cu_ru/sepc [14]),
    .i1(data_csr[14]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [14]));
  AL_MUX \cu_ru/m_s_epc/mux4_b15  (
    .i0(\cu_ru/sepc [15]),
    .i1(data_csr[15]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [15]));
  AL_MUX \cu_ru/m_s_epc/mux4_b16  (
    .i0(\cu_ru/sepc [16]),
    .i1(data_csr[16]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [16]));
  AL_MUX \cu_ru/m_s_epc/mux4_b17  (
    .i0(\cu_ru/sepc [17]),
    .i1(data_csr[17]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [17]));
  AL_MUX \cu_ru/m_s_epc/mux4_b18  (
    .i0(\cu_ru/sepc [18]),
    .i1(data_csr[18]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [18]));
  AL_MUX \cu_ru/m_s_epc/mux4_b19  (
    .i0(\cu_ru/sepc [19]),
    .i1(data_csr[19]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [19]));
  AL_MUX \cu_ru/m_s_epc/mux4_b2  (
    .i0(\cu_ru/sepc [2]),
    .i1(data_csr[2]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [2]));
  AL_MUX \cu_ru/m_s_epc/mux4_b20  (
    .i0(\cu_ru/sepc [20]),
    .i1(data_csr[20]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [20]));
  AL_MUX \cu_ru/m_s_epc/mux4_b21  (
    .i0(\cu_ru/sepc [21]),
    .i1(data_csr[21]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [21]));
  AL_MUX \cu_ru/m_s_epc/mux4_b22  (
    .i0(\cu_ru/sepc [22]),
    .i1(data_csr[22]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [22]));
  AL_MUX \cu_ru/m_s_epc/mux4_b23  (
    .i0(\cu_ru/sepc [23]),
    .i1(data_csr[23]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [23]));
  AL_MUX \cu_ru/m_s_epc/mux4_b24  (
    .i0(\cu_ru/sepc [24]),
    .i1(data_csr[24]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [24]));
  AL_MUX \cu_ru/m_s_epc/mux4_b25  (
    .i0(\cu_ru/sepc [25]),
    .i1(data_csr[25]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [25]));
  AL_MUX \cu_ru/m_s_epc/mux4_b26  (
    .i0(\cu_ru/sepc [26]),
    .i1(data_csr[26]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [26]));
  AL_MUX \cu_ru/m_s_epc/mux4_b27  (
    .i0(\cu_ru/sepc [27]),
    .i1(data_csr[27]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [27]));
  AL_MUX \cu_ru/m_s_epc/mux4_b28  (
    .i0(\cu_ru/sepc [28]),
    .i1(data_csr[28]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [28]));
  AL_MUX \cu_ru/m_s_epc/mux4_b29  (
    .i0(\cu_ru/sepc [29]),
    .i1(data_csr[29]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [29]));
  AL_MUX \cu_ru/m_s_epc/mux4_b3  (
    .i0(\cu_ru/sepc [3]),
    .i1(data_csr[3]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [3]));
  AL_MUX \cu_ru/m_s_epc/mux4_b30  (
    .i0(\cu_ru/sepc [30]),
    .i1(data_csr[30]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [30]));
  AL_MUX \cu_ru/m_s_epc/mux4_b31  (
    .i0(\cu_ru/sepc [31]),
    .i1(data_csr[31]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [31]));
  AL_MUX \cu_ru/m_s_epc/mux4_b32  (
    .i0(\cu_ru/sepc [32]),
    .i1(data_csr[32]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [32]));
  AL_MUX \cu_ru/m_s_epc/mux4_b33  (
    .i0(\cu_ru/sepc [33]),
    .i1(data_csr[33]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [33]));
  AL_MUX \cu_ru/m_s_epc/mux4_b34  (
    .i0(\cu_ru/sepc [34]),
    .i1(data_csr[34]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [34]));
  AL_MUX \cu_ru/m_s_epc/mux4_b35  (
    .i0(\cu_ru/sepc [35]),
    .i1(data_csr[35]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [35]));
  AL_MUX \cu_ru/m_s_epc/mux4_b36  (
    .i0(\cu_ru/sepc [36]),
    .i1(data_csr[36]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [36]));
  AL_MUX \cu_ru/m_s_epc/mux4_b37  (
    .i0(\cu_ru/sepc [37]),
    .i1(data_csr[37]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [37]));
  AL_MUX \cu_ru/m_s_epc/mux4_b38  (
    .i0(\cu_ru/sepc [38]),
    .i1(data_csr[38]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [38]));
  AL_MUX \cu_ru/m_s_epc/mux4_b39  (
    .i0(\cu_ru/sepc [39]),
    .i1(data_csr[39]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [39]));
  AL_MUX \cu_ru/m_s_epc/mux4_b4  (
    .i0(\cu_ru/sepc [4]),
    .i1(data_csr[4]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [4]));
  AL_MUX \cu_ru/m_s_epc/mux4_b40  (
    .i0(\cu_ru/sepc [40]),
    .i1(data_csr[40]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [40]));
  AL_MUX \cu_ru/m_s_epc/mux4_b41  (
    .i0(\cu_ru/sepc [41]),
    .i1(data_csr[41]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [41]));
  AL_MUX \cu_ru/m_s_epc/mux4_b42  (
    .i0(\cu_ru/sepc [42]),
    .i1(data_csr[42]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [42]));
  AL_MUX \cu_ru/m_s_epc/mux4_b43  (
    .i0(\cu_ru/sepc [43]),
    .i1(data_csr[43]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [43]));
  AL_MUX \cu_ru/m_s_epc/mux4_b44  (
    .i0(\cu_ru/sepc [44]),
    .i1(data_csr[44]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [44]));
  AL_MUX \cu_ru/m_s_epc/mux4_b45  (
    .i0(\cu_ru/sepc [45]),
    .i1(data_csr[45]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [45]));
  AL_MUX \cu_ru/m_s_epc/mux4_b46  (
    .i0(\cu_ru/sepc [46]),
    .i1(data_csr[46]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [46]));
  AL_MUX \cu_ru/m_s_epc/mux4_b47  (
    .i0(\cu_ru/sepc [47]),
    .i1(data_csr[47]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [47]));
  AL_MUX \cu_ru/m_s_epc/mux4_b48  (
    .i0(\cu_ru/sepc [48]),
    .i1(data_csr[48]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [48]));
  AL_MUX \cu_ru/m_s_epc/mux4_b49  (
    .i0(\cu_ru/sepc [49]),
    .i1(data_csr[49]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [49]));
  AL_MUX \cu_ru/m_s_epc/mux4_b5  (
    .i0(\cu_ru/sepc [5]),
    .i1(data_csr[5]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [5]));
  AL_MUX \cu_ru/m_s_epc/mux4_b50  (
    .i0(\cu_ru/sepc [50]),
    .i1(data_csr[50]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [50]));
  AL_MUX \cu_ru/m_s_epc/mux4_b51  (
    .i0(\cu_ru/sepc [51]),
    .i1(data_csr[51]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [51]));
  AL_MUX \cu_ru/m_s_epc/mux4_b52  (
    .i0(\cu_ru/sepc [52]),
    .i1(data_csr[52]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [52]));
  AL_MUX \cu_ru/m_s_epc/mux4_b53  (
    .i0(\cu_ru/sepc [53]),
    .i1(data_csr[53]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [53]));
  AL_MUX \cu_ru/m_s_epc/mux4_b54  (
    .i0(\cu_ru/sepc [54]),
    .i1(data_csr[54]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [54]));
  AL_MUX \cu_ru/m_s_epc/mux4_b55  (
    .i0(\cu_ru/sepc [55]),
    .i1(data_csr[55]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [55]));
  AL_MUX \cu_ru/m_s_epc/mux4_b56  (
    .i0(\cu_ru/sepc [56]),
    .i1(data_csr[56]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [56]));
  AL_MUX \cu_ru/m_s_epc/mux4_b57  (
    .i0(\cu_ru/sepc [57]),
    .i1(data_csr[57]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [57]));
  AL_MUX \cu_ru/m_s_epc/mux4_b58  (
    .i0(\cu_ru/sepc [58]),
    .i1(data_csr[58]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [58]));
  AL_MUX \cu_ru/m_s_epc/mux4_b59  (
    .i0(\cu_ru/sepc [59]),
    .i1(data_csr[59]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [59]));
  AL_MUX \cu_ru/m_s_epc/mux4_b6  (
    .i0(\cu_ru/sepc [6]),
    .i1(data_csr[6]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [6]));
  AL_MUX \cu_ru/m_s_epc/mux4_b60  (
    .i0(\cu_ru/sepc [60]),
    .i1(data_csr[60]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [60]));
  AL_MUX \cu_ru/m_s_epc/mux4_b61  (
    .i0(\cu_ru/sepc [61]),
    .i1(data_csr[61]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [61]));
  AL_MUX \cu_ru/m_s_epc/mux4_b62  (
    .i0(\cu_ru/sepc [62]),
    .i1(data_csr[62]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [62]));
  AL_MUX \cu_ru/m_s_epc/mux4_b63  (
    .i0(\cu_ru/sepc [63]),
    .i1(data_csr[63]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [63]));
  AL_MUX \cu_ru/m_s_epc/mux4_b7  (
    .i0(\cu_ru/sepc [7]),
    .i1(data_csr[7]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [7]));
  AL_MUX \cu_ru/m_s_epc/mux4_b8  (
    .i0(\cu_ru/sepc [8]),
    .i1(data_csr[8]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [8]));
  AL_MUX \cu_ru/m_s_epc/mux4_b9  (
    .i0(\cu_ru/sepc [9]),
    .i1(data_csr[9]),
    .sel(\cu_ru/m_s_epc/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n7 [9]));
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b0  (
    .i0(\cu_ru/m_s_epc/n7 [0]),
    .i1(\cu_ru/m_s_epc/n2 [0]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b1  (
    .i0(\cu_ru/m_s_epc/n7 [1]),
    .i1(\cu_ru/m_s_epc/n2 [1]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b10  (
    .i0(\cu_ru/m_s_epc/n7 [10]),
    .i1(\cu_ru/m_s_epc/n2 [10]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b11  (
    .i0(\cu_ru/m_s_epc/n7 [11]),
    .i1(\cu_ru/m_s_epc/n2 [11]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b12  (
    .i0(\cu_ru/m_s_epc/n7 [12]),
    .i1(\cu_ru/m_s_epc/n2 [12]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b13  (
    .i0(\cu_ru/m_s_epc/n7 [13]),
    .i1(\cu_ru/m_s_epc/n2 [13]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b14  (
    .i0(\cu_ru/m_s_epc/n7 [14]),
    .i1(\cu_ru/m_s_epc/n2 [14]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b15  (
    .i0(\cu_ru/m_s_epc/n7 [15]),
    .i1(\cu_ru/m_s_epc/n2 [15]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b16  (
    .i0(\cu_ru/m_s_epc/n7 [16]),
    .i1(\cu_ru/m_s_epc/n2 [16]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b17  (
    .i0(\cu_ru/m_s_epc/n7 [17]),
    .i1(\cu_ru/m_s_epc/n2 [17]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b18  (
    .i0(\cu_ru/m_s_epc/n7 [18]),
    .i1(\cu_ru/m_s_epc/n2 [18]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b19  (
    .i0(\cu_ru/m_s_epc/n7 [19]),
    .i1(\cu_ru/m_s_epc/n2 [19]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b2  (
    .i0(\cu_ru/m_s_epc/n7 [2]),
    .i1(\cu_ru/m_s_epc/n2 [2]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b20  (
    .i0(\cu_ru/m_s_epc/n7 [20]),
    .i1(\cu_ru/m_s_epc/n2 [20]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b21  (
    .i0(\cu_ru/m_s_epc/n7 [21]),
    .i1(\cu_ru/m_s_epc/n2 [21]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b22  (
    .i0(\cu_ru/m_s_epc/n7 [22]),
    .i1(\cu_ru/m_s_epc/n2 [22]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b23  (
    .i0(\cu_ru/m_s_epc/n7 [23]),
    .i1(\cu_ru/m_s_epc/n2 [23]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b24  (
    .i0(\cu_ru/m_s_epc/n7 [24]),
    .i1(\cu_ru/m_s_epc/n2 [24]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b25  (
    .i0(\cu_ru/m_s_epc/n7 [25]),
    .i1(\cu_ru/m_s_epc/n2 [25]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b26  (
    .i0(\cu_ru/m_s_epc/n7 [26]),
    .i1(\cu_ru/m_s_epc/n2 [26]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b27  (
    .i0(\cu_ru/m_s_epc/n7 [27]),
    .i1(\cu_ru/m_s_epc/n2 [27]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b28  (
    .i0(\cu_ru/m_s_epc/n7 [28]),
    .i1(\cu_ru/m_s_epc/n2 [28]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b29  (
    .i0(\cu_ru/m_s_epc/n7 [29]),
    .i1(\cu_ru/m_s_epc/n2 [29]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b3  (
    .i0(\cu_ru/m_s_epc/n7 [3]),
    .i1(\cu_ru/m_s_epc/n2 [3]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b30  (
    .i0(\cu_ru/m_s_epc/n7 [30]),
    .i1(\cu_ru/m_s_epc/n2 [30]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b31  (
    .i0(\cu_ru/m_s_epc/n7 [31]),
    .i1(\cu_ru/m_s_epc/n2 [31]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b32  (
    .i0(\cu_ru/m_s_epc/n7 [32]),
    .i1(\cu_ru/m_s_epc/n2 [32]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b33  (
    .i0(\cu_ru/m_s_epc/n7 [33]),
    .i1(\cu_ru/m_s_epc/n2 [33]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b34  (
    .i0(\cu_ru/m_s_epc/n7 [34]),
    .i1(\cu_ru/m_s_epc/n2 [34]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b35  (
    .i0(\cu_ru/m_s_epc/n7 [35]),
    .i1(\cu_ru/m_s_epc/n2 [35]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b36  (
    .i0(\cu_ru/m_s_epc/n7 [36]),
    .i1(\cu_ru/m_s_epc/n2 [36]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b37  (
    .i0(\cu_ru/m_s_epc/n7 [37]),
    .i1(\cu_ru/m_s_epc/n2 [37]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b38  (
    .i0(\cu_ru/m_s_epc/n7 [38]),
    .i1(\cu_ru/m_s_epc/n2 [38]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b39  (
    .i0(\cu_ru/m_s_epc/n7 [39]),
    .i1(\cu_ru/m_s_epc/n2 [39]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b4  (
    .i0(\cu_ru/m_s_epc/n7 [4]),
    .i1(\cu_ru/m_s_epc/n2 [4]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b40  (
    .i0(\cu_ru/m_s_epc/n7 [40]),
    .i1(\cu_ru/m_s_epc/n2 [40]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b41  (
    .i0(\cu_ru/m_s_epc/n7 [41]),
    .i1(\cu_ru/m_s_epc/n2 [41]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b42  (
    .i0(\cu_ru/m_s_epc/n7 [42]),
    .i1(\cu_ru/m_s_epc/n2 [42]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b43  (
    .i0(\cu_ru/m_s_epc/n7 [43]),
    .i1(\cu_ru/m_s_epc/n2 [43]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b44  (
    .i0(\cu_ru/m_s_epc/n7 [44]),
    .i1(\cu_ru/m_s_epc/n2 [44]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b45  (
    .i0(\cu_ru/m_s_epc/n7 [45]),
    .i1(\cu_ru/m_s_epc/n2 [45]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b46  (
    .i0(\cu_ru/m_s_epc/n7 [46]),
    .i1(\cu_ru/m_s_epc/n2 [46]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b47  (
    .i0(\cu_ru/m_s_epc/n7 [47]),
    .i1(\cu_ru/m_s_epc/n2 [47]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b48  (
    .i0(\cu_ru/m_s_epc/n7 [48]),
    .i1(\cu_ru/m_s_epc/n2 [48]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b49  (
    .i0(\cu_ru/m_s_epc/n7 [49]),
    .i1(\cu_ru/m_s_epc/n2 [49]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b5  (
    .i0(\cu_ru/m_s_epc/n7 [5]),
    .i1(\cu_ru/m_s_epc/n2 [5]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b50  (
    .i0(\cu_ru/m_s_epc/n7 [50]),
    .i1(\cu_ru/m_s_epc/n2 [50]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b51  (
    .i0(\cu_ru/m_s_epc/n7 [51]),
    .i1(\cu_ru/m_s_epc/n2 [51]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b52  (
    .i0(\cu_ru/m_s_epc/n7 [52]),
    .i1(\cu_ru/m_s_epc/n2 [52]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b53  (
    .i0(\cu_ru/m_s_epc/n7 [53]),
    .i1(\cu_ru/m_s_epc/n2 [53]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b54  (
    .i0(\cu_ru/m_s_epc/n7 [54]),
    .i1(\cu_ru/m_s_epc/n2 [54]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b55  (
    .i0(\cu_ru/m_s_epc/n7 [55]),
    .i1(\cu_ru/m_s_epc/n2 [55]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b56  (
    .i0(\cu_ru/m_s_epc/n7 [56]),
    .i1(\cu_ru/m_s_epc/n2 [56]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b57  (
    .i0(\cu_ru/m_s_epc/n7 [57]),
    .i1(\cu_ru/m_s_epc/n2 [57]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b58  (
    .i0(\cu_ru/m_s_epc/n7 [58]),
    .i1(\cu_ru/m_s_epc/n2 [58]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b59  (
    .i0(\cu_ru/m_s_epc/n7 [59]),
    .i1(\cu_ru/m_s_epc/n2 [59]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b6  (
    .i0(\cu_ru/m_s_epc/n7 [6]),
    .i1(\cu_ru/m_s_epc/n2 [6]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b60  (
    .i0(\cu_ru/m_s_epc/n7 [60]),
    .i1(\cu_ru/m_s_epc/n2 [60]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b61  (
    .i0(\cu_ru/m_s_epc/n7 [61]),
    .i1(\cu_ru/m_s_epc/n2 [61]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b62  (
    .i0(\cu_ru/m_s_epc/n7 [62]),
    .i1(\cu_ru/m_s_epc/n2 [62]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b63  (
    .i0(\cu_ru/m_s_epc/n7 [63]),
    .i1(\cu_ru/m_s_epc/n2 [63]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b7  (
    .i0(\cu_ru/m_s_epc/n7 [7]),
    .i1(\cu_ru/m_s_epc/n2 [7]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b8  (
    .i0(\cu_ru/m_s_epc/n7 [8]),
    .i1(\cu_ru/m_s_epc/n2 [8]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux5_b9  (
    .i0(\cu_ru/m_s_epc/n7 [9]),
    .i1(\cu_ru/m_s_epc/n2 [9]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_epc/n8 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  AL_MUX \cu_ru/m_s_epc/mux6_b0  (
    .i0(\cu_ru/mepc [0]),
    .i1(data_csr[0]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [0]));
  and \cu_ru/m_s_epc/mux6_b0_sel_is_2  (\cu_ru/m_s_epc/mux6_b0_sel_is_2_o , \cu_ru/trap_target_s_neg , \cu_ru/m_s_epc/n3 );
  AL_MUX \cu_ru/m_s_epc/mux6_b1  (
    .i0(\cu_ru/mepc [1]),
    .i1(data_csr[1]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [1]));
  AL_MUX \cu_ru/m_s_epc/mux6_b10  (
    .i0(\cu_ru/mepc [10]),
    .i1(data_csr[10]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [10]));
  AL_MUX \cu_ru/m_s_epc/mux6_b11  (
    .i0(\cu_ru/mepc [11]),
    .i1(data_csr[11]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [11]));
  AL_MUX \cu_ru/m_s_epc/mux6_b12  (
    .i0(\cu_ru/mepc [12]),
    .i1(data_csr[12]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [12]));
  AL_MUX \cu_ru/m_s_epc/mux6_b13  (
    .i0(\cu_ru/mepc [13]),
    .i1(data_csr[13]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [13]));
  AL_MUX \cu_ru/m_s_epc/mux6_b14  (
    .i0(\cu_ru/mepc [14]),
    .i1(data_csr[14]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [14]));
  AL_MUX \cu_ru/m_s_epc/mux6_b15  (
    .i0(\cu_ru/mepc [15]),
    .i1(data_csr[15]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [15]));
  AL_MUX \cu_ru/m_s_epc/mux6_b16  (
    .i0(\cu_ru/mepc [16]),
    .i1(data_csr[16]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [16]));
  AL_MUX \cu_ru/m_s_epc/mux6_b17  (
    .i0(\cu_ru/mepc [17]),
    .i1(data_csr[17]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [17]));
  AL_MUX \cu_ru/m_s_epc/mux6_b18  (
    .i0(\cu_ru/mepc [18]),
    .i1(data_csr[18]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [18]));
  AL_MUX \cu_ru/m_s_epc/mux6_b19  (
    .i0(\cu_ru/mepc [19]),
    .i1(data_csr[19]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [19]));
  AL_MUX \cu_ru/m_s_epc/mux6_b2  (
    .i0(\cu_ru/mepc [2]),
    .i1(data_csr[2]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [2]));
  AL_MUX \cu_ru/m_s_epc/mux6_b20  (
    .i0(\cu_ru/mepc [20]),
    .i1(data_csr[20]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [20]));
  AL_MUX \cu_ru/m_s_epc/mux6_b21  (
    .i0(\cu_ru/mepc [21]),
    .i1(data_csr[21]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [21]));
  AL_MUX \cu_ru/m_s_epc/mux6_b22  (
    .i0(\cu_ru/mepc [22]),
    .i1(data_csr[22]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [22]));
  AL_MUX \cu_ru/m_s_epc/mux6_b23  (
    .i0(\cu_ru/mepc [23]),
    .i1(data_csr[23]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [23]));
  AL_MUX \cu_ru/m_s_epc/mux6_b24  (
    .i0(\cu_ru/mepc [24]),
    .i1(data_csr[24]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [24]));
  AL_MUX \cu_ru/m_s_epc/mux6_b25  (
    .i0(\cu_ru/mepc [25]),
    .i1(data_csr[25]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [25]));
  AL_MUX \cu_ru/m_s_epc/mux6_b26  (
    .i0(\cu_ru/mepc [26]),
    .i1(data_csr[26]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [26]));
  AL_MUX \cu_ru/m_s_epc/mux6_b27  (
    .i0(\cu_ru/mepc [27]),
    .i1(data_csr[27]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [27]));
  AL_MUX \cu_ru/m_s_epc/mux6_b28  (
    .i0(\cu_ru/mepc [28]),
    .i1(data_csr[28]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [28]));
  AL_MUX \cu_ru/m_s_epc/mux6_b29  (
    .i0(\cu_ru/mepc [29]),
    .i1(data_csr[29]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [29]));
  AL_MUX \cu_ru/m_s_epc/mux6_b3  (
    .i0(\cu_ru/mepc [3]),
    .i1(data_csr[3]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [3]));
  AL_MUX \cu_ru/m_s_epc/mux6_b30  (
    .i0(\cu_ru/mepc [30]),
    .i1(data_csr[30]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [30]));
  AL_MUX \cu_ru/m_s_epc/mux6_b31  (
    .i0(\cu_ru/mepc [31]),
    .i1(data_csr[31]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [31]));
  AL_MUX \cu_ru/m_s_epc/mux6_b32  (
    .i0(\cu_ru/mepc [32]),
    .i1(data_csr[32]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [32]));
  AL_MUX \cu_ru/m_s_epc/mux6_b33  (
    .i0(\cu_ru/mepc [33]),
    .i1(data_csr[33]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [33]));
  AL_MUX \cu_ru/m_s_epc/mux6_b34  (
    .i0(\cu_ru/mepc [34]),
    .i1(data_csr[34]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [34]));
  AL_MUX \cu_ru/m_s_epc/mux6_b35  (
    .i0(\cu_ru/mepc [35]),
    .i1(data_csr[35]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [35]));
  AL_MUX \cu_ru/m_s_epc/mux6_b36  (
    .i0(\cu_ru/mepc [36]),
    .i1(data_csr[36]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [36]));
  AL_MUX \cu_ru/m_s_epc/mux6_b37  (
    .i0(\cu_ru/mepc [37]),
    .i1(data_csr[37]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [37]));
  AL_MUX \cu_ru/m_s_epc/mux6_b38  (
    .i0(\cu_ru/mepc [38]),
    .i1(data_csr[38]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [38]));
  AL_MUX \cu_ru/m_s_epc/mux6_b39  (
    .i0(\cu_ru/mepc [39]),
    .i1(data_csr[39]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [39]));
  AL_MUX \cu_ru/m_s_epc/mux6_b4  (
    .i0(\cu_ru/mepc [4]),
    .i1(data_csr[4]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [4]));
  AL_MUX \cu_ru/m_s_epc/mux6_b40  (
    .i0(\cu_ru/mepc [40]),
    .i1(data_csr[40]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [40]));
  AL_MUX \cu_ru/m_s_epc/mux6_b41  (
    .i0(\cu_ru/mepc [41]),
    .i1(data_csr[41]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [41]));
  AL_MUX \cu_ru/m_s_epc/mux6_b42  (
    .i0(\cu_ru/mepc [42]),
    .i1(data_csr[42]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [42]));
  AL_MUX \cu_ru/m_s_epc/mux6_b43  (
    .i0(\cu_ru/mepc [43]),
    .i1(data_csr[43]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [43]));
  AL_MUX \cu_ru/m_s_epc/mux6_b44  (
    .i0(\cu_ru/mepc [44]),
    .i1(data_csr[44]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [44]));
  AL_MUX \cu_ru/m_s_epc/mux6_b45  (
    .i0(\cu_ru/mepc [45]),
    .i1(data_csr[45]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [45]));
  AL_MUX \cu_ru/m_s_epc/mux6_b46  (
    .i0(\cu_ru/mepc [46]),
    .i1(data_csr[46]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [46]));
  AL_MUX \cu_ru/m_s_epc/mux6_b47  (
    .i0(\cu_ru/mepc [47]),
    .i1(data_csr[47]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [47]));
  AL_MUX \cu_ru/m_s_epc/mux6_b48  (
    .i0(\cu_ru/mepc [48]),
    .i1(data_csr[48]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [48]));
  AL_MUX \cu_ru/m_s_epc/mux6_b49  (
    .i0(\cu_ru/mepc [49]),
    .i1(data_csr[49]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [49]));
  AL_MUX \cu_ru/m_s_epc/mux6_b5  (
    .i0(\cu_ru/mepc [5]),
    .i1(data_csr[5]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [5]));
  AL_MUX \cu_ru/m_s_epc/mux6_b50  (
    .i0(\cu_ru/mepc [50]),
    .i1(data_csr[50]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [50]));
  AL_MUX \cu_ru/m_s_epc/mux6_b51  (
    .i0(\cu_ru/mepc [51]),
    .i1(data_csr[51]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [51]));
  AL_MUX \cu_ru/m_s_epc/mux6_b52  (
    .i0(\cu_ru/mepc [52]),
    .i1(data_csr[52]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [52]));
  AL_MUX \cu_ru/m_s_epc/mux6_b53  (
    .i0(\cu_ru/mepc [53]),
    .i1(data_csr[53]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [53]));
  AL_MUX \cu_ru/m_s_epc/mux6_b54  (
    .i0(\cu_ru/mepc [54]),
    .i1(data_csr[54]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [54]));
  AL_MUX \cu_ru/m_s_epc/mux6_b55  (
    .i0(\cu_ru/mepc [55]),
    .i1(data_csr[55]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [55]));
  AL_MUX \cu_ru/m_s_epc/mux6_b56  (
    .i0(\cu_ru/mepc [56]),
    .i1(data_csr[56]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [56]));
  AL_MUX \cu_ru/m_s_epc/mux6_b57  (
    .i0(\cu_ru/mepc [57]),
    .i1(data_csr[57]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [57]));
  AL_MUX \cu_ru/m_s_epc/mux6_b58  (
    .i0(\cu_ru/mepc [58]),
    .i1(data_csr[58]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [58]));
  AL_MUX \cu_ru/m_s_epc/mux6_b59  (
    .i0(\cu_ru/mepc [59]),
    .i1(data_csr[59]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [59]));
  AL_MUX \cu_ru/m_s_epc/mux6_b6  (
    .i0(\cu_ru/mepc [6]),
    .i1(data_csr[6]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [6]));
  AL_MUX \cu_ru/m_s_epc/mux6_b60  (
    .i0(\cu_ru/mepc [60]),
    .i1(data_csr[60]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [60]));
  AL_MUX \cu_ru/m_s_epc/mux6_b61  (
    .i0(\cu_ru/mepc [61]),
    .i1(data_csr[61]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [61]));
  AL_MUX \cu_ru/m_s_epc/mux6_b62  (
    .i0(\cu_ru/mepc [62]),
    .i1(data_csr[62]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [62]));
  AL_MUX \cu_ru/m_s_epc/mux6_b63  (
    .i0(\cu_ru/mepc [63]),
    .i1(data_csr[63]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [63]));
  AL_MUX \cu_ru/m_s_epc/mux6_b7  (
    .i0(\cu_ru/mepc [7]),
    .i1(data_csr[7]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [7]));
  AL_MUX \cu_ru/m_s_epc/mux6_b8  (
    .i0(\cu_ru/mepc [8]),
    .i1(data_csr[8]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [8]));
  AL_MUX \cu_ru/m_s_epc/mux6_b9  (
    .i0(\cu_ru/mepc [9]),
    .i1(data_csr[9]),
    .sel(\cu_ru/m_s_epc/mux6_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_epc/n9 [9]));
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b0  (
    .i0(\cu_ru/m_s_epc/n9 [0]),
    .i1(\cu_ru/m_s_epc/n2 [0]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b1  (
    .i0(\cu_ru/m_s_epc/n9 [1]),
    .i1(\cu_ru/m_s_epc/n2 [1]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b10  (
    .i0(\cu_ru/m_s_epc/n9 [10]),
    .i1(\cu_ru/m_s_epc/n2 [10]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b11  (
    .i0(\cu_ru/m_s_epc/n9 [11]),
    .i1(\cu_ru/m_s_epc/n2 [11]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b12  (
    .i0(\cu_ru/m_s_epc/n9 [12]),
    .i1(\cu_ru/m_s_epc/n2 [12]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b13  (
    .i0(\cu_ru/m_s_epc/n9 [13]),
    .i1(\cu_ru/m_s_epc/n2 [13]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b14  (
    .i0(\cu_ru/m_s_epc/n9 [14]),
    .i1(\cu_ru/m_s_epc/n2 [14]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b15  (
    .i0(\cu_ru/m_s_epc/n9 [15]),
    .i1(\cu_ru/m_s_epc/n2 [15]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b16  (
    .i0(\cu_ru/m_s_epc/n9 [16]),
    .i1(\cu_ru/m_s_epc/n2 [16]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b17  (
    .i0(\cu_ru/m_s_epc/n9 [17]),
    .i1(\cu_ru/m_s_epc/n2 [17]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b18  (
    .i0(\cu_ru/m_s_epc/n9 [18]),
    .i1(\cu_ru/m_s_epc/n2 [18]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b19  (
    .i0(\cu_ru/m_s_epc/n9 [19]),
    .i1(\cu_ru/m_s_epc/n2 [19]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b2  (
    .i0(\cu_ru/m_s_epc/n9 [2]),
    .i1(\cu_ru/m_s_epc/n2 [2]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b20  (
    .i0(\cu_ru/m_s_epc/n9 [20]),
    .i1(\cu_ru/m_s_epc/n2 [20]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b21  (
    .i0(\cu_ru/m_s_epc/n9 [21]),
    .i1(\cu_ru/m_s_epc/n2 [21]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b22  (
    .i0(\cu_ru/m_s_epc/n9 [22]),
    .i1(\cu_ru/m_s_epc/n2 [22]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b23  (
    .i0(\cu_ru/m_s_epc/n9 [23]),
    .i1(\cu_ru/m_s_epc/n2 [23]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b24  (
    .i0(\cu_ru/m_s_epc/n9 [24]),
    .i1(\cu_ru/m_s_epc/n2 [24]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b25  (
    .i0(\cu_ru/m_s_epc/n9 [25]),
    .i1(\cu_ru/m_s_epc/n2 [25]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b26  (
    .i0(\cu_ru/m_s_epc/n9 [26]),
    .i1(\cu_ru/m_s_epc/n2 [26]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b27  (
    .i0(\cu_ru/m_s_epc/n9 [27]),
    .i1(\cu_ru/m_s_epc/n2 [27]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b28  (
    .i0(\cu_ru/m_s_epc/n9 [28]),
    .i1(\cu_ru/m_s_epc/n2 [28]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b29  (
    .i0(\cu_ru/m_s_epc/n9 [29]),
    .i1(\cu_ru/m_s_epc/n2 [29]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b3  (
    .i0(\cu_ru/m_s_epc/n9 [3]),
    .i1(\cu_ru/m_s_epc/n2 [3]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b30  (
    .i0(\cu_ru/m_s_epc/n9 [30]),
    .i1(\cu_ru/m_s_epc/n2 [30]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b31  (
    .i0(\cu_ru/m_s_epc/n9 [31]),
    .i1(\cu_ru/m_s_epc/n2 [31]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b32  (
    .i0(\cu_ru/m_s_epc/n9 [32]),
    .i1(\cu_ru/m_s_epc/n2 [32]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b33  (
    .i0(\cu_ru/m_s_epc/n9 [33]),
    .i1(\cu_ru/m_s_epc/n2 [33]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b34  (
    .i0(\cu_ru/m_s_epc/n9 [34]),
    .i1(\cu_ru/m_s_epc/n2 [34]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b35  (
    .i0(\cu_ru/m_s_epc/n9 [35]),
    .i1(\cu_ru/m_s_epc/n2 [35]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b36  (
    .i0(\cu_ru/m_s_epc/n9 [36]),
    .i1(\cu_ru/m_s_epc/n2 [36]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b37  (
    .i0(\cu_ru/m_s_epc/n9 [37]),
    .i1(\cu_ru/m_s_epc/n2 [37]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b38  (
    .i0(\cu_ru/m_s_epc/n9 [38]),
    .i1(\cu_ru/m_s_epc/n2 [38]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b39  (
    .i0(\cu_ru/m_s_epc/n9 [39]),
    .i1(\cu_ru/m_s_epc/n2 [39]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b4  (
    .i0(\cu_ru/m_s_epc/n9 [4]),
    .i1(\cu_ru/m_s_epc/n2 [4]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b40  (
    .i0(\cu_ru/m_s_epc/n9 [40]),
    .i1(\cu_ru/m_s_epc/n2 [40]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b41  (
    .i0(\cu_ru/m_s_epc/n9 [41]),
    .i1(\cu_ru/m_s_epc/n2 [41]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b42  (
    .i0(\cu_ru/m_s_epc/n9 [42]),
    .i1(\cu_ru/m_s_epc/n2 [42]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b43  (
    .i0(\cu_ru/m_s_epc/n9 [43]),
    .i1(\cu_ru/m_s_epc/n2 [43]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b44  (
    .i0(\cu_ru/m_s_epc/n9 [44]),
    .i1(\cu_ru/m_s_epc/n2 [44]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b45  (
    .i0(\cu_ru/m_s_epc/n9 [45]),
    .i1(\cu_ru/m_s_epc/n2 [45]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b46  (
    .i0(\cu_ru/m_s_epc/n9 [46]),
    .i1(\cu_ru/m_s_epc/n2 [46]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b47  (
    .i0(\cu_ru/m_s_epc/n9 [47]),
    .i1(\cu_ru/m_s_epc/n2 [47]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b48  (
    .i0(\cu_ru/m_s_epc/n9 [48]),
    .i1(\cu_ru/m_s_epc/n2 [48]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b49  (
    .i0(\cu_ru/m_s_epc/n9 [49]),
    .i1(\cu_ru/m_s_epc/n2 [49]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b5  (
    .i0(\cu_ru/m_s_epc/n9 [5]),
    .i1(\cu_ru/m_s_epc/n2 [5]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b50  (
    .i0(\cu_ru/m_s_epc/n9 [50]),
    .i1(\cu_ru/m_s_epc/n2 [50]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b51  (
    .i0(\cu_ru/m_s_epc/n9 [51]),
    .i1(\cu_ru/m_s_epc/n2 [51]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b52  (
    .i0(\cu_ru/m_s_epc/n9 [52]),
    .i1(\cu_ru/m_s_epc/n2 [52]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b53  (
    .i0(\cu_ru/m_s_epc/n9 [53]),
    .i1(\cu_ru/m_s_epc/n2 [53]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b54  (
    .i0(\cu_ru/m_s_epc/n9 [54]),
    .i1(\cu_ru/m_s_epc/n2 [54]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b55  (
    .i0(\cu_ru/m_s_epc/n9 [55]),
    .i1(\cu_ru/m_s_epc/n2 [55]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b56  (
    .i0(\cu_ru/m_s_epc/n9 [56]),
    .i1(\cu_ru/m_s_epc/n2 [56]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b57  (
    .i0(\cu_ru/m_s_epc/n9 [57]),
    .i1(\cu_ru/m_s_epc/n2 [57]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b58  (
    .i0(\cu_ru/m_s_epc/n9 [58]),
    .i1(\cu_ru/m_s_epc/n2 [58]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b59  (
    .i0(\cu_ru/m_s_epc/n9 [59]),
    .i1(\cu_ru/m_s_epc/n2 [59]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b6  (
    .i0(\cu_ru/m_s_epc/n9 [6]),
    .i1(\cu_ru/m_s_epc/n2 [6]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b60  (
    .i0(\cu_ru/m_s_epc/n9 [60]),
    .i1(\cu_ru/m_s_epc/n2 [60]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b61  (
    .i0(\cu_ru/m_s_epc/n9 [61]),
    .i1(\cu_ru/m_s_epc/n2 [61]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b62  (
    .i0(\cu_ru/m_s_epc/n9 [62]),
    .i1(\cu_ru/m_s_epc/n2 [62]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b63  (
    .i0(\cu_ru/m_s_epc/n9 [63]),
    .i1(\cu_ru/m_s_epc/n2 [63]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b7  (
    .i0(\cu_ru/m_s_epc/n9 [7]),
    .i1(\cu_ru/m_s_epc/n2 [7]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b8  (
    .i0(\cu_ru/m_s_epc/n9 [8]),
    .i1(\cu_ru/m_s_epc/n2 [8]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  binary_mux_s1_w1 \cu_ru/m_s_epc/mux7_b9  (
    .i0(\cu_ru/m_s_epc/n9 [9]),
    .i1(\cu_ru/m_s_epc/n2 [9]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_epc/n10 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(40)
  not \cu_ru/m_s_epc/n3_inv  (\cu_ru/m_s_epc/n3_neg , \cu_ru/m_s_epc/n3 );
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b0  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [0]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b1  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [1]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b10  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [10]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b11  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [11]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b12  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [12]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b13  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [13]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b14  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [14]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b15  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [15]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b16  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [16]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b17  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [17]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b18  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [18]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b19  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [19]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b2  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [2]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b20  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [20]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b21  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [21]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b22  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [22]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b23  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [23]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b24  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [24]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b25  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [25]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b26  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [26]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b27  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [27]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b28  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [28]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b29  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [29]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b3  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [3]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b30  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [30]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b31  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [31]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b32  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [32]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b33  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [33]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b34  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [34]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b35  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [35]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b36  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [36]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b37  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [37]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b38  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [38]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b39  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [39]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b4  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [4]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b40  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [40]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b41  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [41]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b42  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [42]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b43  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [43]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b44  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [44]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b45  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [45]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b46  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [46]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b47  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [47]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b48  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [48]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b49  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [49]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b5  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [5]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b50  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [50]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b51  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [51]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b52  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [52]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b53  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [53]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b54  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [54]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b55  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [55]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b56  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [56]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b57  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [57]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b58  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [58]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b59  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [59]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b6  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [6]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b60  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [60]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b61  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [61]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b62  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [62]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b63  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [63]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b7  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [7]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b8  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [8]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg0_b9  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n8 [9]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sepc [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b0  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b1  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b10  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b11  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b12  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b13  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b14  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b15  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b16  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b17  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b18  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b19  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b2  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b20  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b21  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b22  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b23  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b24  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b25  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b26  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b27  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b28  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b29  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b3  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b30  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b31  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b32  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b33  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b34  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b35  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b36  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b37  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b38  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b39  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b4  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b40  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b41  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b42  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b43  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b44  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b45  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b46  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b47  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b48  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b49  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b5  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b50  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b51  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b52  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b53  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b54  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b55  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b56  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b57  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b58  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b59  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b6  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b60  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b61  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b62  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b63  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b7  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b8  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  reg_sr_as_w1 \cu_ru/m_s_epc/reg1_b9  (
    .clk(clk),
    .d(\cu_ru/m_s_epc/n10 [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mepc [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(41)
  and \cu_ru/m_s_epc/u2  (\cu_ru/m_s_epc/n3 , \cu_ru/mrw_mepc_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(35)
  and \cu_ru/m_s_epc/u3  (\cu_ru/m_s_epc/n4 , \cu_ru/srw_sepc_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_epc.v(38)
  reg_sr_as_w1 \cu_ru/m_s_ie/meie_reg  (
    .clk(clk),
    .d(data_csr[11]),
    .en(\cu_ru/m_s_ie/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sie [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  reg_sr_as_w1 \cu_ru/m_s_ie/msie_reg  (
    .clk(clk),
    .d(data_csr[3]),
    .en(\cu_ru/m_s_ie/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sie [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  reg_sr_as_w1 \cu_ru/m_s_ie/mtie_reg  (
    .clk(clk),
    .d(data_csr[7]),
    .en(\cu_ru/m_s_ie/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sie [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  not \cu_ru/m_s_ie/n0_inv  (\cu_ru/m_s_ie/n0_neg , \cu_ru/m_s_ie/n0 );
  not \cu_ru/m_s_ie/n1_inv  (\cu_ru/m_s_ie/n1_neg , \cu_ru/m_s_ie/n1 );
  reg_sr_as_w1 \cu_ru/m_s_ie/seie_reg  (
    .clk(clk),
    .d(data_csr[9]),
    .en(~\cu_ru/m_s_ie/u11_sel_is_0_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sie [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  reg_sr_as_w1 \cu_ru/m_s_ie/ssie_reg  (
    .clk(clk),
    .d(data_csr[1]),
    .en(~\cu_ru/m_s_ie/u11_sel_is_0_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sie [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  reg_sr_as_w1 \cu_ru/m_s_ie/stie_reg  (
    .clk(clk),
    .d(data_csr[5]),
    .en(~\cu_ru/m_s_ie/u11_sel_is_0_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sie [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(50)
  and \cu_ru/m_s_ie/u11_sel_is_0  (\cu_ru/m_s_ie/u11_sel_is_0_o , \cu_ru/m_s_ie/n0_neg , \cu_ru/m_s_ie/n1_neg );
  and \cu_ru/m_s_ie/u4  (\cu_ru/m_s_ie/n0 , \cu_ru/mrw_mie_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(35)
  and \cu_ru/m_s_ie/u5  (\cu_ru/m_s_ie/n1 , \cu_ru/srw_sie_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_ie.v(43)
  reg_sr_as_w1 \cu_ru/m_s_ip/meip_reg  (
    .clk(clk),
    .d(m_ext_int),
    .en(~\cu_ru/m_s_ip/u12_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sip [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  reg_sr_as_w1 \cu_ru/m_s_ip/msip_reg  (
    .clk(clk),
    .d(m_soft_int),
    .en(~\cu_ru/m_s_ip/u12_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sip [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  reg_sr_as_w1 \cu_ru/m_s_ip/mtip_reg  (
    .clk(clk),
    .d(m_time_int),
    .en(~\cu_ru/m_s_ip/u12_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sip [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  not \cu_ru/m_s_ip/n0_inv  (\cu_ru/m_s_ip/n0_neg , \cu_ru/m_s_ip/n0 );
  not \cu_ru/m_s_ip/n2_inv  (\cu_ru/m_s_ip/n2_neg , \cu_ru/m_s_ip/n2 );
  reg_sr_as_w1 \cu_ru/m_s_ip/seip_reg  (
    .clk(clk),
    .d(\cu_ru/m_s_ip/n1 ),
    .en(\cu_ru/m_s_ip/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_s_ip/seip ));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  reg_sr_as_w1 \cu_ru/m_s_ip/ssip_reg  (
    .clk(clk),
    .d(data_csr[1]),
    .en(~\cu_ru/m_s_ip/u11_sel_is_0_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sip [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  reg_sr_as_w1 \cu_ru/m_s_ip/stip_reg  (
    .clk(clk),
    .d(data_csr[5]),
    .en(\cu_ru/m_s_ip/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/m_sip [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(57)
  and \cu_ru/m_s_ip/u11_sel_is_0  (\cu_ru/m_s_ip/u11_sel_is_0_o , \cu_ru/m_s_ip/n0_neg , \cu_ru/m_s_ip/n2_neg );
  and \cu_ru/m_s_ip/u12_sel_is_2  (\cu_ru/m_s_ip/u12_sel_is_2_o , \cu_ru/m_s_ip/n0_neg , \cu_ru/m_s_ip/n2 );
  or \cu_ru/m_s_ip/u23  (\cu_ru/m_sip [9], \cu_ru/m_s_ip/seip , s_ext_int);  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(59)
  and \cu_ru/m_s_ip/u4  (\cu_ru/m_s_ip/n0 , \cu_ru/mrw_mip_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(41)
  or \cu_ru/m_s_ip/u5  (\cu_ru/m_s_ip/n1 , data_csr[9], s_ext_int);  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(46)
  and \cu_ru/m_s_ip/u6  (\cu_ru/m_s_ip/n2 , \cu_ru/srw_sip_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_ip.v(49)
  and \cu_ru/m_s_scratch/mux2_b0_sel_is_2  (\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o , \cu_ru/m_s_scratch/n0_neg , \cu_ru/m_s_scratch/n1 );
  not \cu_ru/m_s_scratch/n0_inv  (\cu_ru/m_s_scratch/n0_neg , \cu_ru/m_s_scratch/n0 );
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b0  (
    .clk(clk),
    .d(data_csr[0]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b1  (
    .clk(clk),
    .d(data_csr[1]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b10  (
    .clk(clk),
    .d(data_csr[10]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b11  (
    .clk(clk),
    .d(data_csr[11]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b12  (
    .clk(clk),
    .d(data_csr[12]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b13  (
    .clk(clk),
    .d(data_csr[13]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b14  (
    .clk(clk),
    .d(data_csr[14]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b15  (
    .clk(clk),
    .d(data_csr[15]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b16  (
    .clk(clk),
    .d(data_csr[16]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b17  (
    .clk(clk),
    .d(data_csr[17]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b18  (
    .clk(clk),
    .d(data_csr[18]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b19  (
    .clk(clk),
    .d(data_csr[19]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b2  (
    .clk(clk),
    .d(data_csr[2]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b20  (
    .clk(clk),
    .d(data_csr[20]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b21  (
    .clk(clk),
    .d(data_csr[21]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b22  (
    .clk(clk),
    .d(data_csr[22]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b23  (
    .clk(clk),
    .d(data_csr[23]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b24  (
    .clk(clk),
    .d(data_csr[24]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b25  (
    .clk(clk),
    .d(data_csr[25]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b26  (
    .clk(clk),
    .d(data_csr[26]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b27  (
    .clk(clk),
    .d(data_csr[27]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b28  (
    .clk(clk),
    .d(data_csr[28]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b29  (
    .clk(clk),
    .d(data_csr[29]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b3  (
    .clk(clk),
    .d(data_csr[3]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b30  (
    .clk(clk),
    .d(data_csr[30]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b31  (
    .clk(clk),
    .d(data_csr[31]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b32  (
    .clk(clk),
    .d(data_csr[32]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b33  (
    .clk(clk),
    .d(data_csr[33]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b34  (
    .clk(clk),
    .d(data_csr[34]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b35  (
    .clk(clk),
    .d(data_csr[35]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b36  (
    .clk(clk),
    .d(data_csr[36]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b37  (
    .clk(clk),
    .d(data_csr[37]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b38  (
    .clk(clk),
    .d(data_csr[38]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b39  (
    .clk(clk),
    .d(data_csr[39]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b4  (
    .clk(clk),
    .d(data_csr[4]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b40  (
    .clk(clk),
    .d(data_csr[40]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b41  (
    .clk(clk),
    .d(data_csr[41]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b42  (
    .clk(clk),
    .d(data_csr[42]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b43  (
    .clk(clk),
    .d(data_csr[43]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b44  (
    .clk(clk),
    .d(data_csr[44]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b45  (
    .clk(clk),
    .d(data_csr[45]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b46  (
    .clk(clk),
    .d(data_csr[46]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b47  (
    .clk(clk),
    .d(data_csr[47]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b48  (
    .clk(clk),
    .d(data_csr[48]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b49  (
    .clk(clk),
    .d(data_csr[49]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b5  (
    .clk(clk),
    .d(data_csr[5]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b50  (
    .clk(clk),
    .d(data_csr[50]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b51  (
    .clk(clk),
    .d(data_csr[51]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b52  (
    .clk(clk),
    .d(data_csr[52]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b53  (
    .clk(clk),
    .d(data_csr[53]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b54  (
    .clk(clk),
    .d(data_csr[54]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b55  (
    .clk(clk),
    .d(data_csr[55]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b56  (
    .clk(clk),
    .d(data_csr[56]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b57  (
    .clk(clk),
    .d(data_csr[57]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b58  (
    .clk(clk),
    .d(data_csr[58]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b59  (
    .clk(clk),
    .d(data_csr[59]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b6  (
    .clk(clk),
    .d(data_csr[6]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b60  (
    .clk(clk),
    .d(data_csr[60]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b61  (
    .clk(clk),
    .d(data_csr[61]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b62  (
    .clk(clk),
    .d(data_csr[62]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b63  (
    .clk(clk),
    .d(data_csr[63]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b7  (
    .clk(clk),
    .d(data_csr[7]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b8  (
    .clk(clk),
    .d(data_csr[8]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg0_b9  (
    .clk(clk),
    .d(data_csr[9]),
    .en(\cu_ru/m_s_scratch/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mscratch [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b0  (
    .clk(clk),
    .d(data_csr[0]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b1  (
    .clk(clk),
    .d(data_csr[1]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b10  (
    .clk(clk),
    .d(data_csr[10]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b11  (
    .clk(clk),
    .d(data_csr[11]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b12  (
    .clk(clk),
    .d(data_csr[12]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b13  (
    .clk(clk),
    .d(data_csr[13]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b14  (
    .clk(clk),
    .d(data_csr[14]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b15  (
    .clk(clk),
    .d(data_csr[15]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b16  (
    .clk(clk),
    .d(data_csr[16]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b17  (
    .clk(clk),
    .d(data_csr[17]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b18  (
    .clk(clk),
    .d(data_csr[18]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b19  (
    .clk(clk),
    .d(data_csr[19]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b2  (
    .clk(clk),
    .d(data_csr[2]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b20  (
    .clk(clk),
    .d(data_csr[20]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b21  (
    .clk(clk),
    .d(data_csr[21]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b22  (
    .clk(clk),
    .d(data_csr[22]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b23  (
    .clk(clk),
    .d(data_csr[23]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b24  (
    .clk(clk),
    .d(data_csr[24]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b25  (
    .clk(clk),
    .d(data_csr[25]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b26  (
    .clk(clk),
    .d(data_csr[26]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b27  (
    .clk(clk),
    .d(data_csr[27]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b28  (
    .clk(clk),
    .d(data_csr[28]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b29  (
    .clk(clk),
    .d(data_csr[29]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b3  (
    .clk(clk),
    .d(data_csr[3]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b30  (
    .clk(clk),
    .d(data_csr[30]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b31  (
    .clk(clk),
    .d(data_csr[31]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b32  (
    .clk(clk),
    .d(data_csr[32]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b33  (
    .clk(clk),
    .d(data_csr[33]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b34  (
    .clk(clk),
    .d(data_csr[34]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b35  (
    .clk(clk),
    .d(data_csr[35]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b36  (
    .clk(clk),
    .d(data_csr[36]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b37  (
    .clk(clk),
    .d(data_csr[37]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b38  (
    .clk(clk),
    .d(data_csr[38]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b39  (
    .clk(clk),
    .d(data_csr[39]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b4  (
    .clk(clk),
    .d(data_csr[4]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b40  (
    .clk(clk),
    .d(data_csr[40]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b41  (
    .clk(clk),
    .d(data_csr[41]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b42  (
    .clk(clk),
    .d(data_csr[42]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b43  (
    .clk(clk),
    .d(data_csr[43]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b44  (
    .clk(clk),
    .d(data_csr[44]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b45  (
    .clk(clk),
    .d(data_csr[45]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b46  (
    .clk(clk),
    .d(data_csr[46]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b47  (
    .clk(clk),
    .d(data_csr[47]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b48  (
    .clk(clk),
    .d(data_csr[48]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b49  (
    .clk(clk),
    .d(data_csr[49]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b5  (
    .clk(clk),
    .d(data_csr[5]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b50  (
    .clk(clk),
    .d(data_csr[50]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b51  (
    .clk(clk),
    .d(data_csr[51]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b52  (
    .clk(clk),
    .d(data_csr[52]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b53  (
    .clk(clk),
    .d(data_csr[53]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b54  (
    .clk(clk),
    .d(data_csr[54]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b55  (
    .clk(clk),
    .d(data_csr[55]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b56  (
    .clk(clk),
    .d(data_csr[56]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b57  (
    .clk(clk),
    .d(data_csr[57]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b58  (
    .clk(clk),
    .d(data_csr[58]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b59  (
    .clk(clk),
    .d(data_csr[59]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b6  (
    .clk(clk),
    .d(data_csr[6]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b60  (
    .clk(clk),
    .d(data_csr[60]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b61  (
    .clk(clk),
    .d(data_csr[61]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b62  (
    .clk(clk),
    .d(data_csr[62]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b63  (
    .clk(clk),
    .d(data_csr[63]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b7  (
    .clk(clk),
    .d(data_csr[7]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b8  (
    .clk(clk),
    .d(data_csr[8]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  reg_sr_as_w1 \cu_ru/m_s_scratch/reg1_b9  (
    .clk(clk),
    .d(data_csr[9]),
    .en(\cu_ru/m_s_scratch/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/sscratch [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(26)
  and \cu_ru/m_s_scratch/u1  (\cu_ru/m_s_scratch/n0 , \cu_ru/mrw_mscratch_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(20)
  and \cu_ru/m_s_scratch/u2  (\cu_ru/m_s_scratch/n1 , \cu_ru/srw_sscratch_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_scratch.v(23)
  eq_w2 \cu_ru/m_s_status/eq0  (
    .i0(\cu_ru/mstatus [12:11]),
    .i1(2'b11),
    .o(mod_priv[3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(118)
  eq_w2 \cu_ru/m_s_status/eq1  (
    .i0(\cu_ru/mstatus [12:11]),
    .i1(2'b01),
    .o(mod_priv[1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(118)
  eq_w2 \cu_ru/m_s_status/eq2  (
    .i0(\cu_ru/mstatus [12:11]),
    .i1(2'b00),
    .o(mod_priv[0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(131)
  reg_sr_as_w1 \cu_ru/m_s_status/mie_reg  (
    .clk(clk),
    .d(\cu_ru/m_s_status/n37 ),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mie ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/mpie_reg  (
    .clk(clk),
    .d(\cu_ru/m_s_status/n45 ),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mstatus [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/mprv_reg  (
    .clk(clk),
    .d(data_csr[17]),
    .en(\cu_ru/m_s_status/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(mprv));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux0_b1  (
    .i0(\cu_ru/m_s_status/n4 [1]),
    .i1(1'b0),
    .sel(priv[1]),
    .o(\cu_ru/m_s_status/n5 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(103)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux10_b0  (
    .i0(\cu_ru/m_s_status/n63 [0]),
    .i1(\cu_ru/m_s_status/n61 [0]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(\cu_ru/m_s_status/n64 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(122)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux10_b1  (
    .i0(\cu_ru/m_s_status/n63 [1]),
    .i1(\cu_ru/m_s_status/n61 [1]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(\cu_ru/m_s_status/n64 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(122)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux10_b3  (
    .i0(\cu_ru/m_s_status/n63 [3]),
    .i1(\cu_ru/m_s_status/n61 [3]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(\cu_ru/m_s_status/n64 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(122)
  AL_MUX \cu_ru/m_s_status/mux1_b0  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\cu_ru/m_s_status/mux1_b0_sel_is_0_o ),
    .o(\cu_ru/m_s_status/n6 [0]));
  and \cu_ru/m_s_status/mux1_b0_sel_is_0  (\cu_ru/m_s_status/mux1_b0_sel_is_0_o , \priv[3]_neg , \priv[1]_neg );
  binary_mux_s1_w1 \cu_ru/m_s_status/mux1_b1  (
    .i0(\cu_ru/m_s_status/n5 [1]),
    .i1(1'b1),
    .sel(priv[3]),
    .o(\cu_ru/m_s_status/n6 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(103)
  AL_MUX \cu_ru/m_s_status/mux3_b0  (
    .i0(\cu_ru/mstatus [11]),
    .i1(\cu_ru/m_s_status/n6 [0]),
    .sel(\cu_ru/m_s_status/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_status/n21 [0]));
  and \cu_ru/m_s_status/mux3_b0_sel_is_2  (\cu_ru/m_s_status/mux3_b0_sel_is_2_o , \cu_ru/m_s_status/n3_neg , \cu_ru/trap_target_m );
  AL_MUX \cu_ru/m_s_status/mux3_b1  (
    .i0(\cu_ru/mstatus [12]),
    .i1(\cu_ru/m_s_status/n6 [1]),
    .sel(\cu_ru/m_s_status/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_status/n21 [1]));
  binary_mux_s1_w1 \cu_ru/m_s_status/mux4_b0  (
    .i0(\cu_ru/m_s_status/n21 [0]),
    .i1(1'b0),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(\cu_ru/m_s_status/n24 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux4_b1  (
    .i0(\cu_ru/m_s_status/n21 [1]),
    .i1(1'b0),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(\cu_ru/m_s_status/n24 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux5_b0  (
    .i0(\cu_ru/m_s_status/n24 [0]),
    .i1(\cu_ru/mstatus [11]),
    .sel(\cu_ru/m_s_status/n1 ),
    .o(\cu_ru/m_s_status/n35 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux5_b1  (
    .i0(\cu_ru/m_s_status/n24 [1]),
    .i1(\cu_ru/mstatus [12]),
    .sel(\cu_ru/m_s_status/n1 ),
    .o(\cu_ru/m_s_status/n35 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux6_b0  (
    .i0(\cu_ru/m_s_status/n35 [0]),
    .i1(data_csr[11]),
    .sel(\cu_ru/m_s_status/n0 ),
    .o(\cu_ru/m_s_status/n47 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux6_b1  (
    .i0(\cu_ru/m_s_status/n35 [1]),
    .i1(data_csr[12]),
    .sel(\cu_ru/m_s_status/n0 ),
    .o(\cu_ru/m_s_status/n47 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux8_b0  (
    .i0(\cu_ru/m_s_status/n60 [0]),
    .i1(1'b0),
    .sel(mod_priv[3]),
    .o(\cu_ru/m_s_status/n61 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(118)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux8_b1  (
    .i0(mod_priv[1]),
    .i1(1'b0),
    .sel(mod_priv[3]),
    .o(\cu_ru/m_s_status/n61 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(118)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux8_b3  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(mod_priv[3]),
    .o(\cu_ru/m_s_status/n61 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(118)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux9_b0  (
    .i0(priv[0]),
    .i1(\cu_ru/m_s_status/n62 [0]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/m_s_status/n63 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(122)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux9_b1  (
    .i0(priv[1]),
    .i1(\cu_ru/mstatus [8]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/m_s_status/n63 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(122)
  binary_mux_s1_w1 \cu_ru/m_s_status/mux9_b3  (
    .i0(priv[3]),
    .i1(1'b0),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/m_s_status/n63 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(122)
  reg_sr_as_w1 \cu_ru/m_s_status/mxr_reg  (
    .clk(clk),
    .d(data_csr[19]),
    .en(~\cu_ru/m_s_status/u34_sel_is_0_o ),
    .reset(rst),
    .set(1'b0),
    .q(mxr));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  not \cu_ru/m_s_status/n0_inv  (\cu_ru/m_s_status/n0_neg , \cu_ru/m_s_status/n0 );
  not \cu_ru/m_s_status/n1_inv  (\cu_ru/m_s_status/n1_neg , \cu_ru/m_s_status/n1 );
  not \cu_ru/m_s_status/n3_inv  (\cu_ru/m_s_status/n3_neg , \cu_ru/m_s_status/n3 );
  reg_sr_as_w1 \cu_ru/m_s_status/reg0_b0  (
    .clk(clk),
    .d(\cu_ru/m_s_status/n47 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mstatus [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/reg0_b1  (
    .clk(clk),
    .d(\cu_ru/m_s_status/n47 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mstatus [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/reg1_b0  (
    .clk(clk),
    .d(\cu_ru/m_s_status/n64 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(priv[0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  reg_sr_as_w1 \cu_ru/m_s_status/reg1_b1  (
    .clk(clk),
    .d(\cu_ru/m_s_status/n64 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(priv[1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  reg_ar_ss_w1 \cu_ru/m_s_status/reg1_b3  (
    .clk(clk),
    .d(\cu_ru/m_s_status/n64 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(rst),
    .q(priv[3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(123)
  reg_sr_as_w1 \cu_ru/m_s_status/sie_reg  (
    .clk(clk),
    .d(\cu_ru/m_s_status/n36 ),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mstatus [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/spie_reg  (
    .clk(clk),
    .d(\cu_ru/m_s_status/n44 ),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mstatus [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/spp_reg  (
    .clk(clk),
    .d(\cu_ru/m_s_status/n46 ),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mstatus [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/sum_reg  (
    .clk(clk),
    .d(data_csr[18]),
    .en(~\cu_ru/m_s_status/u34_sel_is_0_o ),
    .reset(rst),
    .set(1'b0),
    .q(sum));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/tsr_reg  (
    .clk(clk),
    .d(data_csr[22]),
    .en(\cu_ru/m_s_status/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(tsr));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/tvm_reg  (
    .clk(clk),
    .d(data_csr[20]),
    .en(\cu_ru/m_s_status/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(tvm));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  reg_sr_as_w1 \cu_ru/m_s_status/tw_reg  (
    .clk(clk),
    .d(data_csr[21]),
    .en(\cu_ru/m_s_status/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(tw));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(110)
  AL_MUX \cu_ru/m_s_status/u14  (
    .i0(\cu_ru/mstatus [5]),
    .i1(\cu_ru/mstatus [1]),
    .sel(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .o(\cu_ru/m_s_status/n13 ));
  and \cu_ru/m_s_status/u14_sel_is_2  (\cu_ru/m_s_status/u14_sel_is_2_o , \cu_ru/trap_target_m_neg , \cu_ru/trap_target_s );
  AL_MUX \cu_ru/m_s_status/u15  (
    .i0(\cu_ru/mstatus [1]),
    .i1(1'b0),
    .sel(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .o(\cu_ru/m_s_status/n14 ));
  AL_MUX \cu_ru/m_s_status/u16  (
    .i0(\cu_ru/mstatus [8]),
    .i1(priv[1]),
    .sel(\cu_ru/m_s_status/u14_sel_is_2_o ),
    .o(\cu_ru/m_s_status/n15 ));
  AL_MUX \cu_ru/m_s_status/u17  (
    .i0(\cu_ru/m_s_status/n14 ),
    .i1(\cu_ru/mstatus [5]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/m_s_status/n16 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u18  (
    .i0(\cu_ru/m_s_status/n13 ),
    .i1(1'b0),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/m_s_status/n17 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u19  (
    .i0(\cu_ru/m_s_status/n15 ),
    .i1(1'b0),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/m_s_status/n18 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u20  (
    .i0(\cu_ru/mstatus [7]),
    .i1(\cu_ru/mie ),
    .sel(\cu_ru/m_s_status/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_status/n19 ));
  AL_MUX \cu_ru/m_s_status/u21  (
    .i0(\cu_ru/mie ),
    .i1(1'b0),
    .sel(\cu_ru/m_s_status/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_status/n20 ));
  AL_MUX \cu_ru/m_s_status/u22  (
    .i0(\cu_ru/m_s_status/n20 ),
    .i1(\cu_ru/mstatus [7]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(\cu_ru/m_s_status/n22 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u23  (
    .i0(\cu_ru/m_s_status/n19 ),
    .i1(1'b0),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(\cu_ru/m_s_status/n23 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u24  (
    .i0(\cu_ru/m_s_status/n16 ),
    .i1(\cu_ru/mstatus [1]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(\cu_ru/m_s_status/n25 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u25  (
    .i0(\cu_ru/m_s_status/n17 ),
    .i1(\cu_ru/mstatus [5]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(\cu_ru/m_s_status/n26 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u26  (
    .i0(\cu_ru/m_s_status/n18 ),
    .i1(\cu_ru/mstatus [8]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(\cu_ru/m_s_status/n27 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u32  (
    .i0(\cu_ru/m_s_status/n22 ),
    .i1(\cu_ru/mie ),
    .sel(\cu_ru/m_s_status/n1 ),
    .o(\cu_ru/m_s_status/n33 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u33  (
    .i0(\cu_ru/m_s_status/n23 ),
    .i1(\cu_ru/mstatus [7]),
    .sel(\cu_ru/m_s_status/n1 ),
    .o(\cu_ru/m_s_status/n34 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u34  (
    .i0(data_csr[1]),
    .i1(\cu_ru/m_s_status/n25 ),
    .sel(\cu_ru/m_s_status/u34_sel_is_0_o ),
    .o(\cu_ru/m_s_status/n36 ));
  and \cu_ru/m_s_status/u34_sel_is_0  (\cu_ru/m_s_status/u34_sel_is_0_o , \cu_ru/m_s_status/n0_neg , \cu_ru/m_s_status/n1_neg );
  AL_MUX \cu_ru/m_s_status/u35  (
    .i0(\cu_ru/m_s_status/n33 ),
    .i1(data_csr[3]),
    .sel(\cu_ru/m_s_status/n0 ),
    .o(\cu_ru/m_s_status/n37 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  and \cu_ru/m_s_status/u4  (\cu_ru/m_s_status/n0 , \cu_ru/mrw_mstatus_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(68)
  AL_MUX \cu_ru/m_s_status/u42  (
    .i0(data_csr[5]),
    .i1(\cu_ru/m_s_status/n26 ),
    .sel(\cu_ru/m_s_status/u34_sel_is_0_o ),
    .o(\cu_ru/m_s_status/n44 ));
  AL_MUX \cu_ru/m_s_status/u43  (
    .i0(\cu_ru/m_s_status/n34 ),
    .i1(data_csr[7]),
    .sel(\cu_ru/m_s_status/n0 ),
    .o(\cu_ru/m_s_status/n45 ));  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(109)
  AL_MUX \cu_ru/m_s_status/u44  (
    .i0(data_csr[8]),
    .i1(\cu_ru/m_s_status/n27 ),
    .sel(\cu_ru/m_s_status/u34_sel_is_0_o ),
    .o(\cu_ru/m_s_status/n46 ));
  and \cu_ru/m_s_status/u5  (\cu_ru/m_s_status/n1 , \cu_ru/srw_sstatus_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(83)
  not \cu_ru/m_s_status/u57  (\cu_ru/m_s_status/n62 [0], \cu_ru/mstatus [8]);  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(121)
  not \cu_ru/m_s_status/u59  (\cu_ru/m_s_status/n4 [1], priv[0]);  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(103)
  and \cu_ru/m_s_status/u6  (\cu_ru/m_s_status/n2 , wb_valid, wb_m_ret);  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(90)
  and \cu_ru/m_s_status/u7  (\cu_ru/m_s_status/n3 , wb_valid, wb_s_ret);  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(95)
  not \cu_ru/m_s_status/u8  (\cu_ru/m_s_status/n60 [0], mod_priv[1]);  // ../../RTL/CPU/CU&RU/csrs/m_s_status.v(118)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b0  (
    .i0(wb_exc_code[0]),
    .i1(wb_ins_pc[0]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b1  (
    .i0(wb_exc_code[1]),
    .i1(wb_ins_pc[1]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b10  (
    .i0(wb_exc_code[10]),
    .i1(wb_ins_pc[10]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b11  (
    .i0(wb_exc_code[11]),
    .i1(wb_ins_pc[11]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b12  (
    .i0(wb_exc_code[12]),
    .i1(wb_ins_pc[12]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b13  (
    .i0(wb_exc_code[13]),
    .i1(wb_ins_pc[13]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b14  (
    .i0(wb_exc_code[14]),
    .i1(wb_ins_pc[14]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b15  (
    .i0(wb_exc_code[15]),
    .i1(wb_ins_pc[15]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b16  (
    .i0(wb_exc_code[16]),
    .i1(wb_ins_pc[16]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b17  (
    .i0(wb_exc_code[17]),
    .i1(wb_ins_pc[17]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b18  (
    .i0(wb_exc_code[18]),
    .i1(wb_ins_pc[18]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b19  (
    .i0(wb_exc_code[19]),
    .i1(wb_ins_pc[19]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b2  (
    .i0(wb_exc_code[2]),
    .i1(wb_ins_pc[2]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b20  (
    .i0(wb_exc_code[20]),
    .i1(wb_ins_pc[20]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b21  (
    .i0(wb_exc_code[21]),
    .i1(wb_ins_pc[21]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b22  (
    .i0(wb_exc_code[22]),
    .i1(wb_ins_pc[22]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b23  (
    .i0(wb_exc_code[23]),
    .i1(wb_ins_pc[23]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b24  (
    .i0(wb_exc_code[24]),
    .i1(wb_ins_pc[24]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b25  (
    .i0(wb_exc_code[25]),
    .i1(wb_ins_pc[25]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b26  (
    .i0(wb_exc_code[26]),
    .i1(wb_ins_pc[26]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b27  (
    .i0(wb_exc_code[27]),
    .i1(wb_ins_pc[27]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b28  (
    .i0(wb_exc_code[28]),
    .i1(wb_ins_pc[28]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b29  (
    .i0(wb_exc_code[29]),
    .i1(wb_ins_pc[29]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b3  (
    .i0(wb_exc_code[3]),
    .i1(wb_ins_pc[3]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b30  (
    .i0(wb_exc_code[30]),
    .i1(wb_ins_pc[30]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b31  (
    .i0(wb_exc_code[31]),
    .i1(wb_ins_pc[31]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b32  (
    .i0(wb_exc_code[32]),
    .i1(wb_ins_pc[32]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b33  (
    .i0(wb_exc_code[33]),
    .i1(wb_ins_pc[33]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b34  (
    .i0(wb_exc_code[34]),
    .i1(wb_ins_pc[34]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b35  (
    .i0(wb_exc_code[35]),
    .i1(wb_ins_pc[35]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b36  (
    .i0(wb_exc_code[36]),
    .i1(wb_ins_pc[36]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b37  (
    .i0(wb_exc_code[37]),
    .i1(wb_ins_pc[37]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b38  (
    .i0(wb_exc_code[38]),
    .i1(wb_ins_pc[38]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b39  (
    .i0(wb_exc_code[39]),
    .i1(wb_ins_pc[39]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b4  (
    .i0(wb_exc_code[4]),
    .i1(wb_ins_pc[4]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b40  (
    .i0(wb_exc_code[40]),
    .i1(wb_ins_pc[40]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b41  (
    .i0(wb_exc_code[41]),
    .i1(wb_ins_pc[41]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b42  (
    .i0(wb_exc_code[42]),
    .i1(wb_ins_pc[42]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b43  (
    .i0(wb_exc_code[43]),
    .i1(wb_ins_pc[43]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b44  (
    .i0(wb_exc_code[44]),
    .i1(wb_ins_pc[44]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b45  (
    .i0(wb_exc_code[45]),
    .i1(wb_ins_pc[45]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b46  (
    .i0(wb_exc_code[46]),
    .i1(wb_ins_pc[46]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b47  (
    .i0(wb_exc_code[47]),
    .i1(wb_ins_pc[47]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b48  (
    .i0(wb_exc_code[48]),
    .i1(wb_ins_pc[48]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b49  (
    .i0(wb_exc_code[49]),
    .i1(wb_ins_pc[49]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b5  (
    .i0(wb_exc_code[5]),
    .i1(wb_ins_pc[5]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b50  (
    .i0(wb_exc_code[50]),
    .i1(wb_ins_pc[50]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b51  (
    .i0(wb_exc_code[51]),
    .i1(wb_ins_pc[51]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b52  (
    .i0(wb_exc_code[52]),
    .i1(wb_ins_pc[52]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b53  (
    .i0(wb_exc_code[53]),
    .i1(wb_ins_pc[53]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b54  (
    .i0(wb_exc_code[54]),
    .i1(wb_ins_pc[54]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b55  (
    .i0(wb_exc_code[55]),
    .i1(wb_ins_pc[55]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b56  (
    .i0(wb_exc_code[56]),
    .i1(wb_ins_pc[56]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b57  (
    .i0(wb_exc_code[57]),
    .i1(wb_ins_pc[57]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b58  (
    .i0(wb_exc_code[58]),
    .i1(wb_ins_pc[58]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b59  (
    .i0(wb_exc_code[59]),
    .i1(wb_ins_pc[59]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b6  (
    .i0(wb_exc_code[6]),
    .i1(wb_ins_pc[6]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b60  (
    .i0(wb_exc_code[60]),
    .i1(wb_ins_pc[60]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b61  (
    .i0(wb_exc_code[61]),
    .i1(wb_ins_pc[61]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b62  (
    .i0(wb_exc_code[62]),
    .i1(wb_ins_pc[62]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b63  (
    .i0(wb_exc_code[63]),
    .i1(wb_ins_pc[63]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b7  (
    .i0(wb_exc_code[7]),
    .i1(wb_ins_pc[7]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b8  (
    .i0(wb_exc_code[8]),
    .i1(wb_ins_pc[8]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux0_b9  (
    .i0(wb_exc_code[9]),
    .i1(wb_ins_pc[9]),
    .sel(\cu_ru/m_s_tval/n2 ),
    .o(\cu_ru/m_s_tval/n3 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  AL_MUX \cu_ru/m_s_tval/mux3_b0  (
    .i0(\cu_ru/stval [0]),
    .i1(data_csr[0]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [0]));
  and \cu_ru/m_s_tval/mux3_b0_sel_is_2  (\cu_ru/m_s_tval/mux3_b0_sel_is_2_o , \cu_ru/m_s_tval/n4_neg , \cu_ru/m_s_tval/n5 );
  AL_MUX \cu_ru/m_s_tval/mux3_b1  (
    .i0(\cu_ru/stval [1]),
    .i1(data_csr[1]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [1]));
  AL_MUX \cu_ru/m_s_tval/mux3_b10  (
    .i0(\cu_ru/stval [10]),
    .i1(data_csr[10]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [10]));
  AL_MUX \cu_ru/m_s_tval/mux3_b11  (
    .i0(\cu_ru/stval [11]),
    .i1(data_csr[11]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [11]));
  AL_MUX \cu_ru/m_s_tval/mux3_b12  (
    .i0(\cu_ru/stval [12]),
    .i1(data_csr[12]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [12]));
  AL_MUX \cu_ru/m_s_tval/mux3_b13  (
    .i0(\cu_ru/stval [13]),
    .i1(data_csr[13]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [13]));
  AL_MUX \cu_ru/m_s_tval/mux3_b14  (
    .i0(\cu_ru/stval [14]),
    .i1(data_csr[14]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [14]));
  AL_MUX \cu_ru/m_s_tval/mux3_b15  (
    .i0(\cu_ru/stval [15]),
    .i1(data_csr[15]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [15]));
  AL_MUX \cu_ru/m_s_tval/mux3_b16  (
    .i0(\cu_ru/stval [16]),
    .i1(data_csr[16]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [16]));
  AL_MUX \cu_ru/m_s_tval/mux3_b17  (
    .i0(\cu_ru/stval [17]),
    .i1(data_csr[17]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [17]));
  AL_MUX \cu_ru/m_s_tval/mux3_b18  (
    .i0(\cu_ru/stval [18]),
    .i1(data_csr[18]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [18]));
  AL_MUX \cu_ru/m_s_tval/mux3_b19  (
    .i0(\cu_ru/stval [19]),
    .i1(data_csr[19]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [19]));
  AL_MUX \cu_ru/m_s_tval/mux3_b2  (
    .i0(\cu_ru/stval [2]),
    .i1(data_csr[2]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [2]));
  AL_MUX \cu_ru/m_s_tval/mux3_b20  (
    .i0(\cu_ru/stval [20]),
    .i1(data_csr[20]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [20]));
  AL_MUX \cu_ru/m_s_tval/mux3_b21  (
    .i0(\cu_ru/stval [21]),
    .i1(data_csr[21]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [21]));
  AL_MUX \cu_ru/m_s_tval/mux3_b22  (
    .i0(\cu_ru/stval [22]),
    .i1(data_csr[22]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [22]));
  AL_MUX \cu_ru/m_s_tval/mux3_b23  (
    .i0(\cu_ru/stval [23]),
    .i1(data_csr[23]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [23]));
  AL_MUX \cu_ru/m_s_tval/mux3_b24  (
    .i0(\cu_ru/stval [24]),
    .i1(data_csr[24]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [24]));
  AL_MUX \cu_ru/m_s_tval/mux3_b25  (
    .i0(\cu_ru/stval [25]),
    .i1(data_csr[25]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [25]));
  AL_MUX \cu_ru/m_s_tval/mux3_b26  (
    .i0(\cu_ru/stval [26]),
    .i1(data_csr[26]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [26]));
  AL_MUX \cu_ru/m_s_tval/mux3_b27  (
    .i0(\cu_ru/stval [27]),
    .i1(data_csr[27]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [27]));
  AL_MUX \cu_ru/m_s_tval/mux3_b28  (
    .i0(\cu_ru/stval [28]),
    .i1(data_csr[28]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [28]));
  AL_MUX \cu_ru/m_s_tval/mux3_b29  (
    .i0(\cu_ru/stval [29]),
    .i1(data_csr[29]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [29]));
  AL_MUX \cu_ru/m_s_tval/mux3_b3  (
    .i0(\cu_ru/stval [3]),
    .i1(data_csr[3]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [3]));
  AL_MUX \cu_ru/m_s_tval/mux3_b30  (
    .i0(\cu_ru/stval [30]),
    .i1(data_csr[30]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [30]));
  AL_MUX \cu_ru/m_s_tval/mux3_b31  (
    .i0(\cu_ru/stval [31]),
    .i1(data_csr[31]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [31]));
  AL_MUX \cu_ru/m_s_tval/mux3_b32  (
    .i0(\cu_ru/stval [32]),
    .i1(data_csr[32]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [32]));
  AL_MUX \cu_ru/m_s_tval/mux3_b33  (
    .i0(\cu_ru/stval [33]),
    .i1(data_csr[33]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [33]));
  AL_MUX \cu_ru/m_s_tval/mux3_b34  (
    .i0(\cu_ru/stval [34]),
    .i1(data_csr[34]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [34]));
  AL_MUX \cu_ru/m_s_tval/mux3_b35  (
    .i0(\cu_ru/stval [35]),
    .i1(data_csr[35]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [35]));
  AL_MUX \cu_ru/m_s_tval/mux3_b36  (
    .i0(\cu_ru/stval [36]),
    .i1(data_csr[36]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [36]));
  AL_MUX \cu_ru/m_s_tval/mux3_b37  (
    .i0(\cu_ru/stval [37]),
    .i1(data_csr[37]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [37]));
  AL_MUX \cu_ru/m_s_tval/mux3_b38  (
    .i0(\cu_ru/stval [38]),
    .i1(data_csr[38]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [38]));
  AL_MUX \cu_ru/m_s_tval/mux3_b39  (
    .i0(\cu_ru/stval [39]),
    .i1(data_csr[39]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [39]));
  AL_MUX \cu_ru/m_s_tval/mux3_b4  (
    .i0(\cu_ru/stval [4]),
    .i1(data_csr[4]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [4]));
  AL_MUX \cu_ru/m_s_tval/mux3_b40  (
    .i0(\cu_ru/stval [40]),
    .i1(data_csr[40]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [40]));
  AL_MUX \cu_ru/m_s_tval/mux3_b41  (
    .i0(\cu_ru/stval [41]),
    .i1(data_csr[41]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [41]));
  AL_MUX \cu_ru/m_s_tval/mux3_b42  (
    .i0(\cu_ru/stval [42]),
    .i1(data_csr[42]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [42]));
  AL_MUX \cu_ru/m_s_tval/mux3_b43  (
    .i0(\cu_ru/stval [43]),
    .i1(data_csr[43]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [43]));
  AL_MUX \cu_ru/m_s_tval/mux3_b44  (
    .i0(\cu_ru/stval [44]),
    .i1(data_csr[44]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [44]));
  AL_MUX \cu_ru/m_s_tval/mux3_b45  (
    .i0(\cu_ru/stval [45]),
    .i1(data_csr[45]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [45]));
  AL_MUX \cu_ru/m_s_tval/mux3_b46  (
    .i0(\cu_ru/stval [46]),
    .i1(data_csr[46]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [46]));
  AL_MUX \cu_ru/m_s_tval/mux3_b47  (
    .i0(\cu_ru/stval [47]),
    .i1(data_csr[47]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [47]));
  AL_MUX \cu_ru/m_s_tval/mux3_b48  (
    .i0(\cu_ru/stval [48]),
    .i1(data_csr[48]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [48]));
  AL_MUX \cu_ru/m_s_tval/mux3_b49  (
    .i0(\cu_ru/stval [49]),
    .i1(data_csr[49]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [49]));
  AL_MUX \cu_ru/m_s_tval/mux3_b5  (
    .i0(\cu_ru/stval [5]),
    .i1(data_csr[5]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [5]));
  AL_MUX \cu_ru/m_s_tval/mux3_b50  (
    .i0(\cu_ru/stval [50]),
    .i1(data_csr[50]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [50]));
  AL_MUX \cu_ru/m_s_tval/mux3_b51  (
    .i0(\cu_ru/stval [51]),
    .i1(data_csr[51]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [51]));
  AL_MUX \cu_ru/m_s_tval/mux3_b52  (
    .i0(\cu_ru/stval [52]),
    .i1(data_csr[52]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [52]));
  AL_MUX \cu_ru/m_s_tval/mux3_b53  (
    .i0(\cu_ru/stval [53]),
    .i1(data_csr[53]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [53]));
  AL_MUX \cu_ru/m_s_tval/mux3_b54  (
    .i0(\cu_ru/stval [54]),
    .i1(data_csr[54]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [54]));
  AL_MUX \cu_ru/m_s_tval/mux3_b55  (
    .i0(\cu_ru/stval [55]),
    .i1(data_csr[55]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [55]));
  AL_MUX \cu_ru/m_s_tval/mux3_b56  (
    .i0(\cu_ru/stval [56]),
    .i1(data_csr[56]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [56]));
  AL_MUX \cu_ru/m_s_tval/mux3_b57  (
    .i0(\cu_ru/stval [57]),
    .i1(data_csr[57]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [57]));
  AL_MUX \cu_ru/m_s_tval/mux3_b58  (
    .i0(\cu_ru/stval [58]),
    .i1(data_csr[58]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [58]));
  AL_MUX \cu_ru/m_s_tval/mux3_b59  (
    .i0(\cu_ru/stval [59]),
    .i1(data_csr[59]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [59]));
  AL_MUX \cu_ru/m_s_tval/mux3_b6  (
    .i0(\cu_ru/stval [6]),
    .i1(data_csr[6]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [6]));
  AL_MUX \cu_ru/m_s_tval/mux3_b60  (
    .i0(\cu_ru/stval [60]),
    .i1(data_csr[60]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [60]));
  AL_MUX \cu_ru/m_s_tval/mux3_b61  (
    .i0(\cu_ru/stval [61]),
    .i1(data_csr[61]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [61]));
  AL_MUX \cu_ru/m_s_tval/mux3_b62  (
    .i0(\cu_ru/stval [62]),
    .i1(data_csr[62]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [62]));
  AL_MUX \cu_ru/m_s_tval/mux3_b63  (
    .i0(\cu_ru/stval [63]),
    .i1(data_csr[63]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [63]));
  AL_MUX \cu_ru/m_s_tval/mux3_b7  (
    .i0(\cu_ru/stval [7]),
    .i1(data_csr[7]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [7]));
  AL_MUX \cu_ru/m_s_tval/mux3_b8  (
    .i0(\cu_ru/stval [8]),
    .i1(data_csr[8]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [8]));
  AL_MUX \cu_ru/m_s_tval/mux3_b9  (
    .i0(\cu_ru/stval [9]),
    .i1(data_csr[9]),
    .sel(\cu_ru/m_s_tval/mux3_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n8 [9]));
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b0  (
    .i0(\cu_ru/m_s_tval/n8 [0]),
    .i1(\cu_ru/m_s_tval/n3 [0]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b1  (
    .i0(\cu_ru/m_s_tval/n8 [1]),
    .i1(\cu_ru/m_s_tval/n3 [1]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b10  (
    .i0(\cu_ru/m_s_tval/n8 [10]),
    .i1(\cu_ru/m_s_tval/n3 [10]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b11  (
    .i0(\cu_ru/m_s_tval/n8 [11]),
    .i1(\cu_ru/m_s_tval/n3 [11]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b12  (
    .i0(\cu_ru/m_s_tval/n8 [12]),
    .i1(\cu_ru/m_s_tval/n3 [12]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b13  (
    .i0(\cu_ru/m_s_tval/n8 [13]),
    .i1(\cu_ru/m_s_tval/n3 [13]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b14  (
    .i0(\cu_ru/m_s_tval/n8 [14]),
    .i1(\cu_ru/m_s_tval/n3 [14]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b15  (
    .i0(\cu_ru/m_s_tval/n8 [15]),
    .i1(\cu_ru/m_s_tval/n3 [15]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b16  (
    .i0(\cu_ru/m_s_tval/n8 [16]),
    .i1(\cu_ru/m_s_tval/n3 [16]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b17  (
    .i0(\cu_ru/m_s_tval/n8 [17]),
    .i1(\cu_ru/m_s_tval/n3 [17]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b18  (
    .i0(\cu_ru/m_s_tval/n8 [18]),
    .i1(\cu_ru/m_s_tval/n3 [18]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b19  (
    .i0(\cu_ru/m_s_tval/n8 [19]),
    .i1(\cu_ru/m_s_tval/n3 [19]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b2  (
    .i0(\cu_ru/m_s_tval/n8 [2]),
    .i1(\cu_ru/m_s_tval/n3 [2]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b20  (
    .i0(\cu_ru/m_s_tval/n8 [20]),
    .i1(\cu_ru/m_s_tval/n3 [20]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b21  (
    .i0(\cu_ru/m_s_tval/n8 [21]),
    .i1(\cu_ru/m_s_tval/n3 [21]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b22  (
    .i0(\cu_ru/m_s_tval/n8 [22]),
    .i1(\cu_ru/m_s_tval/n3 [22]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b23  (
    .i0(\cu_ru/m_s_tval/n8 [23]),
    .i1(\cu_ru/m_s_tval/n3 [23]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b24  (
    .i0(\cu_ru/m_s_tval/n8 [24]),
    .i1(\cu_ru/m_s_tval/n3 [24]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b25  (
    .i0(\cu_ru/m_s_tval/n8 [25]),
    .i1(\cu_ru/m_s_tval/n3 [25]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b26  (
    .i0(\cu_ru/m_s_tval/n8 [26]),
    .i1(\cu_ru/m_s_tval/n3 [26]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b27  (
    .i0(\cu_ru/m_s_tval/n8 [27]),
    .i1(\cu_ru/m_s_tval/n3 [27]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b28  (
    .i0(\cu_ru/m_s_tval/n8 [28]),
    .i1(\cu_ru/m_s_tval/n3 [28]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b29  (
    .i0(\cu_ru/m_s_tval/n8 [29]),
    .i1(\cu_ru/m_s_tval/n3 [29]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b3  (
    .i0(\cu_ru/m_s_tval/n8 [3]),
    .i1(\cu_ru/m_s_tval/n3 [3]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b30  (
    .i0(\cu_ru/m_s_tval/n8 [30]),
    .i1(\cu_ru/m_s_tval/n3 [30]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b31  (
    .i0(\cu_ru/m_s_tval/n8 [31]),
    .i1(\cu_ru/m_s_tval/n3 [31]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b32  (
    .i0(\cu_ru/m_s_tval/n8 [32]),
    .i1(\cu_ru/m_s_tval/n3 [32]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b33  (
    .i0(\cu_ru/m_s_tval/n8 [33]),
    .i1(\cu_ru/m_s_tval/n3 [33]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b34  (
    .i0(\cu_ru/m_s_tval/n8 [34]),
    .i1(\cu_ru/m_s_tval/n3 [34]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b35  (
    .i0(\cu_ru/m_s_tval/n8 [35]),
    .i1(\cu_ru/m_s_tval/n3 [35]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b36  (
    .i0(\cu_ru/m_s_tval/n8 [36]),
    .i1(\cu_ru/m_s_tval/n3 [36]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b37  (
    .i0(\cu_ru/m_s_tval/n8 [37]),
    .i1(\cu_ru/m_s_tval/n3 [37]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b38  (
    .i0(\cu_ru/m_s_tval/n8 [38]),
    .i1(\cu_ru/m_s_tval/n3 [38]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b39  (
    .i0(\cu_ru/m_s_tval/n8 [39]),
    .i1(\cu_ru/m_s_tval/n3 [39]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b4  (
    .i0(\cu_ru/m_s_tval/n8 [4]),
    .i1(\cu_ru/m_s_tval/n3 [4]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b40  (
    .i0(\cu_ru/m_s_tval/n8 [40]),
    .i1(\cu_ru/m_s_tval/n3 [40]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b41  (
    .i0(\cu_ru/m_s_tval/n8 [41]),
    .i1(\cu_ru/m_s_tval/n3 [41]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b42  (
    .i0(\cu_ru/m_s_tval/n8 [42]),
    .i1(\cu_ru/m_s_tval/n3 [42]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b43  (
    .i0(\cu_ru/m_s_tval/n8 [43]),
    .i1(\cu_ru/m_s_tval/n3 [43]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b44  (
    .i0(\cu_ru/m_s_tval/n8 [44]),
    .i1(\cu_ru/m_s_tval/n3 [44]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b45  (
    .i0(\cu_ru/m_s_tval/n8 [45]),
    .i1(\cu_ru/m_s_tval/n3 [45]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b46  (
    .i0(\cu_ru/m_s_tval/n8 [46]),
    .i1(\cu_ru/m_s_tval/n3 [46]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b47  (
    .i0(\cu_ru/m_s_tval/n8 [47]),
    .i1(\cu_ru/m_s_tval/n3 [47]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b48  (
    .i0(\cu_ru/m_s_tval/n8 [48]),
    .i1(\cu_ru/m_s_tval/n3 [48]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b49  (
    .i0(\cu_ru/m_s_tval/n8 [49]),
    .i1(\cu_ru/m_s_tval/n3 [49]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b5  (
    .i0(\cu_ru/m_s_tval/n8 [5]),
    .i1(\cu_ru/m_s_tval/n3 [5]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b50  (
    .i0(\cu_ru/m_s_tval/n8 [50]),
    .i1(\cu_ru/m_s_tval/n3 [50]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b51  (
    .i0(\cu_ru/m_s_tval/n8 [51]),
    .i1(\cu_ru/m_s_tval/n3 [51]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b52  (
    .i0(\cu_ru/m_s_tval/n8 [52]),
    .i1(\cu_ru/m_s_tval/n3 [52]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b53  (
    .i0(\cu_ru/m_s_tval/n8 [53]),
    .i1(\cu_ru/m_s_tval/n3 [53]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b54  (
    .i0(\cu_ru/m_s_tval/n8 [54]),
    .i1(\cu_ru/m_s_tval/n3 [54]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b55  (
    .i0(\cu_ru/m_s_tval/n8 [55]),
    .i1(\cu_ru/m_s_tval/n3 [55]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b56  (
    .i0(\cu_ru/m_s_tval/n8 [56]),
    .i1(\cu_ru/m_s_tval/n3 [56]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b57  (
    .i0(\cu_ru/m_s_tval/n8 [57]),
    .i1(\cu_ru/m_s_tval/n3 [57]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b58  (
    .i0(\cu_ru/m_s_tval/n8 [58]),
    .i1(\cu_ru/m_s_tval/n3 [58]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b59  (
    .i0(\cu_ru/m_s_tval/n8 [59]),
    .i1(\cu_ru/m_s_tval/n3 [59]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b6  (
    .i0(\cu_ru/m_s_tval/n8 [6]),
    .i1(\cu_ru/m_s_tval/n3 [6]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b60  (
    .i0(\cu_ru/m_s_tval/n8 [60]),
    .i1(\cu_ru/m_s_tval/n3 [60]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b61  (
    .i0(\cu_ru/m_s_tval/n8 [61]),
    .i1(\cu_ru/m_s_tval/n3 [61]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b62  (
    .i0(\cu_ru/m_s_tval/n8 [62]),
    .i1(\cu_ru/m_s_tval/n3 [62]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b63  (
    .i0(\cu_ru/m_s_tval/n8 [63]),
    .i1(\cu_ru/m_s_tval/n3 [63]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b7  (
    .i0(\cu_ru/m_s_tval/n8 [7]),
    .i1(\cu_ru/m_s_tval/n3 [7]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b8  (
    .i0(\cu_ru/m_s_tval/n8 [8]),
    .i1(\cu_ru/m_s_tval/n3 [8]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux4_b9  (
    .i0(\cu_ru/m_s_tval/n8 [9]),
    .i1(\cu_ru/m_s_tval/n3 [9]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tval/n9 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  AL_MUX \cu_ru/m_s_tval/mux5_b0  (
    .i0(\cu_ru/mtval [0]),
    .i1(data_csr[0]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [0]));
  and \cu_ru/m_s_tval/mux5_b0_sel_is_2  (\cu_ru/m_s_tval/mux5_b0_sel_is_2_o , \cu_ru/trap_target_s_neg , \cu_ru/m_s_tval/n4 );
  AL_MUX \cu_ru/m_s_tval/mux5_b1  (
    .i0(\cu_ru/mtval [1]),
    .i1(data_csr[1]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [1]));
  AL_MUX \cu_ru/m_s_tval/mux5_b10  (
    .i0(\cu_ru/mtval [10]),
    .i1(data_csr[10]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [10]));
  AL_MUX \cu_ru/m_s_tval/mux5_b11  (
    .i0(\cu_ru/mtval [11]),
    .i1(data_csr[11]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [11]));
  AL_MUX \cu_ru/m_s_tval/mux5_b12  (
    .i0(\cu_ru/mtval [12]),
    .i1(data_csr[12]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [12]));
  AL_MUX \cu_ru/m_s_tval/mux5_b13  (
    .i0(\cu_ru/mtval [13]),
    .i1(data_csr[13]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [13]));
  AL_MUX \cu_ru/m_s_tval/mux5_b14  (
    .i0(\cu_ru/mtval [14]),
    .i1(data_csr[14]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [14]));
  AL_MUX \cu_ru/m_s_tval/mux5_b15  (
    .i0(\cu_ru/mtval [15]),
    .i1(data_csr[15]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [15]));
  AL_MUX \cu_ru/m_s_tval/mux5_b16  (
    .i0(\cu_ru/mtval [16]),
    .i1(data_csr[16]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [16]));
  AL_MUX \cu_ru/m_s_tval/mux5_b17  (
    .i0(\cu_ru/mtval [17]),
    .i1(data_csr[17]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [17]));
  AL_MUX \cu_ru/m_s_tval/mux5_b18  (
    .i0(\cu_ru/mtval [18]),
    .i1(data_csr[18]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [18]));
  AL_MUX \cu_ru/m_s_tval/mux5_b19  (
    .i0(\cu_ru/mtval [19]),
    .i1(data_csr[19]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [19]));
  AL_MUX \cu_ru/m_s_tval/mux5_b2  (
    .i0(\cu_ru/mtval [2]),
    .i1(data_csr[2]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [2]));
  AL_MUX \cu_ru/m_s_tval/mux5_b20  (
    .i0(\cu_ru/mtval [20]),
    .i1(data_csr[20]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [20]));
  AL_MUX \cu_ru/m_s_tval/mux5_b21  (
    .i0(\cu_ru/mtval [21]),
    .i1(data_csr[21]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [21]));
  AL_MUX \cu_ru/m_s_tval/mux5_b22  (
    .i0(\cu_ru/mtval [22]),
    .i1(data_csr[22]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [22]));
  AL_MUX \cu_ru/m_s_tval/mux5_b23  (
    .i0(\cu_ru/mtval [23]),
    .i1(data_csr[23]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [23]));
  AL_MUX \cu_ru/m_s_tval/mux5_b24  (
    .i0(\cu_ru/mtval [24]),
    .i1(data_csr[24]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [24]));
  AL_MUX \cu_ru/m_s_tval/mux5_b25  (
    .i0(\cu_ru/mtval [25]),
    .i1(data_csr[25]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [25]));
  AL_MUX \cu_ru/m_s_tval/mux5_b26  (
    .i0(\cu_ru/mtval [26]),
    .i1(data_csr[26]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [26]));
  AL_MUX \cu_ru/m_s_tval/mux5_b27  (
    .i0(\cu_ru/mtval [27]),
    .i1(data_csr[27]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [27]));
  AL_MUX \cu_ru/m_s_tval/mux5_b28  (
    .i0(\cu_ru/mtval [28]),
    .i1(data_csr[28]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [28]));
  AL_MUX \cu_ru/m_s_tval/mux5_b29  (
    .i0(\cu_ru/mtval [29]),
    .i1(data_csr[29]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [29]));
  AL_MUX \cu_ru/m_s_tval/mux5_b3  (
    .i0(\cu_ru/mtval [3]),
    .i1(data_csr[3]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [3]));
  AL_MUX \cu_ru/m_s_tval/mux5_b30  (
    .i0(\cu_ru/mtval [30]),
    .i1(data_csr[30]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [30]));
  AL_MUX \cu_ru/m_s_tval/mux5_b31  (
    .i0(\cu_ru/mtval [31]),
    .i1(data_csr[31]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [31]));
  AL_MUX \cu_ru/m_s_tval/mux5_b32  (
    .i0(\cu_ru/mtval [32]),
    .i1(data_csr[32]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [32]));
  AL_MUX \cu_ru/m_s_tval/mux5_b33  (
    .i0(\cu_ru/mtval [33]),
    .i1(data_csr[33]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [33]));
  AL_MUX \cu_ru/m_s_tval/mux5_b34  (
    .i0(\cu_ru/mtval [34]),
    .i1(data_csr[34]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [34]));
  AL_MUX \cu_ru/m_s_tval/mux5_b35  (
    .i0(\cu_ru/mtval [35]),
    .i1(data_csr[35]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [35]));
  AL_MUX \cu_ru/m_s_tval/mux5_b36  (
    .i0(\cu_ru/mtval [36]),
    .i1(data_csr[36]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [36]));
  AL_MUX \cu_ru/m_s_tval/mux5_b37  (
    .i0(\cu_ru/mtval [37]),
    .i1(data_csr[37]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [37]));
  AL_MUX \cu_ru/m_s_tval/mux5_b38  (
    .i0(\cu_ru/mtval [38]),
    .i1(data_csr[38]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [38]));
  AL_MUX \cu_ru/m_s_tval/mux5_b39  (
    .i0(\cu_ru/mtval [39]),
    .i1(data_csr[39]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [39]));
  AL_MUX \cu_ru/m_s_tval/mux5_b4  (
    .i0(\cu_ru/mtval [4]),
    .i1(data_csr[4]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [4]));
  AL_MUX \cu_ru/m_s_tval/mux5_b40  (
    .i0(\cu_ru/mtval [40]),
    .i1(data_csr[40]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [40]));
  AL_MUX \cu_ru/m_s_tval/mux5_b41  (
    .i0(\cu_ru/mtval [41]),
    .i1(data_csr[41]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [41]));
  AL_MUX \cu_ru/m_s_tval/mux5_b42  (
    .i0(\cu_ru/mtval [42]),
    .i1(data_csr[42]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [42]));
  AL_MUX \cu_ru/m_s_tval/mux5_b43  (
    .i0(\cu_ru/mtval [43]),
    .i1(data_csr[43]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [43]));
  AL_MUX \cu_ru/m_s_tval/mux5_b44  (
    .i0(\cu_ru/mtval [44]),
    .i1(data_csr[44]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [44]));
  AL_MUX \cu_ru/m_s_tval/mux5_b45  (
    .i0(\cu_ru/mtval [45]),
    .i1(data_csr[45]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [45]));
  AL_MUX \cu_ru/m_s_tval/mux5_b46  (
    .i0(\cu_ru/mtval [46]),
    .i1(data_csr[46]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [46]));
  AL_MUX \cu_ru/m_s_tval/mux5_b47  (
    .i0(\cu_ru/mtval [47]),
    .i1(data_csr[47]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [47]));
  AL_MUX \cu_ru/m_s_tval/mux5_b48  (
    .i0(\cu_ru/mtval [48]),
    .i1(data_csr[48]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [48]));
  AL_MUX \cu_ru/m_s_tval/mux5_b49  (
    .i0(\cu_ru/mtval [49]),
    .i1(data_csr[49]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [49]));
  AL_MUX \cu_ru/m_s_tval/mux5_b5  (
    .i0(\cu_ru/mtval [5]),
    .i1(data_csr[5]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [5]));
  AL_MUX \cu_ru/m_s_tval/mux5_b50  (
    .i0(\cu_ru/mtval [50]),
    .i1(data_csr[50]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [50]));
  AL_MUX \cu_ru/m_s_tval/mux5_b51  (
    .i0(\cu_ru/mtval [51]),
    .i1(data_csr[51]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [51]));
  AL_MUX \cu_ru/m_s_tval/mux5_b52  (
    .i0(\cu_ru/mtval [52]),
    .i1(data_csr[52]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [52]));
  AL_MUX \cu_ru/m_s_tval/mux5_b53  (
    .i0(\cu_ru/mtval [53]),
    .i1(data_csr[53]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [53]));
  AL_MUX \cu_ru/m_s_tval/mux5_b54  (
    .i0(\cu_ru/mtval [54]),
    .i1(data_csr[54]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [54]));
  AL_MUX \cu_ru/m_s_tval/mux5_b55  (
    .i0(\cu_ru/mtval [55]),
    .i1(data_csr[55]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [55]));
  AL_MUX \cu_ru/m_s_tval/mux5_b56  (
    .i0(\cu_ru/mtval [56]),
    .i1(data_csr[56]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [56]));
  AL_MUX \cu_ru/m_s_tval/mux5_b57  (
    .i0(\cu_ru/mtval [57]),
    .i1(data_csr[57]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [57]));
  AL_MUX \cu_ru/m_s_tval/mux5_b58  (
    .i0(\cu_ru/mtval [58]),
    .i1(data_csr[58]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [58]));
  AL_MUX \cu_ru/m_s_tval/mux5_b59  (
    .i0(\cu_ru/mtval [59]),
    .i1(data_csr[59]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [59]));
  AL_MUX \cu_ru/m_s_tval/mux5_b6  (
    .i0(\cu_ru/mtval [6]),
    .i1(data_csr[6]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [6]));
  AL_MUX \cu_ru/m_s_tval/mux5_b60  (
    .i0(\cu_ru/mtval [60]),
    .i1(data_csr[60]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [60]));
  AL_MUX \cu_ru/m_s_tval/mux5_b61  (
    .i0(\cu_ru/mtval [61]),
    .i1(data_csr[61]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [61]));
  AL_MUX \cu_ru/m_s_tval/mux5_b62  (
    .i0(\cu_ru/mtval [62]),
    .i1(data_csr[62]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [62]));
  AL_MUX \cu_ru/m_s_tval/mux5_b63  (
    .i0(\cu_ru/mtval [63]),
    .i1(data_csr[63]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [63]));
  AL_MUX \cu_ru/m_s_tval/mux5_b7  (
    .i0(\cu_ru/mtval [7]),
    .i1(data_csr[7]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [7]));
  AL_MUX \cu_ru/m_s_tval/mux5_b8  (
    .i0(\cu_ru/mtval [8]),
    .i1(data_csr[8]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [8]));
  AL_MUX \cu_ru/m_s_tval/mux5_b9  (
    .i0(\cu_ru/mtval [9]),
    .i1(data_csr[9]),
    .sel(\cu_ru/m_s_tval/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/m_s_tval/n10 [9]));
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b0  (
    .i0(\cu_ru/m_s_tval/n10 [0]),
    .i1(\cu_ru/m_s_tval/n3 [0]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b1  (
    .i0(\cu_ru/m_s_tval/n10 [1]),
    .i1(\cu_ru/m_s_tval/n3 [1]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b10  (
    .i0(\cu_ru/m_s_tval/n10 [10]),
    .i1(\cu_ru/m_s_tval/n3 [10]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b11  (
    .i0(\cu_ru/m_s_tval/n10 [11]),
    .i1(\cu_ru/m_s_tval/n3 [11]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b12  (
    .i0(\cu_ru/m_s_tval/n10 [12]),
    .i1(\cu_ru/m_s_tval/n3 [12]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b13  (
    .i0(\cu_ru/m_s_tval/n10 [13]),
    .i1(\cu_ru/m_s_tval/n3 [13]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b14  (
    .i0(\cu_ru/m_s_tval/n10 [14]),
    .i1(\cu_ru/m_s_tval/n3 [14]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b15  (
    .i0(\cu_ru/m_s_tval/n10 [15]),
    .i1(\cu_ru/m_s_tval/n3 [15]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b16  (
    .i0(\cu_ru/m_s_tval/n10 [16]),
    .i1(\cu_ru/m_s_tval/n3 [16]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b17  (
    .i0(\cu_ru/m_s_tval/n10 [17]),
    .i1(\cu_ru/m_s_tval/n3 [17]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b18  (
    .i0(\cu_ru/m_s_tval/n10 [18]),
    .i1(\cu_ru/m_s_tval/n3 [18]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b19  (
    .i0(\cu_ru/m_s_tval/n10 [19]),
    .i1(\cu_ru/m_s_tval/n3 [19]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b2  (
    .i0(\cu_ru/m_s_tval/n10 [2]),
    .i1(\cu_ru/m_s_tval/n3 [2]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b20  (
    .i0(\cu_ru/m_s_tval/n10 [20]),
    .i1(\cu_ru/m_s_tval/n3 [20]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b21  (
    .i0(\cu_ru/m_s_tval/n10 [21]),
    .i1(\cu_ru/m_s_tval/n3 [21]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b22  (
    .i0(\cu_ru/m_s_tval/n10 [22]),
    .i1(\cu_ru/m_s_tval/n3 [22]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b23  (
    .i0(\cu_ru/m_s_tval/n10 [23]),
    .i1(\cu_ru/m_s_tval/n3 [23]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b24  (
    .i0(\cu_ru/m_s_tval/n10 [24]),
    .i1(\cu_ru/m_s_tval/n3 [24]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b25  (
    .i0(\cu_ru/m_s_tval/n10 [25]),
    .i1(\cu_ru/m_s_tval/n3 [25]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b26  (
    .i0(\cu_ru/m_s_tval/n10 [26]),
    .i1(\cu_ru/m_s_tval/n3 [26]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b27  (
    .i0(\cu_ru/m_s_tval/n10 [27]),
    .i1(\cu_ru/m_s_tval/n3 [27]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b28  (
    .i0(\cu_ru/m_s_tval/n10 [28]),
    .i1(\cu_ru/m_s_tval/n3 [28]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b29  (
    .i0(\cu_ru/m_s_tval/n10 [29]),
    .i1(\cu_ru/m_s_tval/n3 [29]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b3  (
    .i0(\cu_ru/m_s_tval/n10 [3]),
    .i1(\cu_ru/m_s_tval/n3 [3]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b30  (
    .i0(\cu_ru/m_s_tval/n10 [30]),
    .i1(\cu_ru/m_s_tval/n3 [30]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b31  (
    .i0(\cu_ru/m_s_tval/n10 [31]),
    .i1(\cu_ru/m_s_tval/n3 [31]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b32  (
    .i0(\cu_ru/m_s_tval/n10 [32]),
    .i1(\cu_ru/m_s_tval/n3 [32]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b33  (
    .i0(\cu_ru/m_s_tval/n10 [33]),
    .i1(\cu_ru/m_s_tval/n3 [33]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b34  (
    .i0(\cu_ru/m_s_tval/n10 [34]),
    .i1(\cu_ru/m_s_tval/n3 [34]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b35  (
    .i0(\cu_ru/m_s_tval/n10 [35]),
    .i1(\cu_ru/m_s_tval/n3 [35]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b36  (
    .i0(\cu_ru/m_s_tval/n10 [36]),
    .i1(\cu_ru/m_s_tval/n3 [36]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b37  (
    .i0(\cu_ru/m_s_tval/n10 [37]),
    .i1(\cu_ru/m_s_tval/n3 [37]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b38  (
    .i0(\cu_ru/m_s_tval/n10 [38]),
    .i1(\cu_ru/m_s_tval/n3 [38]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b39  (
    .i0(\cu_ru/m_s_tval/n10 [39]),
    .i1(\cu_ru/m_s_tval/n3 [39]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b4  (
    .i0(\cu_ru/m_s_tval/n10 [4]),
    .i1(\cu_ru/m_s_tval/n3 [4]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b40  (
    .i0(\cu_ru/m_s_tval/n10 [40]),
    .i1(\cu_ru/m_s_tval/n3 [40]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b41  (
    .i0(\cu_ru/m_s_tval/n10 [41]),
    .i1(\cu_ru/m_s_tval/n3 [41]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b42  (
    .i0(\cu_ru/m_s_tval/n10 [42]),
    .i1(\cu_ru/m_s_tval/n3 [42]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b43  (
    .i0(\cu_ru/m_s_tval/n10 [43]),
    .i1(\cu_ru/m_s_tval/n3 [43]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b44  (
    .i0(\cu_ru/m_s_tval/n10 [44]),
    .i1(\cu_ru/m_s_tval/n3 [44]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b45  (
    .i0(\cu_ru/m_s_tval/n10 [45]),
    .i1(\cu_ru/m_s_tval/n3 [45]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b46  (
    .i0(\cu_ru/m_s_tval/n10 [46]),
    .i1(\cu_ru/m_s_tval/n3 [46]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b47  (
    .i0(\cu_ru/m_s_tval/n10 [47]),
    .i1(\cu_ru/m_s_tval/n3 [47]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b48  (
    .i0(\cu_ru/m_s_tval/n10 [48]),
    .i1(\cu_ru/m_s_tval/n3 [48]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b49  (
    .i0(\cu_ru/m_s_tval/n10 [49]),
    .i1(\cu_ru/m_s_tval/n3 [49]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b5  (
    .i0(\cu_ru/m_s_tval/n10 [5]),
    .i1(\cu_ru/m_s_tval/n3 [5]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b50  (
    .i0(\cu_ru/m_s_tval/n10 [50]),
    .i1(\cu_ru/m_s_tval/n3 [50]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b51  (
    .i0(\cu_ru/m_s_tval/n10 [51]),
    .i1(\cu_ru/m_s_tval/n3 [51]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b52  (
    .i0(\cu_ru/m_s_tval/n10 [52]),
    .i1(\cu_ru/m_s_tval/n3 [52]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b53  (
    .i0(\cu_ru/m_s_tval/n10 [53]),
    .i1(\cu_ru/m_s_tval/n3 [53]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b54  (
    .i0(\cu_ru/m_s_tval/n10 [54]),
    .i1(\cu_ru/m_s_tval/n3 [54]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b55  (
    .i0(\cu_ru/m_s_tval/n10 [55]),
    .i1(\cu_ru/m_s_tval/n3 [55]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b56  (
    .i0(\cu_ru/m_s_tval/n10 [56]),
    .i1(\cu_ru/m_s_tval/n3 [56]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b57  (
    .i0(\cu_ru/m_s_tval/n10 [57]),
    .i1(\cu_ru/m_s_tval/n3 [57]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b58  (
    .i0(\cu_ru/m_s_tval/n10 [58]),
    .i1(\cu_ru/m_s_tval/n3 [58]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b59  (
    .i0(\cu_ru/m_s_tval/n10 [59]),
    .i1(\cu_ru/m_s_tval/n3 [59]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b6  (
    .i0(\cu_ru/m_s_tval/n10 [6]),
    .i1(\cu_ru/m_s_tval/n3 [6]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b60  (
    .i0(\cu_ru/m_s_tval/n10 [60]),
    .i1(\cu_ru/m_s_tval/n3 [60]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b61  (
    .i0(\cu_ru/m_s_tval/n10 [61]),
    .i1(\cu_ru/m_s_tval/n3 [61]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b62  (
    .i0(\cu_ru/m_s_tval/n10 [62]),
    .i1(\cu_ru/m_s_tval/n3 [62]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b63  (
    .i0(\cu_ru/m_s_tval/n10 [63]),
    .i1(\cu_ru/m_s_tval/n3 [63]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b7  (
    .i0(\cu_ru/m_s_tval/n10 [7]),
    .i1(\cu_ru/m_s_tval/n3 [7]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b8  (
    .i0(\cu_ru/m_s_tval/n10 [8]),
    .i1(\cu_ru/m_s_tval/n3 [8]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  binary_mux_s1_w1 \cu_ru/m_s_tval/mux6_b9  (
    .i0(\cu_ru/m_s_tval/n10 [9]),
    .i1(\cu_ru/m_s_tval/n3 [9]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/m_s_tval/n11 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(55)
  not \cu_ru/m_s_tval/n4_inv  (\cu_ru/m_s_tval/n4_neg , \cu_ru/m_s_tval/n4 );
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b0  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [0]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b1  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [1]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b10  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [10]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b11  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [11]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b12  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [12]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b13  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [13]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b14  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [14]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b15  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [15]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b16  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [16]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b17  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [17]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b18  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [18]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b19  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [19]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b2  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [2]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b20  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [20]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b21  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [21]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b22  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [22]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b23  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [23]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b24  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [24]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b25  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [25]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b26  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [26]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b27  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [27]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b28  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [28]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b29  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [29]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b3  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [3]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b30  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [30]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b31  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [31]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b32  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [32]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b33  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [33]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b34  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [34]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b35  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [35]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b36  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [36]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b37  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [37]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b38  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [38]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b39  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [39]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b4  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [4]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b40  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [40]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b41  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [41]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b42  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [42]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b43  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [43]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b44  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [44]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b45  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [45]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b46  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [46]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b47  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [47]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b48  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [48]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b49  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [49]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b5  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [5]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b50  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [50]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b51  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [51]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b52  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [52]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b53  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [53]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b54  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [54]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b55  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [55]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b56  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [56]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b57  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [57]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b58  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [58]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b59  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [59]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b6  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [6]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b60  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [60]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b61  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [61]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b62  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [62]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b63  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [63]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b7  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [7]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b8  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [8]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg0_b9  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n9 [9]),
    .en(~\cu_ru/trap_target_m ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stval [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b0  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b1  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b10  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b11  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b12  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b13  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b14  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b15  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b16  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b17  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b18  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b19  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b2  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b20  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b21  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b22  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b23  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b24  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b25  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b26  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b27  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b28  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b29  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b3  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b30  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b31  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b32  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b33  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b34  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b35  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b36  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b37  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b38  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b39  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b4  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b40  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b41  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b42  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b43  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b44  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b45  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b46  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b47  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b48  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b49  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b5  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b50  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b51  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b52  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b53  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b54  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b55  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b56  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b57  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b58  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b59  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b6  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b60  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b61  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b62  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b63  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b7  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b8  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  reg_sr_as_w1 \cu_ru/m_s_tval/reg1_b9  (
    .clk(clk),
    .d(\cu_ru/m_s_tval/n11 [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtval [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(56)
  or \cu_ru/m_s_tval/u1  (\cu_ru/m_s_tval/n0 , wb_ins_acc_fault, wb_ins_addr_mis);  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  or \cu_ru/m_s_tval/u2  (\cu_ru/m_s_tval/n1 , \cu_ru/m_s_tval/n0 , wb_ins_page_fault);  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  or \cu_ru/m_s_tval/u3  (\cu_ru/m_s_tval/n2 , \cu_ru/m_s_tval/n1 , wb_ebreak);  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(45)
  and \cu_ru/m_s_tval/u4  (\cu_ru/m_s_tval/n4 , \cu_ru/mrw_mtval_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(50)
  and \cu_ru/m_s_tval/u5  (\cu_ru/m_s_tval/n5 , \cu_ru/srw_stval_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_tval.v(53)
  and \cu_ru/m_s_tvec/mux2_b0_sel_is_2  (\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o , \cu_ru/m_s_tvec/n0_neg , \cu_ru/m_s_tvec/n1 );
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b0  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [0]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b10  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [10]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b11  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [11]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b12  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [12]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b13  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [13]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b14  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [14]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b15  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [15]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b16  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [16]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b17  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [17]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b18  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [18]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b19  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [19]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b2  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [2]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b20  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [20]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b21  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [21]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b22  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [22]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b23  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [23]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b24  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [24]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b25  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [25]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b26  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [26]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b27  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [27]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b28  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [28]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b29  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [29]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b3  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [3]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b30  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [30]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b31  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [31]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b32  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [32]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b33  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [33]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b34  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [34]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b35  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [35]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b36  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [36]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b37  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [37]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b38  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [38]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b39  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [39]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b4  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [4]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b40  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [40]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b41  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [41]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b42  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [42]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b43  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [43]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b44  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [44]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b45  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [45]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b46  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [46]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b47  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [47]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b48  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [48]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b49  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [49]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b5  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [5]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b50  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [50]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b51  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [51]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b52  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [52]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b53  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [53]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b54  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [54]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b55  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [55]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b56  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [56]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b57  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [57]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b58  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [58]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b59  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [59]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b6  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [6]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b60  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [60]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b61  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [61]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b62  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [62]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b63  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [63]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b7  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [7]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b8  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [8]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux5_b9  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [9]),
    .sel(\cu_ru/trap_target_s ),
    .o(\cu_ru/m_s_tvec/n7 [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b0  (
    .i0(\cu_ru/m_s_tvec/n7 [0]),
    .i1(\cu_ru/mtvec [0]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b10  (
    .i0(\cu_ru/m_s_tvec/n7 [10]),
    .i1(\cu_ru/mtvec [10]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b11  (
    .i0(\cu_ru/m_s_tvec/n7 [11]),
    .i1(\cu_ru/mtvec [11]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b12  (
    .i0(\cu_ru/m_s_tvec/n7 [12]),
    .i1(\cu_ru/mtvec [12]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b13  (
    .i0(\cu_ru/m_s_tvec/n7 [13]),
    .i1(\cu_ru/mtvec [13]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b14  (
    .i0(\cu_ru/m_s_tvec/n7 [14]),
    .i1(\cu_ru/mtvec [14]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b15  (
    .i0(\cu_ru/m_s_tvec/n7 [15]),
    .i1(\cu_ru/mtvec [15]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b16  (
    .i0(\cu_ru/m_s_tvec/n7 [16]),
    .i1(\cu_ru/mtvec [16]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b17  (
    .i0(\cu_ru/m_s_tvec/n7 [17]),
    .i1(\cu_ru/mtvec [17]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b18  (
    .i0(\cu_ru/m_s_tvec/n7 [18]),
    .i1(\cu_ru/mtvec [18]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b19  (
    .i0(\cu_ru/m_s_tvec/n7 [19]),
    .i1(\cu_ru/mtvec [19]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b2  (
    .i0(\cu_ru/m_s_tvec/n7 [2]),
    .i1(\cu_ru/mtvec [2]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b20  (
    .i0(\cu_ru/m_s_tvec/n7 [20]),
    .i1(\cu_ru/mtvec [20]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b21  (
    .i0(\cu_ru/m_s_tvec/n7 [21]),
    .i1(\cu_ru/mtvec [21]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b22  (
    .i0(\cu_ru/m_s_tvec/n7 [22]),
    .i1(\cu_ru/mtvec [22]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b23  (
    .i0(\cu_ru/m_s_tvec/n7 [23]),
    .i1(\cu_ru/mtvec [23]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b24  (
    .i0(\cu_ru/m_s_tvec/n7 [24]),
    .i1(\cu_ru/mtvec [24]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b25  (
    .i0(\cu_ru/m_s_tvec/n7 [25]),
    .i1(\cu_ru/mtvec [25]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b26  (
    .i0(\cu_ru/m_s_tvec/n7 [26]),
    .i1(\cu_ru/mtvec [26]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b27  (
    .i0(\cu_ru/m_s_tvec/n7 [27]),
    .i1(\cu_ru/mtvec [27]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b28  (
    .i0(\cu_ru/m_s_tvec/n7 [28]),
    .i1(\cu_ru/mtvec [28]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b29  (
    .i0(\cu_ru/m_s_tvec/n7 [29]),
    .i1(\cu_ru/mtvec [29]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b3  (
    .i0(\cu_ru/m_s_tvec/n7 [3]),
    .i1(\cu_ru/mtvec [3]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b30  (
    .i0(\cu_ru/m_s_tvec/n7 [30]),
    .i1(\cu_ru/mtvec [30]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b31  (
    .i0(\cu_ru/m_s_tvec/n7 [31]),
    .i1(\cu_ru/mtvec [31]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b32  (
    .i0(\cu_ru/m_s_tvec/n7 [32]),
    .i1(\cu_ru/mtvec [32]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b33  (
    .i0(\cu_ru/m_s_tvec/n7 [33]),
    .i1(\cu_ru/mtvec [33]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b34  (
    .i0(\cu_ru/m_s_tvec/n7 [34]),
    .i1(\cu_ru/mtvec [34]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b35  (
    .i0(\cu_ru/m_s_tvec/n7 [35]),
    .i1(\cu_ru/mtvec [35]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b36  (
    .i0(\cu_ru/m_s_tvec/n7 [36]),
    .i1(\cu_ru/mtvec [36]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b37  (
    .i0(\cu_ru/m_s_tvec/n7 [37]),
    .i1(\cu_ru/mtvec [37]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b38  (
    .i0(\cu_ru/m_s_tvec/n7 [38]),
    .i1(\cu_ru/mtvec [38]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b39  (
    .i0(\cu_ru/m_s_tvec/n7 [39]),
    .i1(\cu_ru/mtvec [39]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b4  (
    .i0(\cu_ru/m_s_tvec/n7 [4]),
    .i1(\cu_ru/mtvec [4]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b40  (
    .i0(\cu_ru/m_s_tvec/n7 [40]),
    .i1(\cu_ru/mtvec [40]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b41  (
    .i0(\cu_ru/m_s_tvec/n7 [41]),
    .i1(\cu_ru/mtvec [41]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b42  (
    .i0(\cu_ru/m_s_tvec/n7 [42]),
    .i1(\cu_ru/mtvec [42]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b43  (
    .i0(\cu_ru/m_s_tvec/n7 [43]),
    .i1(\cu_ru/mtvec [43]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b44  (
    .i0(\cu_ru/m_s_tvec/n7 [44]),
    .i1(\cu_ru/mtvec [44]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b45  (
    .i0(\cu_ru/m_s_tvec/n7 [45]),
    .i1(\cu_ru/mtvec [45]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b46  (
    .i0(\cu_ru/m_s_tvec/n7 [46]),
    .i1(\cu_ru/mtvec [46]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b47  (
    .i0(\cu_ru/m_s_tvec/n7 [47]),
    .i1(\cu_ru/mtvec [47]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b48  (
    .i0(\cu_ru/m_s_tvec/n7 [48]),
    .i1(\cu_ru/mtvec [48]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b49  (
    .i0(\cu_ru/m_s_tvec/n7 [49]),
    .i1(\cu_ru/mtvec [49]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b5  (
    .i0(\cu_ru/m_s_tvec/n7 [5]),
    .i1(\cu_ru/mtvec [5]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b50  (
    .i0(\cu_ru/m_s_tvec/n7 [50]),
    .i1(\cu_ru/mtvec [50]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b51  (
    .i0(\cu_ru/m_s_tvec/n7 [51]),
    .i1(\cu_ru/mtvec [51]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b52  (
    .i0(\cu_ru/m_s_tvec/n7 [52]),
    .i1(\cu_ru/mtvec [52]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b53  (
    .i0(\cu_ru/m_s_tvec/n7 [53]),
    .i1(\cu_ru/mtvec [53]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b54  (
    .i0(\cu_ru/m_s_tvec/n7 [54]),
    .i1(\cu_ru/mtvec [54]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b55  (
    .i0(\cu_ru/m_s_tvec/n7 [55]),
    .i1(\cu_ru/mtvec [55]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b56  (
    .i0(\cu_ru/m_s_tvec/n7 [56]),
    .i1(\cu_ru/mtvec [56]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b57  (
    .i0(\cu_ru/m_s_tvec/n7 [57]),
    .i1(\cu_ru/mtvec [57]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b58  (
    .i0(\cu_ru/m_s_tvec/n7 [58]),
    .i1(\cu_ru/mtvec [58]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b59  (
    .i0(\cu_ru/m_s_tvec/n7 [59]),
    .i1(\cu_ru/mtvec [59]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b6  (
    .i0(\cu_ru/m_s_tvec/n7 [6]),
    .i1(\cu_ru/mtvec [6]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b60  (
    .i0(\cu_ru/m_s_tvec/n7 [60]),
    .i1(\cu_ru/mtvec [60]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b61  (
    .i0(\cu_ru/m_s_tvec/n7 [61]),
    .i1(\cu_ru/mtvec [61]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b62  (
    .i0(\cu_ru/m_s_tvec/n7 [62]),
    .i1(\cu_ru/mtvec [62]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b63  (
    .i0(\cu_ru/m_s_tvec/n7 [63]),
    .i1(\cu_ru/mtvec [63]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b7  (
    .i0(\cu_ru/m_s_tvec/n7 [7]),
    .i1(\cu_ru/mtvec [7]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b8  (
    .i0(\cu_ru/m_s_tvec/n7 [8]),
    .i1(\cu_ru/mtvec [8]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  binary_mux_s1_w1 \cu_ru/m_s_tvec/mux6_b9  (
    .i0(\cu_ru/m_s_tvec/n7 [9]),
    .i1(\cu_ru/mtvec [9]),
    .sel(\cu_ru/trap_target_m ),
    .o(\cu_ru/tvec [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(34)
  not \cu_ru/m_s_tvec/n0_inv  (\cu_ru/m_s_tvec/n0_neg , \cu_ru/m_s_tvec/n0 );
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b0  (
    .clk(clk),
    .d(csr_data[0]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b1  (
    .clk(clk),
    .d(csr_data[1]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b10  (
    .clk(clk),
    .d(csr_data[10]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b11  (
    .clk(clk),
    .d(csr_data[11]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b12  (
    .clk(clk),
    .d(csr_data[12]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b13  (
    .clk(clk),
    .d(csr_data[13]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b14  (
    .clk(clk),
    .d(csr_data[14]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b15  (
    .clk(clk),
    .d(csr_data[15]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b16  (
    .clk(clk),
    .d(csr_data[16]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b17  (
    .clk(clk),
    .d(csr_data[17]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b18  (
    .clk(clk),
    .d(csr_data[18]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b19  (
    .clk(clk),
    .d(csr_data[19]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b2  (
    .clk(clk),
    .d(csr_data[2]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b20  (
    .clk(clk),
    .d(csr_data[20]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b21  (
    .clk(clk),
    .d(csr_data[21]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b22  (
    .clk(clk),
    .d(csr_data[22]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b23  (
    .clk(clk),
    .d(csr_data[23]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b24  (
    .clk(clk),
    .d(csr_data[24]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b25  (
    .clk(clk),
    .d(csr_data[25]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b26  (
    .clk(clk),
    .d(csr_data[26]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b27  (
    .clk(clk),
    .d(csr_data[27]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b28  (
    .clk(clk),
    .d(csr_data[28]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b29  (
    .clk(clk),
    .d(csr_data[29]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b3  (
    .clk(clk),
    .d(csr_data[3]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b30  (
    .clk(clk),
    .d(csr_data[30]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b31  (
    .clk(clk),
    .d(csr_data[31]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b32  (
    .clk(clk),
    .d(csr_data[32]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b33  (
    .clk(clk),
    .d(csr_data[33]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b34  (
    .clk(clk),
    .d(csr_data[34]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b35  (
    .clk(clk),
    .d(csr_data[35]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b36  (
    .clk(clk),
    .d(csr_data[36]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b37  (
    .clk(clk),
    .d(csr_data[37]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b38  (
    .clk(clk),
    .d(csr_data[38]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b39  (
    .clk(clk),
    .d(csr_data[39]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b4  (
    .clk(clk),
    .d(csr_data[4]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b40  (
    .clk(clk),
    .d(csr_data[40]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b41  (
    .clk(clk),
    .d(csr_data[41]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b42  (
    .clk(clk),
    .d(csr_data[42]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b43  (
    .clk(clk),
    .d(csr_data[43]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b44  (
    .clk(clk),
    .d(csr_data[44]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b45  (
    .clk(clk),
    .d(csr_data[45]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b46  (
    .clk(clk),
    .d(csr_data[46]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b47  (
    .clk(clk),
    .d(csr_data[47]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b48  (
    .clk(clk),
    .d(csr_data[48]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b49  (
    .clk(clk),
    .d(csr_data[49]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b5  (
    .clk(clk),
    .d(csr_data[5]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b50  (
    .clk(clk),
    .d(csr_data[50]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b51  (
    .clk(clk),
    .d(csr_data[51]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b52  (
    .clk(clk),
    .d(csr_data[52]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b53  (
    .clk(clk),
    .d(csr_data[53]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b54  (
    .clk(clk),
    .d(csr_data[54]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b55  (
    .clk(clk),
    .d(csr_data[55]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b56  (
    .clk(clk),
    .d(csr_data[56]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b57  (
    .clk(clk),
    .d(csr_data[57]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b58  (
    .clk(clk),
    .d(csr_data[58]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b59  (
    .clk(clk),
    .d(csr_data[59]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b6  (
    .clk(clk),
    .d(csr_data[6]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b60  (
    .clk(clk),
    .d(csr_data[60]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b61  (
    .clk(clk),
    .d(csr_data[61]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b62  (
    .clk(clk),
    .d(csr_data[62]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b63  (
    .clk(clk),
    .d(csr_data[63]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b7  (
    .clk(clk),
    .d(csr_data[7]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b8  (
    .clk(clk),
    .d(csr_data[8]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg0_b9  (
    .clk(clk),
    .d(csr_data[9]),
    .en(\cu_ru/m_s_tvec/mux2_b0_sel_is_2_o ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/stvec [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b0  (
    .clk(clk),
    .d(csr_data[0]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [0]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b1  (
    .clk(clk),
    .d(csr_data[1]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [1]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b10  (
    .clk(clk),
    .d(csr_data[10]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [10]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b11  (
    .clk(clk),
    .d(csr_data[11]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [11]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b12  (
    .clk(clk),
    .d(csr_data[12]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [12]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b13  (
    .clk(clk),
    .d(csr_data[13]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [13]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b14  (
    .clk(clk),
    .d(csr_data[14]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [14]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b15  (
    .clk(clk),
    .d(csr_data[15]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [15]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b16  (
    .clk(clk),
    .d(csr_data[16]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [16]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b17  (
    .clk(clk),
    .d(csr_data[17]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [17]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b18  (
    .clk(clk),
    .d(csr_data[18]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [18]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b19  (
    .clk(clk),
    .d(csr_data[19]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [19]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b2  (
    .clk(clk),
    .d(csr_data[2]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [2]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b20  (
    .clk(clk),
    .d(csr_data[20]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [20]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b21  (
    .clk(clk),
    .d(csr_data[21]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [21]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b22  (
    .clk(clk),
    .d(csr_data[22]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [22]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b23  (
    .clk(clk),
    .d(csr_data[23]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [23]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b24  (
    .clk(clk),
    .d(csr_data[24]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [24]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b25  (
    .clk(clk),
    .d(csr_data[25]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [25]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b26  (
    .clk(clk),
    .d(csr_data[26]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [26]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b27  (
    .clk(clk),
    .d(csr_data[27]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [27]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b28  (
    .clk(clk),
    .d(csr_data[28]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [28]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b29  (
    .clk(clk),
    .d(csr_data[29]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [29]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b3  (
    .clk(clk),
    .d(csr_data[3]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [3]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b30  (
    .clk(clk),
    .d(csr_data[30]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [30]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b31  (
    .clk(clk),
    .d(csr_data[31]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [31]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b32  (
    .clk(clk),
    .d(csr_data[32]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [32]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b33  (
    .clk(clk),
    .d(csr_data[33]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [33]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b34  (
    .clk(clk),
    .d(csr_data[34]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [34]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b35  (
    .clk(clk),
    .d(csr_data[35]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [35]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b36  (
    .clk(clk),
    .d(csr_data[36]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [36]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b37  (
    .clk(clk),
    .d(csr_data[37]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [37]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b38  (
    .clk(clk),
    .d(csr_data[38]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [38]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b39  (
    .clk(clk),
    .d(csr_data[39]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [39]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b4  (
    .clk(clk),
    .d(csr_data[4]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [4]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b40  (
    .clk(clk),
    .d(csr_data[40]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [40]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b41  (
    .clk(clk),
    .d(csr_data[41]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [41]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b42  (
    .clk(clk),
    .d(csr_data[42]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [42]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b43  (
    .clk(clk),
    .d(csr_data[43]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [43]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b44  (
    .clk(clk),
    .d(csr_data[44]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [44]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b45  (
    .clk(clk),
    .d(csr_data[45]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [45]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b46  (
    .clk(clk),
    .d(csr_data[46]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [46]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b47  (
    .clk(clk),
    .d(csr_data[47]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [47]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b48  (
    .clk(clk),
    .d(csr_data[48]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [48]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b49  (
    .clk(clk),
    .d(csr_data[49]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [49]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b5  (
    .clk(clk),
    .d(csr_data[5]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [5]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b50  (
    .clk(clk),
    .d(csr_data[50]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [50]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b51  (
    .clk(clk),
    .d(csr_data[51]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [51]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b52  (
    .clk(clk),
    .d(csr_data[52]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [52]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b53  (
    .clk(clk),
    .d(csr_data[53]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [53]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b54  (
    .clk(clk),
    .d(csr_data[54]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [54]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b55  (
    .clk(clk),
    .d(csr_data[55]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [55]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b56  (
    .clk(clk),
    .d(csr_data[56]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [56]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b57  (
    .clk(clk),
    .d(csr_data[57]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [57]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b58  (
    .clk(clk),
    .d(csr_data[58]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [58]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b59  (
    .clk(clk),
    .d(csr_data[59]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [59]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b6  (
    .clk(clk),
    .d(csr_data[6]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [6]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b60  (
    .clk(clk),
    .d(csr_data[60]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [60]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b61  (
    .clk(clk),
    .d(csr_data[61]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [61]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b62  (
    .clk(clk),
    .d(csr_data[62]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [62]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b63  (
    .clk(clk),
    .d(csr_data[63]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [63]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b7  (
    .clk(clk),
    .d(csr_data[7]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [7]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b8  (
    .clk(clk),
    .d(csr_data[8]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [8]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  reg_sr_as_w1 \cu_ru/m_s_tvec/reg1_b9  (
    .clk(clk),
    .d(csr_data[9]),
    .en(\cu_ru/m_s_tvec/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mtvec [9]));  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(32)
  and \cu_ru/m_s_tvec/u1  (\cu_ru/m_s_tvec/n0 , \cu_ru/mrw_mtvec_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(26)
  and \cu_ru/m_s_tvec/u2  (\cu_ru/m_s_tvec/n1 , \cu_ru/srw_stvec_sel , wb_csr_write);  // ../../RTL/CPU/CU&RU/csrs/m_s_tvec.v(29)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dbk_reg  (
    .clk(clk),
    .d(data_csr[3]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [3]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/decs_reg  (
    .clk(clk),
    .d(data_csr[9]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [9]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/decu_reg  (
    .clk(clk),
    .d(data_csr[8]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [8]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/diaf_reg  (
    .clk(clk),
    .d(data_csr[1]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [1]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/diam_reg  (
    .clk(clk),
    .d(data_csr[0]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [0]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dii_reg  (
    .clk(clk),
    .d(data_csr[2]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [2]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dipf_reg  (
    .clk(clk),
    .d(data_csr[12]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [12]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dlaf_reg  (
    .clk(clk),
    .d(data_csr[5]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [5]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dlam_reg  (
    .clk(clk),
    .d(data_csr[4]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [4]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dlpf_reg  (
    .clk(clk),
    .d(data_csr[13]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [13]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dsaf_reg  (
    .clk(clk),
    .d(data_csr[7]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [7]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dsam_reg  (
    .clk(clk),
    .d(data_csr[6]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [6]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  reg_sr_as_w1 \cu_ru/medeleg_exc_ctrl/dspf_reg  (
    .clk(clk),
    .d(data_csr[15]),
    .en(\cu_ru/medeleg_exc_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/medeleg [15]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(133)
  binary_mux_s1_w1 \cu_ru/medeleg_exc_ctrl/mux10_b0  (
    .i0(\cu_ru/medeleg_exc_ctrl/n98 [0]),
    .i1(1'b0),
    .sel(\cu_ru/medeleg_exc_ctrl/n77 ),
    .o(\cu_ru/medeleg_exc_ctrl/n99 [0]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(176)
  and \cu_ru/medeleg_exc_ctrl/mux10_b1_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux10_b1_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n77_neg , \cu_ru/medeleg_exc_ctrl/mux9_b1_sel_is_0_o );
  not \cu_ru/medeleg_exc_ctrl/mux10_b1_sel_is_2_o_inv  (\cu_ru/medeleg_exc_ctrl/mux10_b1_sel_is_2_o_neg , \cu_ru/medeleg_exc_ctrl/mux10_b1_sel_is_2_o );
  binary_mux_s1_w1 \cu_ru/medeleg_exc_ctrl/mux10_b2  (
    .i0(\cu_ru/medeleg_exc_ctrl/n98 [2]),
    .i1(1'b1),
    .sel(\cu_ru/medeleg_exc_ctrl/n77 ),
    .o(\cu_ru/medeleg_exc_ctrl/n99 [2]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(176)
  and \cu_ru/medeleg_exc_ctrl/mux10_b3_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux10_b3_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n77_neg , \cu_ru/medeleg_exc_ctrl/mux9_b3_sel_is_2_o_neg );
  not \cu_ru/medeleg_exc_ctrl/mux10_b3_sel_is_0_o_inv  (\cu_ru/medeleg_exc_ctrl/mux10_b3_sel_is_0_o_neg , \cu_ru/medeleg_exc_ctrl/mux10_b3_sel_is_0_o );
  binary_mux_s1_w1 \cu_ru/medeleg_exc_ctrl/mux11_b0  (
    .i0(\cu_ru/medeleg_exc_ctrl/n99 [0]),
    .i1(1'b1),
    .sel(\cu_ru/medeleg_exc_ctrl/n76 ),
    .o(\cu_ru/exc_cause [0]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(176)
  AL_MUX \cu_ru/medeleg_exc_ctrl/mux11_b1  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\cu_ru/medeleg_exc_ctrl/mux11_b1_sel_is_0_o ),
    .o(\cu_ru/exc_cause [1]));
  and \cu_ru/medeleg_exc_ctrl/mux11_b1_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux11_b1_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n76_neg , \cu_ru/medeleg_exc_ctrl/mux10_b1_sel_is_2_o_neg );
  binary_mux_s1_w1 \cu_ru/medeleg_exc_ctrl/mux11_b2  (
    .i0(\cu_ru/medeleg_exc_ctrl/n99 [2]),
    .i1(1'b0),
    .sel(\cu_ru/medeleg_exc_ctrl/n76 ),
    .o(\cu_ru/exc_cause [2]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(176)
  AL_MUX \cu_ru/medeleg_exc_ctrl/mux11_b3  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\cu_ru/medeleg_exc_ctrl/mux11_b3_sel_is_0_o ),
    .o(\cu_ru/exc_cause [3]));
  and \cu_ru/medeleg_exc_ctrl/mux11_b3_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux11_b3_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n76_neg , \cu_ru/medeleg_exc_ctrl/mux10_b3_sel_is_0_o_neg );
  and \cu_ru/medeleg_exc_ctrl/mux1_b0_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux1_b0_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n86_neg , \cu_ru/medeleg_exc_ctrl/n87_neg );
  and \cu_ru/medeleg_exc_ctrl/mux1_b1_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux1_b1_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n86_neg , \cu_ru/medeleg_exc_ctrl/n87 );
  not \cu_ru/medeleg_exc_ctrl/mux1_b1_sel_is_2_o_inv  (\cu_ru/medeleg_exc_ctrl/mux1_b1_sel_is_2_o_neg , \cu_ru/medeleg_exc_ctrl/mux1_b1_sel_is_2_o );
  AL_MUX \cu_ru/medeleg_exc_ctrl/mux2_b0  (
    .i0(1'b1),
    .i1(\cu_ru/medeleg_exc_ctrl/n88 ),
    .sel(\cu_ru/medeleg_exc_ctrl/mux2_b0_sel_is_2_o ),
    .o(\cu_ru/medeleg_exc_ctrl/n91 [0]));
  and \cu_ru/medeleg_exc_ctrl/mux2_b0_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux2_b0_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n85_neg , \cu_ru/medeleg_exc_ctrl/mux1_b0_sel_is_0_o );
  and \cu_ru/medeleg_exc_ctrl/mux2_b1_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux2_b1_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n85_neg , \cu_ru/medeleg_exc_ctrl/mux1_b1_sel_is_2_o_neg );
  not \cu_ru/medeleg_exc_ctrl/mux2_b1_sel_is_0_o_inv  (\cu_ru/medeleg_exc_ctrl/mux2_b1_sel_is_0_o_neg , \cu_ru/medeleg_exc_ctrl/mux2_b1_sel_is_0_o );
  and \cu_ru/medeleg_exc_ctrl/mux2_b3_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux2_b3_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n85_neg , \cu_ru/medeleg_exc_ctrl/n86_neg );
  not \cu_ru/medeleg_exc_ctrl/mux2_b3_sel_is_0_o_inv  (\cu_ru/medeleg_exc_ctrl/mux2_b3_sel_is_0_o_neg , \cu_ru/medeleg_exc_ctrl/mux2_b3_sel_is_0_o );
  and \cu_ru/medeleg_exc_ctrl/mux3_b1_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux3_b1_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n84_neg , \cu_ru/medeleg_exc_ctrl/mux2_b1_sel_is_0_o_neg );
  not \cu_ru/medeleg_exc_ctrl/mux3_b1_sel_is_0_o_inv  (\cu_ru/medeleg_exc_ctrl/mux3_b1_sel_is_0_o_neg , \cu_ru/medeleg_exc_ctrl/mux3_b1_sel_is_0_o );
  and \cu_ru/medeleg_exc_ctrl/mux3_b3_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux3_b3_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n84_neg , \cu_ru/medeleg_exc_ctrl/mux2_b3_sel_is_0_o_neg );
  and \cu_ru/medeleg_exc_ctrl/mux4_b0_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux4_b0_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n83_neg , \cu_ru/medeleg_exc_ctrl/n84_neg );
  and \cu_ru/medeleg_exc_ctrl/mux4_b1_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux4_b1_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n83_neg , \cu_ru/medeleg_exc_ctrl/mux3_b1_sel_is_0_o_neg );
  not \cu_ru/medeleg_exc_ctrl/mux4_b1_sel_is_0_o_inv  (\cu_ru/medeleg_exc_ctrl/mux4_b1_sel_is_0_o_neg , \cu_ru/medeleg_exc_ctrl/mux4_b1_sel_is_0_o );
  AL_MUX \cu_ru/medeleg_exc_ctrl/mux4_b2  (
    .i0(1'b1),
    .i1(\cu_ru/medeleg_exc_ctrl/n91 [0]),
    .sel(\cu_ru/medeleg_exc_ctrl/mux4_b0_sel_is_0_o ),
    .o(\cu_ru/medeleg_exc_ctrl/n93 [2]));
  and \cu_ru/medeleg_exc_ctrl/mux4_b3_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux4_b3_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n83_neg , \cu_ru/medeleg_exc_ctrl/mux3_b3_sel_is_0_o );
  not \cu_ru/medeleg_exc_ctrl/mux4_b3_sel_is_2_o_inv  (\cu_ru/medeleg_exc_ctrl/mux4_b3_sel_is_2_o_neg , \cu_ru/medeleg_exc_ctrl/mux4_b3_sel_is_2_o );
  AL_MUX \cu_ru/medeleg_exc_ctrl/mux5_b0  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg_exc_ctrl/n91 [0]),
    .sel(\cu_ru/medeleg_exc_ctrl/mux5_b0_sel_is_2_o ),
    .o(\cu_ru/medeleg_exc_ctrl/n94 [0]));
  and \cu_ru/medeleg_exc_ctrl/mux5_b0_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux5_b0_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n82_neg , \cu_ru/medeleg_exc_ctrl/mux4_b0_sel_is_0_o );
  and \cu_ru/medeleg_exc_ctrl/mux5_b1_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux5_b1_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n82_neg , \cu_ru/medeleg_exc_ctrl/mux4_b1_sel_is_0_o_neg );
  and \cu_ru/medeleg_exc_ctrl/mux5_b3_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux5_b3_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n82_neg , \cu_ru/medeleg_exc_ctrl/mux4_b3_sel_is_2_o_neg );
  binary_mux_s1_w1 \cu_ru/medeleg_exc_ctrl/mux6_b0  (
    .i0(\cu_ru/medeleg_exc_ctrl/n94 [0]),
    .i1(1'b1),
    .sel(\cu_ru/medeleg_exc_ctrl/n81 ),
    .o(\cu_ru/medeleg_exc_ctrl/n95 [0]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(176)
  and \cu_ru/medeleg_exc_ctrl/mux6_b1_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux6_b1_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n81_neg , \cu_ru/medeleg_exc_ctrl/mux5_b1_sel_is_0_o );
  and \cu_ru/medeleg_exc_ctrl/mux6_b2_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux6_b2_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n81_neg , \cu_ru/medeleg_exc_ctrl/n82_neg );
  and \cu_ru/medeleg_exc_ctrl/mux6_b3_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux6_b3_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n81_neg , \cu_ru/medeleg_exc_ctrl/mux5_b3_sel_is_0_o );
  not \cu_ru/medeleg_exc_ctrl/mux6_b3_sel_is_2_o_inv  (\cu_ru/medeleg_exc_ctrl/mux6_b3_sel_is_2_o_neg , \cu_ru/medeleg_exc_ctrl/mux6_b3_sel_is_2_o );
  and \cu_ru/medeleg_exc_ctrl/mux7_b1_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux7_b1_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n80_neg , \cu_ru/medeleg_exc_ctrl/mux6_b1_sel_is_2_o );
  not \cu_ru/medeleg_exc_ctrl/mux7_b1_sel_is_2_o_inv  (\cu_ru/medeleg_exc_ctrl/mux7_b1_sel_is_2_o_neg , \cu_ru/medeleg_exc_ctrl/mux7_b1_sel_is_2_o );
  and \cu_ru/medeleg_exc_ctrl/mux7_b2_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux7_b2_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n80_neg , \cu_ru/medeleg_exc_ctrl/mux6_b2_sel_is_0_o );
  and \cu_ru/medeleg_exc_ctrl/mux7_b3_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux7_b3_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n80_neg , \cu_ru/medeleg_exc_ctrl/mux6_b3_sel_is_2_o_neg );
  AL_MUX \cu_ru/medeleg_exc_ctrl/mux8_b0  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg_exc_ctrl/n95 [0]),
    .sel(\cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o ),
    .o(\cu_ru/medeleg_exc_ctrl/n97 [0]));
  and \cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux8_b0_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n79_neg , \cu_ru/medeleg_exc_ctrl/n80_neg );
  and \cu_ru/medeleg_exc_ctrl/mux8_b1_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux8_b1_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n79_neg , \cu_ru/medeleg_exc_ctrl/mux7_b1_sel_is_2_o_neg );
  not \cu_ru/medeleg_exc_ctrl/mux8_b1_sel_is_0_o_inv  (\cu_ru/medeleg_exc_ctrl/mux8_b1_sel_is_0_o_neg , \cu_ru/medeleg_exc_ctrl/mux8_b1_sel_is_0_o );
  and \cu_ru/medeleg_exc_ctrl/mux8_b2_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux8_b2_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n79_neg , \cu_ru/medeleg_exc_ctrl/mux7_b2_sel_is_2_o );
  and \cu_ru/medeleg_exc_ctrl/mux8_b3_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux8_b3_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n79_neg , \cu_ru/medeleg_exc_ctrl/mux7_b3_sel_is_0_o );
  binary_mux_s1_w1 \cu_ru/medeleg_exc_ctrl/mux9_b0  (
    .i0(\cu_ru/medeleg_exc_ctrl/n97 [0]),
    .i1(1'b1),
    .sel(\cu_ru/medeleg_exc_ctrl/n78 ),
    .o(\cu_ru/medeleg_exc_ctrl/n98 [0]));  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(176)
  and \cu_ru/medeleg_exc_ctrl/mux9_b1_sel_is_0  (\cu_ru/medeleg_exc_ctrl/mux9_b1_sel_is_0_o , \cu_ru/medeleg_exc_ctrl/n78_neg , \cu_ru/medeleg_exc_ctrl/mux8_b1_sel_is_0_o_neg );
  AL_MUX \cu_ru/medeleg_exc_ctrl/mux9_b2  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg_exc_ctrl/n93 [2]),
    .sel(\cu_ru/medeleg_exc_ctrl/mux9_b2_sel_is_2_o ),
    .o(\cu_ru/medeleg_exc_ctrl/n98 [2]));
  and \cu_ru/medeleg_exc_ctrl/mux9_b2_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux9_b2_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n78_neg , \cu_ru/medeleg_exc_ctrl/mux8_b2_sel_is_2_o );
  and \cu_ru/medeleg_exc_ctrl/mux9_b3_sel_is_2  (\cu_ru/medeleg_exc_ctrl/mux9_b3_sel_is_2_o , \cu_ru/medeleg_exc_ctrl/n78_neg , \cu_ru/medeleg_exc_ctrl/mux8_b3_sel_is_2_o );
  not \cu_ru/medeleg_exc_ctrl/mux9_b3_sel_is_2_o_inv  (\cu_ru/medeleg_exc_ctrl/mux9_b3_sel_is_2_o_neg , \cu_ru/medeleg_exc_ctrl/mux9_b3_sel_is_2_o );
  not \cu_ru/medeleg_exc_ctrl/n76_inv  (\cu_ru/medeleg_exc_ctrl/n76_neg , \cu_ru/medeleg_exc_ctrl/n76 );
  not \cu_ru/medeleg_exc_ctrl/n77_inv  (\cu_ru/medeleg_exc_ctrl/n77_neg , \cu_ru/medeleg_exc_ctrl/n77 );
  not \cu_ru/medeleg_exc_ctrl/n78_inv  (\cu_ru/medeleg_exc_ctrl/n78_neg , \cu_ru/medeleg_exc_ctrl/n78 );
  not \cu_ru/medeleg_exc_ctrl/n79_inv  (\cu_ru/medeleg_exc_ctrl/n79_neg , \cu_ru/medeleg_exc_ctrl/n79 );
  not \cu_ru/medeleg_exc_ctrl/n80_inv  (\cu_ru/medeleg_exc_ctrl/n80_neg , \cu_ru/medeleg_exc_ctrl/n80 );
  not \cu_ru/medeleg_exc_ctrl/n81_inv  (\cu_ru/medeleg_exc_ctrl/n81_neg , \cu_ru/medeleg_exc_ctrl/n81 );
  not \cu_ru/medeleg_exc_ctrl/n82_inv  (\cu_ru/medeleg_exc_ctrl/n82_neg , \cu_ru/medeleg_exc_ctrl/n82 );
  not \cu_ru/medeleg_exc_ctrl/n83_inv  (\cu_ru/medeleg_exc_ctrl/n83_neg , \cu_ru/medeleg_exc_ctrl/n83 );
  not \cu_ru/medeleg_exc_ctrl/n84_inv  (\cu_ru/medeleg_exc_ctrl/n84_neg , \cu_ru/medeleg_exc_ctrl/n84 );
  not \cu_ru/medeleg_exc_ctrl/n85_inv  (\cu_ru/medeleg_exc_ctrl/n85_neg , \cu_ru/medeleg_exc_ctrl/n85 );
  not \cu_ru/medeleg_exc_ctrl/n86_inv  (\cu_ru/medeleg_exc_ctrl/n86_neg , \cu_ru/medeleg_exc_ctrl/n86 );
  not \cu_ru/medeleg_exc_ctrl/n87_inv  (\cu_ru/medeleg_exc_ctrl/n87_neg , \cu_ru/medeleg_exc_ctrl/n87 );
  and \cu_ru/medeleg_exc_ctrl/u100  (\cu_ru/medeleg_exc_ctrl/n70 , \cu_ru/medeleg_exc_ctrl/n64 , wb_ld_acc_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(154)
  and \cu_ru/medeleg_exc_ctrl/u101  (\cu_ru/medeleg_exc_ctrl/laf_target_s , \cu_ru/medeleg_exc_ctrl/n70 , \cu_ru/medeleg [5]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(154)
  and \cu_ru/medeleg_exc_ctrl/u103  (\cu_ru/medeleg_exc_ctrl/n71 , \cu_ru/medeleg_exc_ctrl/n64 , wb_st_addr_mis);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(155)
  and \cu_ru/medeleg_exc_ctrl/u104  (\cu_ru/medeleg_exc_ctrl/sam_target_s , \cu_ru/medeleg_exc_ctrl/n71 , \cu_ru/medeleg [6]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(155)
  and \cu_ru/medeleg_exc_ctrl/u106  (\cu_ru/medeleg_exc_ctrl/n72 , \cu_ru/medeleg_exc_ctrl/n64 , wb_st_acc_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(156)
  and \cu_ru/medeleg_exc_ctrl/u107  (\cu_ru/medeleg_exc_ctrl/saf_target_s , \cu_ru/medeleg_exc_ctrl/n72 , \cu_ru/medeleg [7]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(156)
  and \cu_ru/medeleg_exc_ctrl/u109  (\cu_ru/medeleg_exc_ctrl/ecu_target_s , \cu_ru/medeleg_exc_ctrl/n51 , \cu_ru/medeleg [8]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(157)
  and \cu_ru/medeleg_exc_ctrl/u111  (\cu_ru/medeleg_exc_ctrl/ecs_target_s , \cu_ru/medeleg_exc_ctrl/n53 , \cu_ru/medeleg [9]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(158)
  and \cu_ru/medeleg_exc_ctrl/u113  (\cu_ru/medeleg_exc_ctrl/n73 , \cu_ru/medeleg_exc_ctrl/n64 , wb_ins_page_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(159)
  and \cu_ru/medeleg_exc_ctrl/u114  (\cu_ru/medeleg_exc_ctrl/ipf_target_s , \cu_ru/medeleg_exc_ctrl/n73 , \cu_ru/medeleg [12]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(159)
  and \cu_ru/medeleg_exc_ctrl/u116  (\cu_ru/medeleg_exc_ctrl/n74 , \cu_ru/medeleg_exc_ctrl/n64 , wb_ld_page_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(160)
  and \cu_ru/medeleg_exc_ctrl/u117  (\cu_ru/medeleg_exc_ctrl/lpf_target_s , \cu_ru/medeleg_exc_ctrl/n74 , \cu_ru/medeleg [13]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(160)
  and \cu_ru/medeleg_exc_ctrl/u119  (\cu_ru/medeleg_exc_ctrl/n75 , \cu_ru/medeleg_exc_ctrl/n64 , wb_st_page_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(161)
  and \cu_ru/medeleg_exc_ctrl/u120  (\cu_ru/medeleg_exc_ctrl/spf_target_s , \cu_ru/medeleg_exc_ctrl/n75 , \cu_ru/medeleg [15]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(161)
  or \cu_ru/medeleg_exc_ctrl/u121  (\cu_ru/medeleg_exc_ctrl/n76 , \cu_ru/medeleg_exc_ctrl/bk_target_m , \cu_ru/medeleg_exc_ctrl/bk_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(164)
  or \cu_ru/medeleg_exc_ctrl/u122  (\cu_ru/medeleg_exc_ctrl/n77 , \cu_ru/medeleg_exc_ctrl/ipf_target_m , \cu_ru/medeleg_exc_ctrl/ipf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(165)
  or \cu_ru/medeleg_exc_ctrl/u123  (\cu_ru/medeleg_exc_ctrl/n78 , \cu_ru/medeleg_exc_ctrl/iaf_target_m , \cu_ru/medeleg_exc_ctrl/iaf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(166)
  or \cu_ru/medeleg_exc_ctrl/u124  (\cu_ru/medeleg_exc_ctrl/n79 , \cu_ru/medeleg_exc_ctrl/ii_target_m , \cu_ru/medeleg_exc_ctrl/ii_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(167)
  or \cu_ru/medeleg_exc_ctrl/u125  (\cu_ru/medeleg_exc_ctrl/n80 , \cu_ru/medeleg_exc_ctrl/iam_target_m , \cu_ru/medeleg_exc_ctrl/iam_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(168)
  or \cu_ru/medeleg_exc_ctrl/u126  (\cu_ru/medeleg_exc_ctrl/n81 , \cu_ru/medeleg_exc_ctrl/ecs_target_m , \cu_ru/medeleg_exc_ctrl/ecs_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(169)
  or \cu_ru/medeleg_exc_ctrl/u127  (\cu_ru/medeleg_exc_ctrl/n82 , \cu_ru/medeleg_exc_ctrl/ecu_target_m , \cu_ru/medeleg_exc_ctrl/ecu_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(170)
  or \cu_ru/medeleg_exc_ctrl/u128  (\cu_ru/medeleg_exc_ctrl/n83 , \cu_ru/medeleg_exc_ctrl/sam_target_m , \cu_ru/medeleg_exc_ctrl/sam_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(171)
  or \cu_ru/medeleg_exc_ctrl/u129  (\cu_ru/medeleg_exc_ctrl/n84 , \cu_ru/medeleg_exc_ctrl/lam_target_m , \cu_ru/medeleg_exc_ctrl/lam_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(172)
  or \cu_ru/medeleg_exc_ctrl/u130  (\cu_ru/medeleg_exc_ctrl/n85 , \cu_ru/medeleg_exc_ctrl/spf_target_m , \cu_ru/medeleg_exc_ctrl/spf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(173)
  or \cu_ru/medeleg_exc_ctrl/u131  (\cu_ru/medeleg_exc_ctrl/n86 , \cu_ru/medeleg_exc_ctrl/lpf_target_m , \cu_ru/medeleg_exc_ctrl/lpf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(174)
  or \cu_ru/medeleg_exc_ctrl/u132  (\cu_ru/medeleg_exc_ctrl/n87 , \cu_ru/medeleg_exc_ctrl/saf_target_m , \cu_ru/medeleg_exc_ctrl/saf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(175)
  or \cu_ru/medeleg_exc_ctrl/u133  (\cu_ru/medeleg_exc_ctrl/n88 , \cu_ru/medeleg_exc_ctrl/laf_target_m , \cu_ru/medeleg_exc_ctrl/laf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(176)
  or \cu_ru/medeleg_exc_ctrl/u196  (\cu_ru/medeleg_exc_ctrl/n100 , \cu_ru/medeleg_exc_ctrl/iam_target_m , \cu_ru/medeleg_exc_ctrl/iaf_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(181)
  or \cu_ru/medeleg_exc_ctrl/u197  (\cu_ru/medeleg_exc_ctrl/n101 , \cu_ru/medeleg_exc_ctrl/n100 , \cu_ru/medeleg_exc_ctrl/ii_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(181)
  or \cu_ru/medeleg_exc_ctrl/u198  (\cu_ru/medeleg_exc_ctrl/n102 , \cu_ru/medeleg_exc_ctrl/n101 , \cu_ru/medeleg_exc_ctrl/bk_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(181)
  or \cu_ru/medeleg_exc_ctrl/u199  (\cu_ru/medeleg_exc_ctrl/n103 , \cu_ru/medeleg_exc_ctrl/n102 , \cu_ru/medeleg_exc_ctrl/lam_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(181)
  or \cu_ru/medeleg_exc_ctrl/u200  (\cu_ru/medeleg_exc_ctrl/n104 , \cu_ru/medeleg_exc_ctrl/n103 , \cu_ru/medeleg_exc_ctrl/laf_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(181)
  or \cu_ru/medeleg_exc_ctrl/u201  (\cu_ru/medeleg_exc_ctrl/n105 , \cu_ru/medeleg_exc_ctrl/n104 , \cu_ru/medeleg_exc_ctrl/sam_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(181)
  or \cu_ru/medeleg_exc_ctrl/u202  (\cu_ru/medeleg_exc_ctrl/n106 , \cu_ru/medeleg_exc_ctrl/n105 , \cu_ru/medeleg_exc_ctrl/saf_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(181)
  or \cu_ru/medeleg_exc_ctrl/u203  (\cu_ru/medeleg_exc_ctrl/n107 , \cu_ru/medeleg_exc_ctrl/n106 , \cu_ru/medeleg_exc_ctrl/ecu_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(182)
  or \cu_ru/medeleg_exc_ctrl/u204  (\cu_ru/medeleg_exc_ctrl/n108 , \cu_ru/medeleg_exc_ctrl/n107 , \cu_ru/medeleg_exc_ctrl/ecs_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(182)
  or \cu_ru/medeleg_exc_ctrl/u205  (\cu_ru/medeleg_exc_ctrl/n109 , \cu_ru/medeleg_exc_ctrl/n108 , \cu_ru/medeleg_exc_ctrl/ipf_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(182)
  or \cu_ru/medeleg_exc_ctrl/u206  (\cu_ru/medeleg_exc_ctrl/n110 , \cu_ru/medeleg_exc_ctrl/n109 , \cu_ru/medeleg_exc_ctrl/lpf_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(182)
  or \cu_ru/medeleg_exc_ctrl/u207  (\cu_ru/medeleg_exc_ctrl/n111 , \cu_ru/medeleg_exc_ctrl/n110 , \cu_ru/medeleg_exc_ctrl/spf_target_m );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(182)
  and \cu_ru/medeleg_exc_ctrl/u208  (\cu_ru/exc_target_m , wb_valid, \cu_ru/medeleg_exc_ctrl/n111 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(182)
  or \cu_ru/medeleg_exc_ctrl/u209  (\cu_ru/medeleg_exc_ctrl/n112 , \cu_ru/medeleg_exc_ctrl/iam_target_s , \cu_ru/medeleg_exc_ctrl/iaf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(183)
  or \cu_ru/medeleg_exc_ctrl/u210  (\cu_ru/medeleg_exc_ctrl/n113 , \cu_ru/medeleg_exc_ctrl/n112 , \cu_ru/medeleg_exc_ctrl/ii_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(183)
  or \cu_ru/medeleg_exc_ctrl/u211  (\cu_ru/medeleg_exc_ctrl/n114 , \cu_ru/medeleg_exc_ctrl/n113 , \cu_ru/medeleg_exc_ctrl/bk_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(183)
  or \cu_ru/medeleg_exc_ctrl/u212  (\cu_ru/medeleg_exc_ctrl/n115 , \cu_ru/medeleg_exc_ctrl/n114 , \cu_ru/medeleg_exc_ctrl/lam_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(183)
  or \cu_ru/medeleg_exc_ctrl/u213  (\cu_ru/medeleg_exc_ctrl/n116 , \cu_ru/medeleg_exc_ctrl/n115 , \cu_ru/medeleg_exc_ctrl/laf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(183)
  or \cu_ru/medeleg_exc_ctrl/u214  (\cu_ru/medeleg_exc_ctrl/n117 , \cu_ru/medeleg_exc_ctrl/n116 , \cu_ru/medeleg_exc_ctrl/sam_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(183)
  or \cu_ru/medeleg_exc_ctrl/u215  (\cu_ru/medeleg_exc_ctrl/n118 , \cu_ru/medeleg_exc_ctrl/n117 , \cu_ru/medeleg_exc_ctrl/saf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(183)
  or \cu_ru/medeleg_exc_ctrl/u216  (\cu_ru/medeleg_exc_ctrl/n119 , \cu_ru/medeleg_exc_ctrl/n118 , \cu_ru/medeleg_exc_ctrl/ecu_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(184)
  or \cu_ru/medeleg_exc_ctrl/u217  (\cu_ru/medeleg_exc_ctrl/n120 , \cu_ru/medeleg_exc_ctrl/n119 , \cu_ru/medeleg_exc_ctrl/ecs_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(184)
  or \cu_ru/medeleg_exc_ctrl/u218  (\cu_ru/medeleg_exc_ctrl/n121 , \cu_ru/medeleg_exc_ctrl/n120 , \cu_ru/medeleg_exc_ctrl/ipf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(184)
  or \cu_ru/medeleg_exc_ctrl/u219  (\cu_ru/medeleg_exc_ctrl/n122 , \cu_ru/medeleg_exc_ctrl/n121 , \cu_ru/medeleg_exc_ctrl/lpf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(184)
  or \cu_ru/medeleg_exc_ctrl/u220  (\cu_ru/medeleg_exc_ctrl/n123 , \cu_ru/medeleg_exc_ctrl/n122 , \cu_ru/medeleg_exc_ctrl/spf_target_s );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(184)
  and \cu_ru/medeleg_exc_ctrl/u221  (\cu_ru/exc_target_s , wb_valid, \cu_ru/medeleg_exc_ctrl/n123 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(184)
  and \cu_ru/medeleg_exc_ctrl/u34  (\cu_ru/medeleg_exc_ctrl/n27 , priv[3], wb_ins_addr_mis);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(135)
  not \cu_ru/medeleg_exc_ctrl/u35  (\cu_ru/medeleg_exc_ctrl/n28 , \cu_ru/medeleg [0]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(135)
  and \cu_ru/medeleg_exc_ctrl/u36  (\cu_ru/medeleg_exc_ctrl/n29 , wb_ins_addr_mis, \cu_ru/medeleg_exc_ctrl/n28 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(135)
  or \cu_ru/medeleg_exc_ctrl/u37  (\cu_ru/medeleg_exc_ctrl/iam_target_m , \cu_ru/medeleg_exc_ctrl/n27 , \cu_ru/medeleg_exc_ctrl/n29 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(135)
  and \cu_ru/medeleg_exc_ctrl/u38  (\cu_ru/medeleg_exc_ctrl/n30 , priv[3], wb_ins_acc_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(136)
  not \cu_ru/medeleg_exc_ctrl/u39  (\cu_ru/medeleg_exc_ctrl/n31 , \cu_ru/medeleg [1]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(136)
  and \cu_ru/medeleg_exc_ctrl/u40  (\cu_ru/medeleg_exc_ctrl/n32 , wb_ins_acc_fault, \cu_ru/medeleg_exc_ctrl/n31 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(136)
  or \cu_ru/medeleg_exc_ctrl/u41  (\cu_ru/medeleg_exc_ctrl/iaf_target_m , \cu_ru/medeleg_exc_ctrl/n30 , \cu_ru/medeleg_exc_ctrl/n32 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(136)
  and \cu_ru/medeleg_exc_ctrl/u42  (\cu_ru/medeleg_exc_ctrl/n33 , priv[3], wb_ill_ins);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(137)
  not \cu_ru/medeleg_exc_ctrl/u43  (\cu_ru/medeleg_exc_ctrl/n34 , \cu_ru/medeleg [2]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(137)
  and \cu_ru/medeleg_exc_ctrl/u44  (\cu_ru/medeleg_exc_ctrl/n35 , wb_ill_ins, \cu_ru/medeleg_exc_ctrl/n34 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(137)
  or \cu_ru/medeleg_exc_ctrl/u45  (\cu_ru/medeleg_exc_ctrl/ii_target_m , \cu_ru/medeleg_exc_ctrl/n33 , \cu_ru/medeleg_exc_ctrl/n35 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(137)
  and \cu_ru/medeleg_exc_ctrl/u46  (\cu_ru/medeleg_exc_ctrl/n36 , priv[3], wb_ebreak);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(138)
  not \cu_ru/medeleg_exc_ctrl/u47  (\cu_ru/medeleg_exc_ctrl/n37 , \cu_ru/medeleg [3]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(138)
  and \cu_ru/medeleg_exc_ctrl/u48  (\cu_ru/medeleg_exc_ctrl/n38 , wb_ebreak, \cu_ru/medeleg_exc_ctrl/n37 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(138)
  or \cu_ru/medeleg_exc_ctrl/u49  (\cu_ru/medeleg_exc_ctrl/bk_target_m , \cu_ru/medeleg_exc_ctrl/n36 , \cu_ru/medeleg_exc_ctrl/n38 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(138)
  and \cu_ru/medeleg_exc_ctrl/u50  (\cu_ru/medeleg_exc_ctrl/n39 , priv[3], wb_ld_addr_mis);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(139)
  not \cu_ru/medeleg_exc_ctrl/u51  (\cu_ru/medeleg_exc_ctrl/n40 , \cu_ru/medeleg [4]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(139)
  and \cu_ru/medeleg_exc_ctrl/u52  (\cu_ru/medeleg_exc_ctrl/n41 , wb_ld_addr_mis, \cu_ru/medeleg_exc_ctrl/n40 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(139)
  or \cu_ru/medeleg_exc_ctrl/u53  (\cu_ru/medeleg_exc_ctrl/lam_target_m , \cu_ru/medeleg_exc_ctrl/n39 , \cu_ru/medeleg_exc_ctrl/n41 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(139)
  and \cu_ru/medeleg_exc_ctrl/u54  (\cu_ru/medeleg_exc_ctrl/n42 , priv[3], wb_ld_acc_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(140)
  not \cu_ru/medeleg_exc_ctrl/u55  (\cu_ru/medeleg_exc_ctrl/n43 , \cu_ru/medeleg [5]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(140)
  and \cu_ru/medeleg_exc_ctrl/u56  (\cu_ru/medeleg_exc_ctrl/n44 , wb_ld_acc_fault, \cu_ru/medeleg_exc_ctrl/n43 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(140)
  or \cu_ru/medeleg_exc_ctrl/u57  (\cu_ru/medeleg_exc_ctrl/laf_target_m , \cu_ru/medeleg_exc_ctrl/n42 , \cu_ru/medeleg_exc_ctrl/n44 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(140)
  and \cu_ru/medeleg_exc_ctrl/u58  (\cu_ru/medeleg_exc_ctrl/n45 , priv[3], wb_st_addr_mis);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(141)
  not \cu_ru/medeleg_exc_ctrl/u59  (\cu_ru/medeleg_exc_ctrl/n46 , \cu_ru/medeleg [6]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(141)
  and \cu_ru/medeleg_exc_ctrl/u60  (\cu_ru/medeleg_exc_ctrl/n47 , wb_st_addr_mis, \cu_ru/medeleg_exc_ctrl/n46 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(141)
  or \cu_ru/medeleg_exc_ctrl/u61  (\cu_ru/medeleg_exc_ctrl/sam_target_m , \cu_ru/medeleg_exc_ctrl/n45 , \cu_ru/medeleg_exc_ctrl/n47 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(141)
  and \cu_ru/medeleg_exc_ctrl/u62  (\cu_ru/medeleg_exc_ctrl/n48 , priv[3], wb_st_acc_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(142)
  not \cu_ru/medeleg_exc_ctrl/u63  (\cu_ru/medeleg_exc_ctrl/n49 , \cu_ru/medeleg [7]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(142)
  and \cu_ru/medeleg_exc_ctrl/u64  (\cu_ru/medeleg_exc_ctrl/n50 , wb_st_acc_fault, \cu_ru/medeleg_exc_ctrl/n49 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(142)
  or \cu_ru/medeleg_exc_ctrl/u65  (\cu_ru/medeleg_exc_ctrl/saf_target_m , \cu_ru/medeleg_exc_ctrl/n48 , \cu_ru/medeleg_exc_ctrl/n50 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(142)
  and \cu_ru/medeleg_exc_ctrl/u66  (\cu_ru/medeleg_exc_ctrl/n51 , priv[0], wb_ecall);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(143)
  not \cu_ru/medeleg_exc_ctrl/u67  (\cu_ru/medeleg_exc_ctrl/n52 , \cu_ru/medeleg [8]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(143)
  and \cu_ru/medeleg_exc_ctrl/u68  (\cu_ru/medeleg_exc_ctrl/ecu_target_m , \cu_ru/medeleg_exc_ctrl/n51 , \cu_ru/medeleg_exc_ctrl/n52 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(143)
  and \cu_ru/medeleg_exc_ctrl/u69  (\cu_ru/medeleg_exc_ctrl/n53 , priv[1], wb_ecall);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(144)
  and \cu_ru/medeleg_exc_ctrl/u7  (\cu_ru/medeleg_exc_ctrl/n0 , wb_csr_write, \cu_ru/mrw_medeleg_sel );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(118)
  not \cu_ru/medeleg_exc_ctrl/u70  (\cu_ru/medeleg_exc_ctrl/n54 , \cu_ru/medeleg [9]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(144)
  and \cu_ru/medeleg_exc_ctrl/u71  (\cu_ru/medeleg_exc_ctrl/ecs_target_m , \cu_ru/medeleg_exc_ctrl/n53 , \cu_ru/medeleg_exc_ctrl/n54 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(144)
  and \cu_ru/medeleg_exc_ctrl/u72  (\cu_ru/medeleg_exc_ctrl/n55 , priv[3], wb_ins_page_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(145)
  not \cu_ru/medeleg_exc_ctrl/u73  (\cu_ru/medeleg_exc_ctrl/n56 , \cu_ru/medeleg [12]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(145)
  and \cu_ru/medeleg_exc_ctrl/u74  (\cu_ru/medeleg_exc_ctrl/n57 , wb_ins_page_fault, \cu_ru/medeleg_exc_ctrl/n56 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(145)
  or \cu_ru/medeleg_exc_ctrl/u75  (\cu_ru/medeleg_exc_ctrl/ipf_target_m , \cu_ru/medeleg_exc_ctrl/n55 , \cu_ru/medeleg_exc_ctrl/n57 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(145)
  and \cu_ru/medeleg_exc_ctrl/u76  (\cu_ru/medeleg_exc_ctrl/n58 , priv[3], wb_ld_page_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(146)
  not \cu_ru/medeleg_exc_ctrl/u77  (\cu_ru/medeleg_exc_ctrl/n59 , \cu_ru/medeleg [13]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(146)
  and \cu_ru/medeleg_exc_ctrl/u78  (\cu_ru/medeleg_exc_ctrl/n60 , wb_ld_page_fault, \cu_ru/medeleg_exc_ctrl/n59 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(146)
  or \cu_ru/medeleg_exc_ctrl/u79  (\cu_ru/medeleg_exc_ctrl/lpf_target_m , \cu_ru/medeleg_exc_ctrl/n58 , \cu_ru/medeleg_exc_ctrl/n60 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(146)
  and \cu_ru/medeleg_exc_ctrl/u80  (\cu_ru/medeleg_exc_ctrl/n61 , priv[3], wb_st_page_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(147)
  not \cu_ru/medeleg_exc_ctrl/u81  (\cu_ru/medeleg_exc_ctrl/n62 , \cu_ru/medeleg [15]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(147)
  and \cu_ru/medeleg_exc_ctrl/u82  (\cu_ru/medeleg_exc_ctrl/n63 , wb_st_page_fault, \cu_ru/medeleg_exc_ctrl/n62 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(147)
  or \cu_ru/medeleg_exc_ctrl/u83  (\cu_ru/medeleg_exc_ctrl/spf_target_m , \cu_ru/medeleg_exc_ctrl/n61 , \cu_ru/medeleg_exc_ctrl/n63 );  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(147)
  or \cu_ru/medeleg_exc_ctrl/u84  (\cu_ru/medeleg_exc_ctrl/n64 , priv[1], priv[0]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(149)
  and \cu_ru/medeleg_exc_ctrl/u85  (\cu_ru/medeleg_exc_ctrl/n65 , \cu_ru/medeleg_exc_ctrl/n64 , wb_ins_addr_mis);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(149)
  and \cu_ru/medeleg_exc_ctrl/u86  (\cu_ru/medeleg_exc_ctrl/iam_target_s , \cu_ru/medeleg_exc_ctrl/n65 , \cu_ru/medeleg [0]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(149)
  and \cu_ru/medeleg_exc_ctrl/u88  (\cu_ru/medeleg_exc_ctrl/n66 , \cu_ru/medeleg_exc_ctrl/n64 , wb_ins_acc_fault);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(150)
  and \cu_ru/medeleg_exc_ctrl/u89  (\cu_ru/medeleg_exc_ctrl/iaf_target_s , \cu_ru/medeleg_exc_ctrl/n66 , \cu_ru/medeleg [1]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(150)
  and \cu_ru/medeleg_exc_ctrl/u91  (\cu_ru/medeleg_exc_ctrl/n67 , \cu_ru/medeleg_exc_ctrl/n64 , wb_ill_ins);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(151)
  and \cu_ru/medeleg_exc_ctrl/u92  (\cu_ru/medeleg_exc_ctrl/ii_target_s , \cu_ru/medeleg_exc_ctrl/n67 , \cu_ru/medeleg [2]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(151)
  and \cu_ru/medeleg_exc_ctrl/u94  (\cu_ru/medeleg_exc_ctrl/n68 , \cu_ru/medeleg_exc_ctrl/n64 , wb_ebreak);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(152)
  and \cu_ru/medeleg_exc_ctrl/u95  (\cu_ru/medeleg_exc_ctrl/bk_target_s , \cu_ru/medeleg_exc_ctrl/n68 , \cu_ru/medeleg [3]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(152)
  and \cu_ru/medeleg_exc_ctrl/u97  (\cu_ru/medeleg_exc_ctrl/n69 , \cu_ru/medeleg_exc_ctrl/n64 , wb_ld_addr_mis);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(153)
  and \cu_ru/medeleg_exc_ctrl/u98  (\cu_ru/medeleg_exc_ctrl/lam_target_s , \cu_ru/medeleg_exc_ctrl/n69 , \cu_ru/medeleg [4]);  // ../../RTL/CPU/CU&RU/csrs/medeleg_exc_ctrl.v(153)
  reg_sr_as_w1 \cu_ru/mideleg_int_ctrl/dsei_reg  (
    .clk(clk),
    .d(data_csr[9]),
    .en(\cu_ru/mideleg_int_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mideleg [9]));  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  reg_sr_as_w1 \cu_ru/mideleg_int_ctrl/dssi_reg  (
    .clk(clk),
    .d(data_csr[1]),
    .en(\cu_ru/mideleg_int_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mideleg [1]));  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  reg_sr_as_w1 \cu_ru/mideleg_int_ctrl/dsti_reg  (
    .clk(clk),
    .d(data_csr[5]),
    .en(\cu_ru/mideleg_int_ctrl/n0 ),
    .reset(rst),
    .set(1'b0),
    .q(\cu_ru/mideleg [5]));  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(81)
  not \cu_ru/mideleg_int_ctrl/mei_ack_m_inv  (\cu_ru/mideleg_int_ctrl/mei_ack_m_neg , \cu_ru/mideleg_int_ctrl/mei_ack_m );
  not \cu_ru/mideleg_int_ctrl/msi_ack_m_inv  (\cu_ru/mideleg_int_ctrl/msi_ack_m_neg , \cu_ru/mideleg_int_ctrl/msi_ack_m );
  not \cu_ru/mideleg_int_ctrl/mti_ack_m_inv  (\cu_ru/mideleg_int_ctrl/mti_ack_m_neg , \cu_ru/mideleg_int_ctrl/mti_ack_m );
  and \cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0  (\cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o , \cu_ru/mideleg_int_ctrl/n33_neg , \cu_ru/mideleg_int_ctrl/n34_neg );
  AL_MUX \cu_ru/mideleg_int_ctrl/mux1_b2  (
    .i0(1'b0),
    .i1(\cu_ru/mideleg_int_ctrl/n35 ),
    .sel(\cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o ),
    .o(\cu_ru/mideleg_int_ctrl/n37 [2]));
  and \cu_ru/mideleg_int_ctrl/mux2_b0_sel_is_2  (\cu_ru/mideleg_int_ctrl/mux2_b0_sel_is_2_o , \cu_ru/mideleg_int_ctrl/mti_ack_m_neg , \cu_ru/mideleg_int_ctrl/mux1_b0_sel_is_0_o );
  binary_mux_s1_w1 \cu_ru/mideleg_int_ctrl/mux2_b2  (
    .i0(\cu_ru/mideleg_int_ctrl/n37 [2]),
    .i1(1'b1),
    .sel(\cu_ru/mideleg_int_ctrl/mti_ack_m ),
    .o(\cu_ru/mideleg_int_ctrl/n38 [2]));  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(105)
  and \cu_ru/mideleg_int_ctrl/mux2_b3_sel_is_2  (\cu_ru/mideleg_int_ctrl/mux2_b3_sel_is_2_o , \cu_ru/mideleg_int_ctrl/mti_ack_m_neg , \cu_ru/mideleg_int_ctrl/n33 );
  and \cu_ru/mideleg_int_ctrl/mux3_b0_sel_is_2  (\cu_ru/mideleg_int_ctrl/mux3_b0_sel_is_2_o , \cu_ru/mideleg_int_ctrl/msi_ack_m_neg , \cu_ru/mideleg_int_ctrl/mux2_b0_sel_is_2_o );
  and \cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0  (\cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o , \cu_ru/mideleg_int_ctrl/msi_ack_m_neg , \cu_ru/mideleg_int_ctrl/mti_ack_m_neg );
  and \cu_ru/mideleg_int_ctrl/mux3_b3_sel_is_2  (\cu_ru/mideleg_int_ctrl/mux3_b3_sel_is_2_o , \cu_ru/mideleg_int_ctrl/msi_ack_m_neg , \cu_ru/mideleg_int_ctrl/mux2_b3_sel_is_2_o );
  not \cu_ru/mideleg_int_ctrl/mux3_b3_sel_is_2_o_inv  (\cu_ru/mideleg_int_ctrl/mux3_b3_sel_is_2_o_neg , \cu_ru/mideleg_int_ctrl/mux3_b3_sel_is_2_o );
  AL_MUX \cu_ru/mideleg_int_ctrl/mux4_b0  (
    .i0(1'b1),
    .i1(\cu_ru/mideleg_int_ctrl/n35 ),
    .sel(\cu_ru/mideleg_int_ctrl/mux4_b0_sel_is_2_o ),
    .o(\cu_ru/int_cause [63]));
  and \cu_ru/mideleg_int_ctrl/mux4_b0_sel_is_2  (\cu_ru/mideleg_int_ctrl/mux4_b0_sel_is_2_o , \cu_ru/mideleg_int_ctrl/mei_ack_m_neg , \cu_ru/mideleg_int_ctrl/mux3_b0_sel_is_2_o );
  AL_MUX \cu_ru/mideleg_int_ctrl/mux4_b1  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\cu_ru/mideleg_int_ctrl/mux4_b1_sel_is_2_o ),
    .o(\cu_ru/int_cause [1]));
  and \cu_ru/mideleg_int_ctrl/mux4_b1_sel_is_2  (\cu_ru/mideleg_int_ctrl/mux4_b1_sel_is_2_o , \cu_ru/mideleg_int_ctrl/mei_ack_m_neg , \cu_ru/mideleg_int_ctrl/mux3_b1_sel_is_0_o );
  AL_MUX \cu_ru/mideleg_int_ctrl/mux4_b2  (
    .i0(1'b0),
    .i1(\cu_ru/mideleg_int_ctrl/n38 [2]),
    .sel(\cu_ru/mideleg_int_ctrl/mux4_b2_sel_is_0_o ),
    .o(\cu_ru/int_cause [2]));
  and \cu_ru/mideleg_int_ctrl/mux4_b2_sel_is_0  (\cu_ru/mideleg_int_ctrl/mux4_b2_sel_is_0_o , \cu_ru/mideleg_int_ctrl/mei_ack_m_neg , \cu_ru/mideleg_int_ctrl/msi_ack_m_neg );
  AL_MUX \cu_ru/mideleg_int_ctrl/mux4_b3  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\cu_ru/mideleg_int_ctrl/mux4_b3_sel_is_0_o ),
    .o(\cu_ru/int_cause [3]));
  and \cu_ru/mideleg_int_ctrl/mux4_b3_sel_is_0  (\cu_ru/mideleg_int_ctrl/mux4_b3_sel_is_0_o , \cu_ru/mideleg_int_ctrl/mei_ack_m_neg , \cu_ru/mideleg_int_ctrl/mux3_b3_sel_is_2_o_neg );
  not \cu_ru/mideleg_int_ctrl/n33_inv  (\cu_ru/mideleg_int_ctrl/n33_neg , \cu_ru/mideleg_int_ctrl/n33 );
  not \cu_ru/mideleg_int_ctrl/n34_inv  (\cu_ru/mideleg_int_ctrl/n34_neg , \cu_ru/mideleg_int_ctrl/n34 );
  and \cu_ru/mideleg_int_ctrl/u12  (\cu_ru/mideleg_int_ctrl/n7 , \cu_ru/mie , \cu_ru/m_sip [11]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(84)
  and \cu_ru/mideleg_int_ctrl/u13  (\cu_ru/mideleg_int_ctrl/mei_ack_m , \cu_ru/mideleg_int_ctrl/n7 , \cu_ru/m_sie [11]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(84)
  and \cu_ru/mideleg_int_ctrl/u14  (\cu_ru/mideleg_int_ctrl/n8 , \cu_ru/mie , \cu_ru/m_sip [3]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(85)
  and \cu_ru/mideleg_int_ctrl/u15  (\cu_ru/mideleg_int_ctrl/msi_ack_m , \cu_ru/mideleg_int_ctrl/n8 , \cu_ru/m_sie [3]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(85)
  and \cu_ru/mideleg_int_ctrl/u16  (\cu_ru/mideleg_int_ctrl/n9 , \cu_ru/mie , \cu_ru/m_sip [7]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(86)
  and \cu_ru/mideleg_int_ctrl/u17  (\cu_ru/mideleg_int_ctrl/mti_ack_m , \cu_ru/mideleg_int_ctrl/n9 , \cu_ru/m_sie [7]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(86)
  not \cu_ru/mideleg_int_ctrl/u18  (\cu_ru/mideleg_int_ctrl/n10 , \cu_ru/mideleg [9]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(87)
  and \cu_ru/mideleg_int_ctrl/u19  (\cu_ru/mideleg_int_ctrl/n11 , \cu_ru/mie , \cu_ru/mideleg_int_ctrl/n10 );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(87)
  or \cu_ru/mideleg_int_ctrl/u20  (\cu_ru/mideleg_int_ctrl/n12 , \cu_ru/m_sip [9], s_ext_int);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(87)
  and \cu_ru/mideleg_int_ctrl/u21  (\cu_ru/mideleg_int_ctrl/sei_ack_m , \cu_ru/mideleg_int_ctrl/n11 , \cu_ru/mideleg_int_ctrl/n12 );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(87)
  not \cu_ru/mideleg_int_ctrl/u22  (\cu_ru/mideleg_int_ctrl/n13 , \cu_ru/mideleg [1]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(88)
  and \cu_ru/mideleg_int_ctrl/u23  (\cu_ru/mideleg_int_ctrl/n14 , \cu_ru/mie , \cu_ru/mideleg_int_ctrl/n13 );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(88)
  and \cu_ru/mideleg_int_ctrl/u24  (\cu_ru/mideleg_int_ctrl/ssi_ack_m , \cu_ru/mideleg_int_ctrl/n14 , \cu_ru/m_sip [1]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(88)
  not \cu_ru/mideleg_int_ctrl/u25  (\cu_ru/mideleg_int_ctrl/n15 , \cu_ru/mideleg [5]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(89)
  and \cu_ru/mideleg_int_ctrl/u26  (\cu_ru/mideleg_int_ctrl/n16 , \cu_ru/mie , \cu_ru/mideleg_int_ctrl/n15 );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(89)
  and \cu_ru/mideleg_int_ctrl/u27  (\cu_ru/mideleg_int_ctrl/sti_ack_m , \cu_ru/mideleg_int_ctrl/n16 , \cu_ru/m_sip [5]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(89)
  and \cu_ru/mideleg_int_ctrl/u29  (\cu_ru/mideleg_int_ctrl/n18 , \cu_ru/mstatus [1], \cu_ru/medeleg_exc_ctrl/n64 );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(91)
  and \cu_ru/mideleg_int_ctrl/u31  (\cu_ru/mideleg_int_ctrl/n19 , \cu_ru/mideleg_int_ctrl/n18 , \cu_ru/mideleg_int_ctrl/n12 );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(91)
  and \cu_ru/mideleg_int_ctrl/u32  (\cu_ru/mideleg_int_ctrl/n20 , \cu_ru/mideleg_int_ctrl/n19 , \cu_ru/m_sie [9]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(91)
  and \cu_ru/mideleg_int_ctrl/u33  (\cu_ru/mideleg_int_ctrl/sei_ack_s , \cu_ru/mideleg_int_ctrl/n20 , \cu_ru/mideleg [9]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(91)
  and \cu_ru/mideleg_int_ctrl/u36  (\cu_ru/mideleg_int_ctrl/n21 , \cu_ru/mideleg_int_ctrl/n18 , \cu_ru/m_sip [1]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(92)
  and \cu_ru/mideleg_int_ctrl/u37  (\cu_ru/mideleg_int_ctrl/n22 , \cu_ru/mideleg_int_ctrl/n21 , \cu_ru/m_sie [1]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(92)
  and \cu_ru/mideleg_int_ctrl/u38  (\cu_ru/mideleg_int_ctrl/ssi_ack_s , \cu_ru/mideleg_int_ctrl/n22 , \cu_ru/mideleg [1]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(92)
  and \cu_ru/mideleg_int_ctrl/u4  (\cu_ru/mideleg_int_ctrl/n0 , wb_csr_write, \cu_ru/mrw_mideleg_sel );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(76)
  and \cu_ru/mideleg_int_ctrl/u41  (\cu_ru/mideleg_int_ctrl/n23 , \cu_ru/mideleg_int_ctrl/n18 , \cu_ru/m_sip [5]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(93)
  and \cu_ru/mideleg_int_ctrl/u42  (\cu_ru/mideleg_int_ctrl/n24 , \cu_ru/mideleg_int_ctrl/n23 , \cu_ru/m_sie [5]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(93)
  and \cu_ru/mideleg_int_ctrl/u43  (\cu_ru/mideleg_int_ctrl/sti_ack_s , \cu_ru/mideleg_int_ctrl/n24 , \cu_ru/mideleg [5]);  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(93)
  or \cu_ru/mideleg_int_ctrl/u47  (\cu_ru/mideleg_int_ctrl/n25 , \cu_ru/mideleg_int_ctrl/msi_ack_m , \cu_ru/mideleg_int_ctrl/mti_ack_m );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(100)
  or \cu_ru/mideleg_int_ctrl/u48  (\cu_ru/mideleg_int_ctrl/n26 , \cu_ru/mideleg_int_ctrl/n25 , \cu_ru/mideleg_int_ctrl/sei_ack_m );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(100)
  or \cu_ru/mideleg_int_ctrl/u49  (\cu_ru/mideleg_int_ctrl/n27 , \cu_ru/mideleg_int_ctrl/n26 , \cu_ru/mideleg_int_ctrl/ssi_ack_m );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(100)
  or \cu_ru/mideleg_int_ctrl/u50  (\cu_ru/int_target_m , \cu_ru/mideleg_int_ctrl/n27 , \cu_ru/mideleg_int_ctrl/sti_ack_m );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(100)
  not \cu_ru/mideleg_int_ctrl/u51  (\cu_ru/mideleg_int_ctrl/n28 , \cu_ru/int_target_m );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(101)
  or \cu_ru/mideleg_int_ctrl/u52  (\cu_ru/mideleg_int_ctrl/n29 , \cu_ru/mideleg_int_ctrl/sei_ack_s , \cu_ru/mideleg_int_ctrl/ssi_ack_s );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(101)
  or \cu_ru/mideleg_int_ctrl/u53  (\cu_ru/mideleg_int_ctrl/n30 , \cu_ru/mideleg_int_ctrl/n29 , \cu_ru/mideleg_int_ctrl/sti_ack_s );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(101)
  and \cu_ru/mideleg_int_ctrl/u54  (\cu_ru/int_target_s , \cu_ru/mideleg_int_ctrl/n28 , \cu_ru/mideleg_int_ctrl/n30 );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(101)
  or \cu_ru/mideleg_int_ctrl/u59  (\cu_ru/mideleg_int_ctrl/n31 , \cu_ru/int_target_m , \cu_ru/mideleg_int_ctrl/sei_ack_s );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(103)
  or \cu_ru/mideleg_int_ctrl/u60  (\cu_ru/mideleg_int_ctrl/n32 , \cu_ru/mideleg_int_ctrl/n31 , \cu_ru/mideleg_int_ctrl/ssi_ack_s );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(103)
  or \cu_ru/mideleg_int_ctrl/u61  (int_req, \cu_ru/mideleg_int_ctrl/n32 , \cu_ru/mideleg_int_ctrl/sti_ack_s );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(103)
  or \cu_ru/mideleg_int_ctrl/u62  (\cu_ru/mideleg_int_ctrl/n33 , \cu_ru/mideleg_int_ctrl/sei_ack_m , \cu_ru/mideleg_int_ctrl/sei_ack_s );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(105)
  or \cu_ru/mideleg_int_ctrl/u63  (\cu_ru/mideleg_int_ctrl/n34 , \cu_ru/mideleg_int_ctrl/ssi_ack_m , \cu_ru/mideleg_int_ctrl/ssi_ack_s );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(105)
  or \cu_ru/mideleg_int_ctrl/u64  (\cu_ru/mideleg_int_ctrl/n35 , \cu_ru/mideleg_int_ctrl/sti_ack_m , \cu_ru/mideleg_int_ctrl/sti_ack_s );  // ../../RTL/CPU/CU&RU/csrs/mideleg_int_ctrl.v(105)
  binary_mux_s1_w1 \cu_ru/mux0_b0  (
    .i0(\cu_ru/int_cause [63]),
    .i1(\cu_ru/exc_cause [0]),
    .sel(\cu_ru/exception ),
    .o(\cu_ru/trap_cause [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(350)
  binary_mux_s1_w1 \cu_ru/mux0_b1  (
    .i0(\cu_ru/int_cause [1]),
    .i1(\cu_ru/exc_cause [1]),
    .sel(\cu_ru/exception ),
    .o(\cu_ru/trap_cause [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(350)
  binary_mux_s1_w1 \cu_ru/mux0_b2  (
    .i0(\cu_ru/int_cause [2]),
    .i1(\cu_ru/exc_cause [2]),
    .sel(\cu_ru/exception ),
    .o(\cu_ru/trap_cause [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(350)
  binary_mux_s1_w1 \cu_ru/mux0_b3  (
    .i0(\cu_ru/int_cause [3]),
    .i1(\cu_ru/exc_cause [3]),
    .sel(\cu_ru/exception ),
    .o(\cu_ru/trap_cause [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(350)
  binary_mux_s1_w1 \cu_ru/mux0_b63  (
    .i0(\cu_ru/int_cause [63]),
    .i1(1'b0),
    .sel(\cu_ru/exception ),
    .o(\cu_ru/trap_cause [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(350)
  binary_mux_s1_w1 \cu_ru/mux10_b1  (
    .i0(1'b0),
    .i1(\cu_ru/mstatus [1]),
    .sel(\cu_ru/read_sstatus_sel ),
    .o(\cu_ru/n64 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  binary_mux_s1_w1 \cu_ru/mux10_b18  (
    .i0(1'b0),
    .i1(sum),
    .sel(\cu_ru/read_sstatus_sel ),
    .o(\cu_ru/n64 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  binary_mux_s1_w1 \cu_ru/mux10_b19  (
    .i0(1'b0),
    .i1(mxr),
    .sel(\cu_ru/read_sstatus_sel ),
    .o(\cu_ru/n64 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  binary_mux_s1_w1 \cu_ru/mux10_b32  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\cu_ru/read_sstatus_sel ),
    .o(\cu_ru/n64 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  binary_mux_s1_w1 \cu_ru/mux10_b5  (
    .i0(1'b0),
    .i1(\cu_ru/mstatus [5]),
    .sel(\cu_ru/read_sstatus_sel ),
    .o(\cu_ru/n64 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  binary_mux_s1_w1 \cu_ru/mux10_b8  (
    .i0(1'b0),
    .i1(\cu_ru/mstatus [8]),
    .sel(\cu_ru/read_sstatus_sel ),
    .o(\cu_ru/n64 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  binary_mux_s1_w1 \cu_ru/mux11_b0  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [0]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b1  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [1]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b10  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [10]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b11  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [11]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b12  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [12]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b13  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [13]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b14  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [14]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b15  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [15]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b16  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [16]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b17  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [17]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b18  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [18]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b19  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [19]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b2  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [2]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b20  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [20]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b21  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [21]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b22  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [22]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b23  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [23]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b24  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [24]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b25  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [25]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b26  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [26]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b27  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [27]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b28  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [28]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b29  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [29]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b3  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [3]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b30  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [30]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b31  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [31]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b32  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [32]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b33  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [33]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b34  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [34]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b35  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [35]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b36  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [36]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b37  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [37]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b38  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [38]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b39  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [39]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b4  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [4]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b40  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [40]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b41  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [41]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b42  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [42]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b43  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [43]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b44  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [44]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b45  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [45]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b46  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [46]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b47  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [47]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b48  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [48]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b49  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [49]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b5  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [5]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b50  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [50]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b51  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [51]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b52  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [52]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b53  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [53]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b54  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [54]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b55  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [55]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b56  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [56]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b57  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [57]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b58  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [58]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b59  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [59]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b6  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [6]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b60  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [60]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b61  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [61]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b62  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [62]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b63  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [63]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b7  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [7]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b8  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [8]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux11_b9  (
    .i0(1'b0),
    .i1(\cu_ru/stvec [9]),
    .sel(\cu_ru/read_stvec_sel ),
    .o(\cu_ru/n68 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  binary_mux_s1_w1 \cu_ru/mux12_b0  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [0]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b1  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [1]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b10  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [10]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b11  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [11]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b12  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [12]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b13  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [13]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b14  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [14]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b15  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [15]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b16  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [16]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b17  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [17]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b18  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [18]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b19  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [19]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b2  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [2]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b20  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [20]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b21  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [21]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b22  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [22]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b23  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [23]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b24  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [24]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b25  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [25]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b26  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [26]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b27  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [27]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b28  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [28]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b29  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [29]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b3  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [3]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b30  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [30]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b31  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [31]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b32  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [32]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b33  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [33]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b34  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [34]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b35  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [35]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b36  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [36]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b37  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [37]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b38  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [38]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b39  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [39]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b4  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [4]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b40  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [40]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b41  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [41]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b42  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [42]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b43  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [43]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b44  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [44]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b45  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [45]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b46  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [46]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b47  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [47]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b48  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [48]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b49  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [49]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b5  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [5]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b50  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [50]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b51  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [51]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b52  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [52]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b53  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [53]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b54  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [54]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b55  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [55]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b56  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [56]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b57  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [57]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b58  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [58]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b59  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [59]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b6  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [6]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b60  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [60]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b61  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [61]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b62  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [62]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b63  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [63]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b7  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [7]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b8  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [8]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux12_b9  (
    .i0(1'b0),
    .i1(\cu_ru/sscratch [9]),
    .sel(\cu_ru/read_sscratch_sel ),
    .o(\cu_ru/n70 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  binary_mux_s1_w1 \cu_ru/mux13_b0  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [0]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b1  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [1]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b10  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [10]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b11  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [11]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b12  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [12]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b13  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [13]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b14  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [14]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b15  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [15]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b16  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [16]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b17  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [17]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b18  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [18]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b19  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [19]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b2  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [2]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b20  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [20]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b21  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [21]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b22  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [22]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b23  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [23]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b24  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [24]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b25  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [25]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b26  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [26]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b27  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [27]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b28  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [28]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b29  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [29]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b3  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [3]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b30  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [30]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b31  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [31]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b32  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [32]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b33  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [33]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b34  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [34]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b35  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [35]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b36  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [36]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b37  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [37]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b38  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [38]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b39  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [39]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b4  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [4]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b40  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [40]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b41  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [41]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b42  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [42]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b43  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [43]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b44  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [44]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b45  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [45]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b46  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [46]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b47  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [47]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b48  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [48]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b49  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [49]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b5  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [5]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b50  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [50]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b51  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [51]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b52  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [52]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b53  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [53]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b54  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [54]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b55  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [55]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b56  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [56]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b57  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [57]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b58  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [58]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b59  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [59]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b6  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [6]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b60  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [60]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b61  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [61]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b62  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [62]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b63  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [63]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b7  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [7]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b8  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [8]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux13_b9  (
    .i0(1'b0),
    .i1(\cu_ru/sepc [9]),
    .sel(\cu_ru/read_sepc_sel ),
    .o(\cu_ru/n72 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  binary_mux_s1_w1 \cu_ru/mux14_b0  (
    .i0(1'b0),
    .i1(\cu_ru/scause [0]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b1  (
    .i0(1'b0),
    .i1(\cu_ru/scause [1]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b10  (
    .i0(1'b0),
    .i1(\cu_ru/scause [10]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b11  (
    .i0(1'b0),
    .i1(\cu_ru/scause [11]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b12  (
    .i0(1'b0),
    .i1(\cu_ru/scause [12]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b13  (
    .i0(1'b0),
    .i1(\cu_ru/scause [13]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b14  (
    .i0(1'b0),
    .i1(\cu_ru/scause [14]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b15  (
    .i0(1'b0),
    .i1(\cu_ru/scause [15]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b16  (
    .i0(1'b0),
    .i1(\cu_ru/scause [16]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b17  (
    .i0(1'b0),
    .i1(\cu_ru/scause [17]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b18  (
    .i0(1'b0),
    .i1(\cu_ru/scause [18]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b19  (
    .i0(1'b0),
    .i1(\cu_ru/scause [19]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b2  (
    .i0(1'b0),
    .i1(\cu_ru/scause [2]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b20  (
    .i0(1'b0),
    .i1(\cu_ru/scause [20]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b21  (
    .i0(1'b0),
    .i1(\cu_ru/scause [21]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b22  (
    .i0(1'b0),
    .i1(\cu_ru/scause [22]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b23  (
    .i0(1'b0),
    .i1(\cu_ru/scause [23]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b24  (
    .i0(1'b0),
    .i1(\cu_ru/scause [24]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b25  (
    .i0(1'b0),
    .i1(\cu_ru/scause [25]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b26  (
    .i0(1'b0),
    .i1(\cu_ru/scause [26]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b27  (
    .i0(1'b0),
    .i1(\cu_ru/scause [27]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b28  (
    .i0(1'b0),
    .i1(\cu_ru/scause [28]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b29  (
    .i0(1'b0),
    .i1(\cu_ru/scause [29]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b3  (
    .i0(1'b0),
    .i1(\cu_ru/scause [3]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b30  (
    .i0(1'b0),
    .i1(\cu_ru/scause [30]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b31  (
    .i0(1'b0),
    .i1(\cu_ru/scause [31]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b32  (
    .i0(1'b0),
    .i1(\cu_ru/scause [32]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b33  (
    .i0(1'b0),
    .i1(\cu_ru/scause [33]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b34  (
    .i0(1'b0),
    .i1(\cu_ru/scause [34]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b35  (
    .i0(1'b0),
    .i1(\cu_ru/scause [35]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b36  (
    .i0(1'b0),
    .i1(\cu_ru/scause [36]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b37  (
    .i0(1'b0),
    .i1(\cu_ru/scause [37]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b38  (
    .i0(1'b0),
    .i1(\cu_ru/scause [38]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b39  (
    .i0(1'b0),
    .i1(\cu_ru/scause [39]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b4  (
    .i0(1'b0),
    .i1(\cu_ru/scause [4]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b40  (
    .i0(1'b0),
    .i1(\cu_ru/scause [40]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b41  (
    .i0(1'b0),
    .i1(\cu_ru/scause [41]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b42  (
    .i0(1'b0),
    .i1(\cu_ru/scause [42]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b43  (
    .i0(1'b0),
    .i1(\cu_ru/scause [43]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b44  (
    .i0(1'b0),
    .i1(\cu_ru/scause [44]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b45  (
    .i0(1'b0),
    .i1(\cu_ru/scause [45]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b46  (
    .i0(1'b0),
    .i1(\cu_ru/scause [46]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b47  (
    .i0(1'b0),
    .i1(\cu_ru/scause [47]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b48  (
    .i0(1'b0),
    .i1(\cu_ru/scause [48]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b49  (
    .i0(1'b0),
    .i1(\cu_ru/scause [49]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b5  (
    .i0(1'b0),
    .i1(\cu_ru/scause [5]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b50  (
    .i0(1'b0),
    .i1(\cu_ru/scause [50]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b51  (
    .i0(1'b0),
    .i1(\cu_ru/scause [51]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b52  (
    .i0(1'b0),
    .i1(\cu_ru/scause [52]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b53  (
    .i0(1'b0),
    .i1(\cu_ru/scause [53]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b54  (
    .i0(1'b0),
    .i1(\cu_ru/scause [54]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b55  (
    .i0(1'b0),
    .i1(\cu_ru/scause [55]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b56  (
    .i0(1'b0),
    .i1(\cu_ru/scause [56]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b57  (
    .i0(1'b0),
    .i1(\cu_ru/scause [57]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b58  (
    .i0(1'b0),
    .i1(\cu_ru/scause [58]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b59  (
    .i0(1'b0),
    .i1(\cu_ru/scause [59]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b6  (
    .i0(1'b0),
    .i1(\cu_ru/scause [6]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b60  (
    .i0(1'b0),
    .i1(\cu_ru/scause [60]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b61  (
    .i0(1'b0),
    .i1(\cu_ru/scause [61]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b62  (
    .i0(1'b0),
    .i1(\cu_ru/scause [62]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b63  (
    .i0(1'b0),
    .i1(\cu_ru/scause [63]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b7  (
    .i0(1'b0),
    .i1(\cu_ru/scause [7]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b8  (
    .i0(1'b0),
    .i1(\cu_ru/scause [8]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux14_b9  (
    .i0(1'b0),
    .i1(\cu_ru/scause [9]),
    .sel(\cu_ru/read_scause_sel ),
    .o(\cu_ru/n74 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  binary_mux_s1_w1 \cu_ru/mux15_b0  (
    .i0(1'b0),
    .i1(\cu_ru/stval [0]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b1  (
    .i0(1'b0),
    .i1(\cu_ru/stval [1]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b10  (
    .i0(1'b0),
    .i1(\cu_ru/stval [10]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b11  (
    .i0(1'b0),
    .i1(\cu_ru/stval [11]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b12  (
    .i0(1'b0),
    .i1(\cu_ru/stval [12]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b13  (
    .i0(1'b0),
    .i1(\cu_ru/stval [13]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b14  (
    .i0(1'b0),
    .i1(\cu_ru/stval [14]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b15  (
    .i0(1'b0),
    .i1(\cu_ru/stval [15]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b16  (
    .i0(1'b0),
    .i1(\cu_ru/stval [16]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b17  (
    .i0(1'b0),
    .i1(\cu_ru/stval [17]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b18  (
    .i0(1'b0),
    .i1(\cu_ru/stval [18]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b19  (
    .i0(1'b0),
    .i1(\cu_ru/stval [19]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b2  (
    .i0(1'b0),
    .i1(\cu_ru/stval [2]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b20  (
    .i0(1'b0),
    .i1(\cu_ru/stval [20]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b21  (
    .i0(1'b0),
    .i1(\cu_ru/stval [21]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b22  (
    .i0(1'b0),
    .i1(\cu_ru/stval [22]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b23  (
    .i0(1'b0),
    .i1(\cu_ru/stval [23]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b24  (
    .i0(1'b0),
    .i1(\cu_ru/stval [24]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b25  (
    .i0(1'b0),
    .i1(\cu_ru/stval [25]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b26  (
    .i0(1'b0),
    .i1(\cu_ru/stval [26]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b27  (
    .i0(1'b0),
    .i1(\cu_ru/stval [27]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b28  (
    .i0(1'b0),
    .i1(\cu_ru/stval [28]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b29  (
    .i0(1'b0),
    .i1(\cu_ru/stval [29]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b3  (
    .i0(1'b0),
    .i1(\cu_ru/stval [3]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b30  (
    .i0(1'b0),
    .i1(\cu_ru/stval [30]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b31  (
    .i0(1'b0),
    .i1(\cu_ru/stval [31]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b32  (
    .i0(1'b0),
    .i1(\cu_ru/stval [32]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b33  (
    .i0(1'b0),
    .i1(\cu_ru/stval [33]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b34  (
    .i0(1'b0),
    .i1(\cu_ru/stval [34]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b35  (
    .i0(1'b0),
    .i1(\cu_ru/stval [35]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b36  (
    .i0(1'b0),
    .i1(\cu_ru/stval [36]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b37  (
    .i0(1'b0),
    .i1(\cu_ru/stval [37]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b38  (
    .i0(1'b0),
    .i1(\cu_ru/stval [38]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b39  (
    .i0(1'b0),
    .i1(\cu_ru/stval [39]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b4  (
    .i0(1'b0),
    .i1(\cu_ru/stval [4]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b40  (
    .i0(1'b0),
    .i1(\cu_ru/stval [40]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b41  (
    .i0(1'b0),
    .i1(\cu_ru/stval [41]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b42  (
    .i0(1'b0),
    .i1(\cu_ru/stval [42]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b43  (
    .i0(1'b0),
    .i1(\cu_ru/stval [43]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b44  (
    .i0(1'b0),
    .i1(\cu_ru/stval [44]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b45  (
    .i0(1'b0),
    .i1(\cu_ru/stval [45]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b46  (
    .i0(1'b0),
    .i1(\cu_ru/stval [46]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b47  (
    .i0(1'b0),
    .i1(\cu_ru/stval [47]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b48  (
    .i0(1'b0),
    .i1(\cu_ru/stval [48]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b49  (
    .i0(1'b0),
    .i1(\cu_ru/stval [49]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b5  (
    .i0(1'b0),
    .i1(\cu_ru/stval [5]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b50  (
    .i0(1'b0),
    .i1(\cu_ru/stval [50]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b51  (
    .i0(1'b0),
    .i1(\cu_ru/stval [51]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b52  (
    .i0(1'b0),
    .i1(\cu_ru/stval [52]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b53  (
    .i0(1'b0),
    .i1(\cu_ru/stval [53]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b54  (
    .i0(1'b0),
    .i1(\cu_ru/stval [54]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b55  (
    .i0(1'b0),
    .i1(\cu_ru/stval [55]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b56  (
    .i0(1'b0),
    .i1(\cu_ru/stval [56]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b57  (
    .i0(1'b0),
    .i1(\cu_ru/stval [57]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b58  (
    .i0(1'b0),
    .i1(\cu_ru/stval [58]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b59  (
    .i0(1'b0),
    .i1(\cu_ru/stval [59]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b6  (
    .i0(1'b0),
    .i1(\cu_ru/stval [6]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b60  (
    .i0(1'b0),
    .i1(\cu_ru/stval [60]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b61  (
    .i0(1'b0),
    .i1(\cu_ru/stval [61]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b62  (
    .i0(1'b0),
    .i1(\cu_ru/stval [62]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b63  (
    .i0(1'b0),
    .i1(\cu_ru/stval [63]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b7  (
    .i0(1'b0),
    .i1(\cu_ru/stval [7]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b8  (
    .i0(1'b0),
    .i1(\cu_ru/stval [8]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux15_b9  (
    .i0(1'b0),
    .i1(\cu_ru/stval [9]),
    .sel(\cu_ru/read_stval_sel ),
    .o(\cu_ru/n76 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  binary_mux_s1_w1 \cu_ru/mux16_b1  (
    .i0(1'b0),
    .i1(\cu_ru/m_sip [1]),
    .sel(\cu_ru/read_sip_sel ),
    .o(\cu_ru/n78 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(684)
  binary_mux_s1_w1 \cu_ru/mux16_b5  (
    .i0(1'b0),
    .i1(\cu_ru/m_sip [5]),
    .sel(\cu_ru/read_sip_sel ),
    .o(\cu_ru/n78 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(684)
  binary_mux_s1_w1 \cu_ru/mux16_b9  (
    .i0(1'b0),
    .i1(\cu_ru/m_sip [9]),
    .sel(\cu_ru/read_sip_sel ),
    .o(\cu_ru/n78 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(684)
  binary_mux_s1_w1 \cu_ru/mux17_b0  (
    .i0(1'b0),
    .i1(satp[0]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b1  (
    .i0(1'b0),
    .i1(satp[1]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b10  (
    .i0(1'b0),
    .i1(satp[10]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b11  (
    .i0(1'b0),
    .i1(satp[11]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b12  (
    .i0(1'b0),
    .i1(satp[12]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b13  (
    .i0(1'b0),
    .i1(satp[13]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b14  (
    .i0(1'b0),
    .i1(satp[14]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b15  (
    .i0(1'b0),
    .i1(satp[15]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b16  (
    .i0(1'b0),
    .i1(satp[16]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b17  (
    .i0(1'b0),
    .i1(satp[17]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b18  (
    .i0(1'b0),
    .i1(satp[18]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b19  (
    .i0(1'b0),
    .i1(satp[19]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b2  (
    .i0(1'b0),
    .i1(satp[2]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b20  (
    .i0(1'b0),
    .i1(satp[20]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b21  (
    .i0(1'b0),
    .i1(satp[21]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b22  (
    .i0(1'b0),
    .i1(satp[22]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b23  (
    .i0(1'b0),
    .i1(satp[23]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b24  (
    .i0(1'b0),
    .i1(satp[24]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b25  (
    .i0(1'b0),
    .i1(satp[25]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b26  (
    .i0(1'b0),
    .i1(satp[26]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b27  (
    .i0(1'b0),
    .i1(satp[27]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b28  (
    .i0(1'b0),
    .i1(satp[28]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b29  (
    .i0(1'b0),
    .i1(satp[29]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b3  (
    .i0(1'b0),
    .i1(satp[3]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b30  (
    .i0(1'b0),
    .i1(satp[30]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b31  (
    .i0(1'b0),
    .i1(satp[31]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b32  (
    .i0(1'b0),
    .i1(satp[32]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b33  (
    .i0(1'b0),
    .i1(satp[33]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b34  (
    .i0(1'b0),
    .i1(satp[34]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b35  (
    .i0(1'b0),
    .i1(satp[35]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b36  (
    .i0(1'b0),
    .i1(satp[36]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b37  (
    .i0(1'b0),
    .i1(satp[37]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b38  (
    .i0(1'b0),
    .i1(satp[38]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b39  (
    .i0(1'b0),
    .i1(satp[39]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b4  (
    .i0(1'b0),
    .i1(satp[4]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b40  (
    .i0(1'b0),
    .i1(satp[40]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b41  (
    .i0(1'b0),
    .i1(satp[41]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b42  (
    .i0(1'b0),
    .i1(satp[42]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b43  (
    .i0(1'b0),
    .i1(satp[43]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b5  (
    .i0(1'b0),
    .i1(satp[5]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b6  (
    .i0(1'b0),
    .i1(satp[6]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b60  (
    .i0(1'b0),
    .i1(satp[60]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b61  (
    .i0(1'b0),
    .i1(satp[61]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b62  (
    .i0(1'b0),
    .i1(satp[62]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b63  (
    .i0(1'b0),
    .i1(satp[63]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b7  (
    .i0(1'b0),
    .i1(satp[7]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b8  (
    .i0(1'b0),
    .i1(satp[8]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux17_b9  (
    .i0(1'b0),
    .i1(satp[9]),
    .sel(\cu_ru/read_satp_sel ),
    .o(\cu_ru/n80 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  binary_mux_s1_w1 \cu_ru/mux18_b14  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\cu_ru/read_mvendorid_sel ),
    .o(\cu_ru/n82 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  binary_mux_s1_w1 \cu_ru/mux19_b10  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\cu_ru/read_marchid_sel ),
    .o(\cu_ru/n84 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  binary_mux_s1_w1 \cu_ru/mux20_b2  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\cu_ru/read_mimp_sel ),
    .o(\cu_ru/n86 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(688)
  binary_mux_s1_w1 \cu_ru/mux22_b1  (
    .i0(1'b0),
    .i1(\cu_ru/mstatus [1]),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b11  (
    .i0(1'b0),
    .i1(\cu_ru/mstatus [11]),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b12  (
    .i0(1'b0),
    .i1(\cu_ru/mstatus [12]),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b17  (
    .i0(1'b0),
    .i1(mprv),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b18  (
    .i0(1'b0),
    .i1(sum),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b19  (
    .i0(1'b0),
    .i1(mxr),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b20  (
    .i0(1'b0),
    .i1(tvm),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b21  (
    .i0(1'b0),
    .i1(tw),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b22  (
    .i0(1'b0),
    .i1(tsr),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b3  (
    .i0(1'b0),
    .i1(\cu_ru/mie ),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b32  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b5  (
    .i0(1'b0),
    .i1(\cu_ru/mstatus [5]),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b7  (
    .i0(1'b0),
    .i1(\cu_ru/mstatus [7]),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux22_b8  (
    .i0(1'b0),
    .i1(\cu_ru/mstatus [8]),
    .sel(\cu_ru/read_mstatus_sel ),
    .o(\cu_ru/n90 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  binary_mux_s1_w1 \cu_ru/mux24_b0  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [0]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b1  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [1]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b12  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [12]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b13  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [13]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b15  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [15]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b2  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [2]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b3  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [3]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b4  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [4]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b5  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [5]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b6  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [6]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b7  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [7]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b8  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [8]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux24_b9  (
    .i0(1'b0),
    .i1(\cu_ru/medeleg [9]),
    .sel(\cu_ru/read_medeleg_sel ),
    .o(\cu_ru/n94 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  binary_mux_s1_w1 \cu_ru/mux25_b1  (
    .i0(1'b0),
    .i1(\cu_ru/mideleg [1]),
    .sel(\cu_ru/read_mideleg_sel ),
    .o(\cu_ru/n96 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(693)
  binary_mux_s1_w1 \cu_ru/mux25_b5  (
    .i0(1'b0),
    .i1(\cu_ru/mideleg [5]),
    .sel(\cu_ru/read_mideleg_sel ),
    .o(\cu_ru/n96 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(693)
  binary_mux_s1_w1 \cu_ru/mux25_b9  (
    .i0(1'b0),
    .i1(\cu_ru/mideleg [9]),
    .sel(\cu_ru/read_mideleg_sel ),
    .o(\cu_ru/n96 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(693)
  binary_mux_s1_w1 \cu_ru/mux26_b0  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [0]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b1  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [1]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b10  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [10]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b11  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [11]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b12  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [12]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b13  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [13]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b14  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [14]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b15  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [15]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b16  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [16]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b17  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [17]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b18  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [18]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b19  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [19]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b2  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [2]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b20  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [20]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b21  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [21]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b22  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [22]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b23  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [23]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b24  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [24]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b25  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [25]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b26  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [26]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b27  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [27]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b28  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [28]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b29  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [29]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b3  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [3]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b30  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [30]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b31  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [31]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b32  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [32]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b33  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [33]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b34  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [34]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b35  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [35]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b36  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [36]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b37  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [37]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b38  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [38]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b39  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [39]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b4  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [4]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b40  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [40]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b41  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [41]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b42  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [42]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b43  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [43]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b44  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [44]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b45  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [45]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b46  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [46]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b47  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [47]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b48  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [48]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b49  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [49]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b5  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [5]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b50  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [50]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b51  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [51]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b52  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [52]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b53  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [53]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b54  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [54]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b55  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [55]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b56  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [56]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b57  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [57]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b58  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [58]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b59  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [59]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b6  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [6]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b60  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [60]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b61  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [61]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b62  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [62]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b63  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [63]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b7  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [7]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b8  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [8]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux26_b9  (
    .i0(1'b0),
    .i1(\cu_ru/mtvec [9]),
    .sel(\cu_ru/read_mtvec_sel ),
    .o(\cu_ru/n100 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  binary_mux_s1_w1 \cu_ru/mux27_b0  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [0]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b1  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [1]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b10  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [10]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b11  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [11]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b12  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [12]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b13  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [13]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b14  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [14]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b15  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [15]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b16  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [16]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b17  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [17]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b18  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [18]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b19  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [19]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b2  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [2]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b20  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [20]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b21  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [21]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b22  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [22]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b23  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [23]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b24  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [24]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b25  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [25]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b26  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [26]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b27  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [27]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b28  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [28]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b29  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [29]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b3  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [3]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b30  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [30]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b31  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [31]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b32  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [32]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b33  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [33]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b34  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [34]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b35  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [35]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b36  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [36]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b37  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [37]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b38  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [38]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b39  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [39]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b4  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [4]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b40  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [40]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b41  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [41]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b42  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [42]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b43  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [43]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b44  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [44]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b45  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [45]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b46  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [46]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b47  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [47]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b48  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [48]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b49  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [49]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b5  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [5]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b50  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [50]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b51  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [51]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b52  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [52]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b53  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [53]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b54  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [54]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b55  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [55]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b56  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [56]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b57  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [57]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b58  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [58]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b59  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [59]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b6  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [6]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b60  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [60]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b61  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [61]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b62  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [62]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b63  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [63]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b7  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [7]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b8  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [8]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux27_b9  (
    .i0(1'b0),
    .i1(\cu_ru/mscratch [9]),
    .sel(\cu_ru/read_mscratch_sel ),
    .o(\cu_ru/n102 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  binary_mux_s1_w1 \cu_ru/mux28_b0  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [0]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b1  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [1]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b10  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [10]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b11  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [11]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b12  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [12]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b13  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [13]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b14  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [14]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b15  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [15]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b16  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [16]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b17  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [17]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b18  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [18]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b19  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [19]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b2  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [2]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b20  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [20]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b21  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [21]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b22  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [22]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b23  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [23]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b24  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [24]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b25  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [25]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b26  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [26]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b27  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [27]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b28  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [28]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b29  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [29]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b3  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [3]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b30  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [30]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b31  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [31]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b32  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [32]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b33  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [33]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b34  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [34]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b35  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [35]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b36  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [36]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b37  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [37]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b38  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [38]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b39  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [39]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b4  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [4]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b40  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [40]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b41  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [41]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b42  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [42]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b43  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [43]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b44  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [44]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b45  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [45]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b46  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [46]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b47  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [47]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b48  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [48]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b49  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [49]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b5  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [5]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b50  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [50]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b51  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [51]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b52  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [52]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b53  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [53]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b54  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [54]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b55  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [55]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b56  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [56]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b57  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [57]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b58  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [58]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b59  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [59]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b6  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [6]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b60  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [60]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b61  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [61]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b62  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [62]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b63  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [63]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b7  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [7]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b8  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [8]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux28_b9  (
    .i0(1'b0),
    .i1(\cu_ru/mepc [9]),
    .sel(\cu_ru/read_mepc_sel ),
    .o(\cu_ru/n104 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  binary_mux_s1_w1 \cu_ru/mux29_b0  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [0]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b1  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [1]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b10  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [10]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b11  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [11]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b12  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [12]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b13  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [13]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b14  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [14]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b15  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [15]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b16  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [16]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b17  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [17]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b18  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [18]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b19  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [19]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b2  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [2]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b20  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [20]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b21  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [21]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b22  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [22]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b23  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [23]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b24  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [24]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b25  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [25]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b26  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [26]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b27  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [27]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b28  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [28]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b29  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [29]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b3  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [3]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b30  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [30]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b31  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [31]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b32  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [32]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b33  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [33]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b34  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [34]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b35  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [35]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b36  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [36]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b37  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [37]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b38  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [38]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b39  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [39]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b4  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [4]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b40  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [40]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b41  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [41]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b42  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [42]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b43  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [43]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b44  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [44]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b45  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [45]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b46  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [46]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b47  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [47]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b48  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [48]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b49  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [49]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b5  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [5]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b50  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [50]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b51  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [51]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b52  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [52]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b53  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [53]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b54  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [54]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b55  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [55]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b56  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [56]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b57  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [57]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b58  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [58]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b59  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [59]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b6  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [6]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b60  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [60]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b61  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [61]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b62  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [62]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b63  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [63]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b7  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [7]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b8  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [8]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux29_b9  (
    .i0(1'b0),
    .i1(\cu_ru/mcause [9]),
    .sel(\cu_ru/read_mcause_sel ),
    .o(\cu_ru/n106 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  binary_mux_s1_w1 \cu_ru/mux2_b0  (
    .i0(\cu_ru/n47 [0]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b1  (
    .i0(\cu_ru/n47 [1]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b10  (
    .i0(\cu_ru/n47 [10]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b11  (
    .i0(\cu_ru/n47 [11]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b12  (
    .i0(\cu_ru/n47 [12]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b13  (
    .i0(\cu_ru/n47 [13]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b14  (
    .i0(\cu_ru/n47 [14]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b15  (
    .i0(\cu_ru/n47 [15]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b16  (
    .i0(\cu_ru/n47 [16]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b17  (
    .i0(\cu_ru/n47 [17]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b18  (
    .i0(\cu_ru/n47 [18]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b19  (
    .i0(\cu_ru/n47 [19]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b2  (
    .i0(\cu_ru/n47 [2]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b20  (
    .i0(\cu_ru/n47 [20]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b21  (
    .i0(\cu_ru/n47 [21]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b22  (
    .i0(\cu_ru/n47 [22]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b23  (
    .i0(\cu_ru/n47 [23]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b24  (
    .i0(\cu_ru/n47 [24]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b25  (
    .i0(\cu_ru/n47 [25]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b26  (
    .i0(\cu_ru/n47 [26]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b27  (
    .i0(\cu_ru/n47 [27]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b28  (
    .i0(\cu_ru/n47 [28]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b29  (
    .i0(\cu_ru/n47 [29]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b3  (
    .i0(\cu_ru/n47 [3]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b30  (
    .i0(\cu_ru/n47 [30]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b31  (
    .i0(\cu_ru/n47 [31]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b32  (
    .i0(\cu_ru/n47 [32]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b33  (
    .i0(\cu_ru/n47 [33]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b34  (
    .i0(\cu_ru/n47 [34]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b35  (
    .i0(\cu_ru/n47 [35]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b36  (
    .i0(\cu_ru/n47 [36]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b37  (
    .i0(\cu_ru/n47 [37]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b38  (
    .i0(\cu_ru/n47 [38]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b39  (
    .i0(\cu_ru/n47 [39]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b4  (
    .i0(\cu_ru/n47 [4]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b40  (
    .i0(\cu_ru/n47 [40]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b41  (
    .i0(\cu_ru/n47 [41]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b42  (
    .i0(\cu_ru/n47 [42]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b43  (
    .i0(\cu_ru/n47 [43]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b44  (
    .i0(\cu_ru/n47 [44]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b45  (
    .i0(\cu_ru/n47 [45]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b46  (
    .i0(\cu_ru/n47 [46]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b47  (
    .i0(\cu_ru/n47 [47]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b48  (
    .i0(\cu_ru/n47 [48]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b49  (
    .i0(\cu_ru/n47 [49]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b5  (
    .i0(\cu_ru/n47 [5]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b50  (
    .i0(\cu_ru/n47 [50]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b51  (
    .i0(\cu_ru/n47 [51]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b52  (
    .i0(\cu_ru/n47 [52]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b53  (
    .i0(\cu_ru/n47 [53]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b54  (
    .i0(\cu_ru/n47 [54]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b55  (
    .i0(\cu_ru/n47 [55]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b56  (
    .i0(\cu_ru/n47 [56]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b57  (
    .i0(\cu_ru/n47 [57]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b58  (
    .i0(\cu_ru/n47 [58]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b59  (
    .i0(\cu_ru/n47 [59]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b6  (
    .i0(\cu_ru/n47 [6]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b60  (
    .i0(\cu_ru/n47 [60]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b61  (
    .i0(\cu_ru/n47 [61]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b62  (
    .i0(\cu_ru/n47 [62]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b63  (
    .i0(\cu_ru/n47 [63]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b7  (
    .i0(\cu_ru/n47 [7]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b8  (
    .i0(\cu_ru/n47 [8]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux2_b9  (
    .i0(\cu_ru/n47 [9]),
    .i1(1'b0),
    .sel(\cu_ru/n45 ),
    .o(rs1_data[9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  binary_mux_s1_w1 \cu_ru/mux30_b0  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [0]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b1  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [1]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b10  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [10]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b11  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [11]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b12  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [12]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b13  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [13]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b14  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [14]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b15  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [15]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b16  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [16]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b17  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [17]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b18  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [18]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b19  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [19]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b2  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [2]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b20  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [20]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b21  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [21]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b22  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [22]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b23  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [23]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b24  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [24]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b25  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [25]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b26  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [26]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b27  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [27]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b28  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [28]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b29  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [29]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b3  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [3]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b30  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [30]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b31  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [31]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b32  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [32]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b33  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [33]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b34  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [34]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b35  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [35]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b36  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [36]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b37  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [37]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b38  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [38]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b39  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [39]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b4  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [4]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b40  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [40]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b41  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [41]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b42  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [42]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b43  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [43]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b44  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [44]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b45  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [45]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b46  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [46]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b47  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [47]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b48  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [48]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b49  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [49]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b5  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [5]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b50  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [50]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b51  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [51]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b52  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [52]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b53  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [53]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b54  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [54]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b55  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [55]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b56  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [56]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b57  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [57]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b58  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [58]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b59  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [59]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b6  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [6]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b60  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [60]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b61  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [61]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b62  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [62]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b63  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [63]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b7  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [7]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b8  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [8]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux30_b9  (
    .i0(1'b0),
    .i1(\cu_ru/mtval [9]),
    .sel(\cu_ru/read_mtval_sel ),
    .o(\cu_ru/n108 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  binary_mux_s1_w1 \cu_ru/mux31_b1  (
    .i0(1'b0),
    .i1(\cu_ru/m_sip [1]),
    .sel(\cu_ru/read_mip_sel ),
    .o(\cu_ru/n110 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  binary_mux_s1_w1 \cu_ru/mux31_b11  (
    .i0(1'b0),
    .i1(\cu_ru/m_sip [11]),
    .sel(\cu_ru/read_mip_sel ),
    .o(\cu_ru/n110 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  binary_mux_s1_w1 \cu_ru/mux31_b3  (
    .i0(1'b0),
    .i1(\cu_ru/m_sip [3]),
    .sel(\cu_ru/read_mip_sel ),
    .o(\cu_ru/n110 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  binary_mux_s1_w1 \cu_ru/mux31_b5  (
    .i0(1'b0),
    .i1(\cu_ru/m_sip [5]),
    .sel(\cu_ru/read_mip_sel ),
    .o(\cu_ru/n110 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  binary_mux_s1_w1 \cu_ru/mux31_b7  (
    .i0(1'b0),
    .i1(\cu_ru/m_sip [7]),
    .sel(\cu_ru/read_mip_sel ),
    .o(\cu_ru/n110 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  binary_mux_s1_w1 \cu_ru/mux31_b9  (
    .i0(1'b0),
    .i1(\cu_ru/m_sip [9]),
    .sel(\cu_ru/read_mip_sel ),
    .o(\cu_ru/n110 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  binary_mux_s1_w1 \cu_ru/mux32_b0  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [0]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b1  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [1]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b10  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [10]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b11  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [11]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b12  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [12]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b13  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [13]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b14  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [14]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b15  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [15]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b16  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [16]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b17  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [17]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b18  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [18]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b19  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [19]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b2  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [2]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b20  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [20]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b21  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [21]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b22  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [22]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b23  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [23]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b24  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [24]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b25  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [25]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b26  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [26]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b27  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [27]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b28  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [28]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b29  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [29]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b3  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [3]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b30  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [30]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b31  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [31]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b32  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [32]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b33  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [33]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b34  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [34]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b35  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [35]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b36  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [36]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b37  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [37]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b38  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [38]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b39  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [39]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b4  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [4]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b40  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [40]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b41  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [41]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b42  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [42]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b43  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [43]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b44  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [44]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b45  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [45]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b46  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [46]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b47  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [47]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b48  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [48]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b49  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [49]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b5  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [5]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b50  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [50]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b51  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [51]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b52  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [52]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b53  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [53]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b54  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [54]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b55  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [55]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b56  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [56]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b57  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [57]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b58  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [58]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b59  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [59]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b6  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [6]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b60  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [60]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b61  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [61]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b62  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [62]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b63  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [63]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b7  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [7]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b8  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [8]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux32_b9  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [9]),
    .sel(\cu_ru/read_mcycle_sel ),
    .o(\cu_ru/n112 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  binary_mux_s1_w1 \cu_ru/mux33_b0  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [0]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b1  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [1]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b10  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [10]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b11  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [11]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b12  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [12]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b13  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [13]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b14  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [14]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b15  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [15]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b16  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [16]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b17  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [17]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b18  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [18]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b19  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [19]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b2  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [2]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b20  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [20]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b21  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [21]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b22  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [22]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b23  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [23]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b24  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [24]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b25  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [25]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b26  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [26]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b27  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [27]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b28  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [28]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b29  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [29]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b3  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [3]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b30  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [30]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b31  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [31]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b32  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [32]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b33  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [33]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b34  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [34]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b35  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [35]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b36  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [36]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b37  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [37]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b38  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [38]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b39  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [39]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b4  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [4]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b40  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [40]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b41  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [41]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b42  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [42]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b43  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [43]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b44  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [44]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b45  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [45]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b46  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [46]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b47  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [47]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b48  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [48]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b49  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [49]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b5  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [5]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b50  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [50]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b51  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [51]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b52  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [52]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b53  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [53]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b54  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [54]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b55  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [55]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b56  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [56]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b57  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [57]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b58  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [58]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b59  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [59]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b6  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [6]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b60  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [60]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b61  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [61]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b62  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [62]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b63  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [63]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b7  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [7]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b8  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [8]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  binary_mux_s1_w1 \cu_ru/mux33_b9  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [9]),
    .sel(\cu_ru/read_minstret_sel ),
    .o(\cu_ru/n114 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  AL_MUX \cu_ru/mux34_b0  (
    .i0(\cu_ru/tvec [4]),
    .i1(\cu_ru/n43 [0]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [2]));
  and \cu_ru/mux34_b0_sel_is_2  (\cu_ru/mux34_b0_sel_is_2_o , \cu_ru/exception_neg , \cu_ru/tvec [0]);
  AL_MUX \cu_ru/mux34_b1  (
    .i0(\cu_ru/tvec [5]),
    .i1(\cu_ru/n43 [1]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [3]));
  AL_MUX \cu_ru/mux34_b10  (
    .i0(\cu_ru/tvec [14]),
    .i1(\cu_ru/n43 [10]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [12]));
  AL_MUX \cu_ru/mux34_b11  (
    .i0(\cu_ru/tvec [15]),
    .i1(\cu_ru/n43 [11]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [13]));
  AL_MUX \cu_ru/mux34_b12  (
    .i0(\cu_ru/tvec [16]),
    .i1(\cu_ru/n43 [12]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [14]));
  AL_MUX \cu_ru/mux34_b13  (
    .i0(\cu_ru/tvec [17]),
    .i1(\cu_ru/n43 [13]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [15]));
  AL_MUX \cu_ru/mux34_b14  (
    .i0(\cu_ru/tvec [18]),
    .i1(\cu_ru/n43 [14]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [16]));
  AL_MUX \cu_ru/mux34_b15  (
    .i0(\cu_ru/tvec [19]),
    .i1(\cu_ru/n43 [15]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [17]));
  AL_MUX \cu_ru/mux34_b16  (
    .i0(\cu_ru/tvec [20]),
    .i1(\cu_ru/n43 [16]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [18]));
  AL_MUX \cu_ru/mux34_b17  (
    .i0(\cu_ru/tvec [21]),
    .i1(\cu_ru/n43 [17]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [19]));
  AL_MUX \cu_ru/mux34_b18  (
    .i0(\cu_ru/tvec [22]),
    .i1(\cu_ru/n43 [18]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [20]));
  AL_MUX \cu_ru/mux34_b19  (
    .i0(\cu_ru/tvec [23]),
    .i1(\cu_ru/n43 [19]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [21]));
  AL_MUX \cu_ru/mux34_b2  (
    .i0(\cu_ru/tvec [6]),
    .i1(\cu_ru/n43 [2]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [4]));
  AL_MUX \cu_ru/mux34_b20  (
    .i0(\cu_ru/tvec [24]),
    .i1(\cu_ru/n43 [20]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [22]));
  AL_MUX \cu_ru/mux34_b21  (
    .i0(\cu_ru/tvec [25]),
    .i1(\cu_ru/n43 [21]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [23]));
  AL_MUX \cu_ru/mux34_b22  (
    .i0(\cu_ru/tvec [26]),
    .i1(\cu_ru/n43 [22]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [24]));
  AL_MUX \cu_ru/mux34_b23  (
    .i0(\cu_ru/tvec [27]),
    .i1(\cu_ru/n43 [23]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [25]));
  AL_MUX \cu_ru/mux34_b24  (
    .i0(\cu_ru/tvec [28]),
    .i1(\cu_ru/n43 [24]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [26]));
  AL_MUX \cu_ru/mux34_b25  (
    .i0(\cu_ru/tvec [29]),
    .i1(\cu_ru/n43 [25]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [27]));
  AL_MUX \cu_ru/mux34_b26  (
    .i0(\cu_ru/tvec [30]),
    .i1(\cu_ru/n43 [26]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [28]));
  AL_MUX \cu_ru/mux34_b27  (
    .i0(\cu_ru/tvec [31]),
    .i1(\cu_ru/n43 [27]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [29]));
  AL_MUX \cu_ru/mux34_b28  (
    .i0(\cu_ru/tvec [32]),
    .i1(\cu_ru/n43 [28]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [30]));
  AL_MUX \cu_ru/mux34_b29  (
    .i0(\cu_ru/tvec [33]),
    .i1(\cu_ru/n43 [29]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [31]));
  AL_MUX \cu_ru/mux34_b3  (
    .i0(\cu_ru/tvec [7]),
    .i1(\cu_ru/n43 [3]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [5]));
  AL_MUX \cu_ru/mux34_b30  (
    .i0(\cu_ru/tvec [34]),
    .i1(\cu_ru/n43 [30]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [32]));
  AL_MUX \cu_ru/mux34_b31  (
    .i0(\cu_ru/tvec [35]),
    .i1(\cu_ru/n43 [31]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [33]));
  AL_MUX \cu_ru/mux34_b32  (
    .i0(\cu_ru/tvec [36]),
    .i1(\cu_ru/n43 [32]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [34]));
  AL_MUX \cu_ru/mux34_b33  (
    .i0(\cu_ru/tvec [37]),
    .i1(\cu_ru/n43 [33]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [35]));
  AL_MUX \cu_ru/mux34_b34  (
    .i0(\cu_ru/tvec [38]),
    .i1(\cu_ru/n43 [34]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [36]));
  AL_MUX \cu_ru/mux34_b35  (
    .i0(\cu_ru/tvec [39]),
    .i1(\cu_ru/n43 [35]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [37]));
  AL_MUX \cu_ru/mux34_b36  (
    .i0(\cu_ru/tvec [40]),
    .i1(\cu_ru/n43 [36]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [38]));
  AL_MUX \cu_ru/mux34_b37  (
    .i0(\cu_ru/tvec [41]),
    .i1(\cu_ru/n43 [37]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [39]));
  AL_MUX \cu_ru/mux34_b38  (
    .i0(\cu_ru/tvec [42]),
    .i1(\cu_ru/n43 [38]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [40]));
  AL_MUX \cu_ru/mux34_b39  (
    .i0(\cu_ru/tvec [43]),
    .i1(\cu_ru/n43 [39]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [41]));
  AL_MUX \cu_ru/mux34_b4  (
    .i0(\cu_ru/tvec [8]),
    .i1(\cu_ru/n43 [4]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [6]));
  AL_MUX \cu_ru/mux34_b40  (
    .i0(\cu_ru/tvec [44]),
    .i1(\cu_ru/n43 [40]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [42]));
  AL_MUX \cu_ru/mux34_b41  (
    .i0(\cu_ru/tvec [45]),
    .i1(\cu_ru/n43 [41]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [43]));
  AL_MUX \cu_ru/mux34_b42  (
    .i0(\cu_ru/tvec [46]),
    .i1(\cu_ru/n43 [42]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [44]));
  AL_MUX \cu_ru/mux34_b43  (
    .i0(\cu_ru/tvec [47]),
    .i1(\cu_ru/n43 [43]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [45]));
  AL_MUX \cu_ru/mux34_b44  (
    .i0(\cu_ru/tvec [48]),
    .i1(\cu_ru/n43 [44]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [46]));
  AL_MUX \cu_ru/mux34_b45  (
    .i0(\cu_ru/tvec [49]),
    .i1(\cu_ru/n43 [45]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [47]));
  AL_MUX \cu_ru/mux34_b46  (
    .i0(\cu_ru/tvec [50]),
    .i1(\cu_ru/n43 [46]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [48]));
  AL_MUX \cu_ru/mux34_b47  (
    .i0(\cu_ru/tvec [51]),
    .i1(\cu_ru/n43 [47]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [49]));
  AL_MUX \cu_ru/mux34_b48  (
    .i0(\cu_ru/tvec [52]),
    .i1(\cu_ru/n43 [48]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [50]));
  AL_MUX \cu_ru/mux34_b49  (
    .i0(\cu_ru/tvec [53]),
    .i1(\cu_ru/n43 [49]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [51]));
  AL_MUX \cu_ru/mux34_b5  (
    .i0(\cu_ru/tvec [9]),
    .i1(\cu_ru/n43 [5]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [7]));
  AL_MUX \cu_ru/mux34_b50  (
    .i0(\cu_ru/tvec [54]),
    .i1(\cu_ru/n43 [50]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [52]));
  AL_MUX \cu_ru/mux34_b51  (
    .i0(\cu_ru/tvec [55]),
    .i1(\cu_ru/n43 [51]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [53]));
  AL_MUX \cu_ru/mux34_b52  (
    .i0(\cu_ru/tvec [56]),
    .i1(\cu_ru/n43 [52]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [54]));
  AL_MUX \cu_ru/mux34_b53  (
    .i0(\cu_ru/tvec [57]),
    .i1(\cu_ru/n43 [53]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [55]));
  AL_MUX \cu_ru/mux34_b54  (
    .i0(\cu_ru/tvec [58]),
    .i1(\cu_ru/n43 [54]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [56]));
  AL_MUX \cu_ru/mux34_b55  (
    .i0(\cu_ru/tvec [59]),
    .i1(\cu_ru/n43 [55]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [57]));
  AL_MUX \cu_ru/mux34_b56  (
    .i0(\cu_ru/tvec [60]),
    .i1(\cu_ru/n43 [56]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [58]));
  AL_MUX \cu_ru/mux34_b57  (
    .i0(\cu_ru/tvec [61]),
    .i1(\cu_ru/n43 [57]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [59]));
  AL_MUX \cu_ru/mux34_b58  (
    .i0(\cu_ru/tvec [62]),
    .i1(\cu_ru/n43 [58]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [60]));
  AL_MUX \cu_ru/mux34_b59  (
    .i0(\cu_ru/tvec [63]),
    .i1(\cu_ru/n43 [59]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [61]));
  AL_MUX \cu_ru/mux34_b6  (
    .i0(\cu_ru/tvec [10]),
    .i1(\cu_ru/n43 [6]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [8]));
  AL_MUX \cu_ru/mux34_b60  (
    .i0(1'b0),
    .i1(\cu_ru/add0_2_co ),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [62]));
  AL_MUX \cu_ru/mux34_b7  (
    .i0(\cu_ru/tvec [11]),
    .i1(\cu_ru/n43 [7]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [9]));
  AL_MUX \cu_ru/mux34_b8  (
    .i0(\cu_ru/tvec [12]),
    .i1(\cu_ru/n43 [8]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [10]));
  AL_MUX \cu_ru/mux34_b9  (
    .i0(\cu_ru/tvec [13]),
    .i1(\cu_ru/n43 [9]),
    .sel(\cu_ru/mux34_b0_sel_is_2_o ),
    .o(\cu_ru/vec_pc [11]));
  binary_mux_s1_w1 \cu_ru/mux3_b0  (
    .i0(\cu_ru/n50 [0]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b1  (
    .i0(\cu_ru/n50 [1]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b10  (
    .i0(\cu_ru/n50 [10]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b11  (
    .i0(\cu_ru/n50 [11]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b12  (
    .i0(\cu_ru/n50 [12]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b13  (
    .i0(\cu_ru/n50 [13]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b14  (
    .i0(\cu_ru/n50 [14]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b15  (
    .i0(\cu_ru/n50 [15]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b16  (
    .i0(\cu_ru/n50 [16]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b17  (
    .i0(\cu_ru/n50 [17]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b18  (
    .i0(\cu_ru/n50 [18]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b19  (
    .i0(\cu_ru/n50 [19]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b2  (
    .i0(\cu_ru/n50 [2]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b20  (
    .i0(\cu_ru/n50 [20]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b21  (
    .i0(\cu_ru/n50 [21]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b22  (
    .i0(\cu_ru/n50 [22]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b23  (
    .i0(\cu_ru/n50 [23]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b24  (
    .i0(\cu_ru/n50 [24]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b25  (
    .i0(\cu_ru/n50 [25]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b26  (
    .i0(\cu_ru/n50 [26]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b27  (
    .i0(\cu_ru/n50 [27]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b28  (
    .i0(\cu_ru/n50 [28]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b29  (
    .i0(\cu_ru/n50 [29]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b3  (
    .i0(\cu_ru/n50 [3]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b30  (
    .i0(\cu_ru/n50 [30]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b31  (
    .i0(\cu_ru/n50 [31]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b32  (
    .i0(\cu_ru/n50 [32]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b33  (
    .i0(\cu_ru/n50 [33]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b34  (
    .i0(\cu_ru/n50 [34]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b35  (
    .i0(\cu_ru/n50 [35]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b36  (
    .i0(\cu_ru/n50 [36]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b37  (
    .i0(\cu_ru/n50 [37]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b38  (
    .i0(\cu_ru/n50 [38]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b39  (
    .i0(\cu_ru/n50 [39]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b4  (
    .i0(\cu_ru/n50 [4]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b40  (
    .i0(\cu_ru/n50 [40]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b41  (
    .i0(\cu_ru/n50 [41]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b42  (
    .i0(\cu_ru/n50 [42]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b43  (
    .i0(\cu_ru/n50 [43]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b44  (
    .i0(\cu_ru/n50 [44]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b45  (
    .i0(\cu_ru/n50 [45]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b46  (
    .i0(\cu_ru/n50 [46]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b47  (
    .i0(\cu_ru/n50 [47]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b48  (
    .i0(\cu_ru/n50 [48]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b49  (
    .i0(\cu_ru/n50 [49]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b5  (
    .i0(\cu_ru/n50 [5]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b50  (
    .i0(\cu_ru/n50 [50]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b51  (
    .i0(\cu_ru/n50 [51]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b52  (
    .i0(\cu_ru/n50 [52]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b53  (
    .i0(\cu_ru/n50 [53]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b54  (
    .i0(\cu_ru/n50 [54]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b55  (
    .i0(\cu_ru/n50 [55]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b56  (
    .i0(\cu_ru/n50 [56]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b57  (
    .i0(\cu_ru/n50 [57]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b58  (
    .i0(\cu_ru/n50 [58]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b59  (
    .i0(\cu_ru/n50 [59]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b6  (
    .i0(\cu_ru/n50 [6]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b60  (
    .i0(\cu_ru/n50 [60]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b61  (
    .i0(\cu_ru/n50 [61]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b62  (
    .i0(\cu_ru/n50 [62]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b63  (
    .i0(\cu_ru/n50 [63]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b7  (
    .i0(\cu_ru/n50 [7]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b8  (
    .i0(\cu_ru/n50 [8]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux3_b9  (
    .i0(\cu_ru/n50 [9]),
    .i1(1'b0),
    .sel(\cu_ru/n48 ),
    .o(rs2_data[9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  binary_mux_s1_w1 \cu_ru/mux4_b0  (
    .i0(new_pc[0]),
    .i1(\cu_ru/tvec [2]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b1  (
    .i0(new_pc[1]),
    .i1(\cu_ru/tvec [3]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b10  (
    .i0(new_pc[10]),
    .i1(\cu_ru/vec_pc [10]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b11  (
    .i0(new_pc[11]),
    .i1(\cu_ru/vec_pc [11]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b12  (
    .i0(new_pc[12]),
    .i1(\cu_ru/vec_pc [12]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b13  (
    .i0(new_pc[13]),
    .i1(\cu_ru/vec_pc [13]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b14  (
    .i0(new_pc[14]),
    .i1(\cu_ru/vec_pc [14]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b15  (
    .i0(new_pc[15]),
    .i1(\cu_ru/vec_pc [15]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b16  (
    .i0(new_pc[16]),
    .i1(\cu_ru/vec_pc [16]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b17  (
    .i0(new_pc[17]),
    .i1(\cu_ru/vec_pc [17]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b18  (
    .i0(new_pc[18]),
    .i1(\cu_ru/vec_pc [18]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b19  (
    .i0(new_pc[19]),
    .i1(\cu_ru/vec_pc [19]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b2  (
    .i0(new_pc[2]),
    .i1(\cu_ru/vec_pc [2]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b20  (
    .i0(new_pc[20]),
    .i1(\cu_ru/vec_pc [20]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b21  (
    .i0(new_pc[21]),
    .i1(\cu_ru/vec_pc [21]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b22  (
    .i0(new_pc[22]),
    .i1(\cu_ru/vec_pc [22]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b23  (
    .i0(new_pc[23]),
    .i1(\cu_ru/vec_pc [23]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b24  (
    .i0(new_pc[24]),
    .i1(\cu_ru/vec_pc [24]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b25  (
    .i0(new_pc[25]),
    .i1(\cu_ru/vec_pc [25]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b26  (
    .i0(new_pc[26]),
    .i1(\cu_ru/vec_pc [26]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b27  (
    .i0(new_pc[27]),
    .i1(\cu_ru/vec_pc [27]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b28  (
    .i0(new_pc[28]),
    .i1(\cu_ru/vec_pc [28]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b29  (
    .i0(new_pc[29]),
    .i1(\cu_ru/vec_pc [29]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b3  (
    .i0(new_pc[3]),
    .i1(\cu_ru/vec_pc [3]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b30  (
    .i0(new_pc[30]),
    .i1(\cu_ru/vec_pc [30]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b31  (
    .i0(new_pc[31]),
    .i1(\cu_ru/vec_pc [31]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b32  (
    .i0(new_pc[32]),
    .i1(\cu_ru/vec_pc [32]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b33  (
    .i0(new_pc[33]),
    .i1(\cu_ru/vec_pc [33]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b34  (
    .i0(new_pc[34]),
    .i1(\cu_ru/vec_pc [34]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b35  (
    .i0(new_pc[35]),
    .i1(\cu_ru/vec_pc [35]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b36  (
    .i0(new_pc[36]),
    .i1(\cu_ru/vec_pc [36]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b37  (
    .i0(new_pc[37]),
    .i1(\cu_ru/vec_pc [37]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b38  (
    .i0(new_pc[38]),
    .i1(\cu_ru/vec_pc [38]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b39  (
    .i0(new_pc[39]),
    .i1(\cu_ru/vec_pc [39]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b4  (
    .i0(new_pc[4]),
    .i1(\cu_ru/vec_pc [4]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b40  (
    .i0(new_pc[40]),
    .i1(\cu_ru/vec_pc [40]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b41  (
    .i0(new_pc[41]),
    .i1(\cu_ru/vec_pc [41]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b42  (
    .i0(new_pc[42]),
    .i1(\cu_ru/vec_pc [42]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b43  (
    .i0(new_pc[43]),
    .i1(\cu_ru/vec_pc [43]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b44  (
    .i0(new_pc[44]),
    .i1(\cu_ru/vec_pc [44]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b45  (
    .i0(new_pc[45]),
    .i1(\cu_ru/vec_pc [45]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b46  (
    .i0(new_pc[46]),
    .i1(\cu_ru/vec_pc [46]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b47  (
    .i0(new_pc[47]),
    .i1(\cu_ru/vec_pc [47]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b48  (
    .i0(new_pc[48]),
    .i1(\cu_ru/vec_pc [48]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b49  (
    .i0(new_pc[49]),
    .i1(\cu_ru/vec_pc [49]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b5  (
    .i0(new_pc[5]),
    .i1(\cu_ru/vec_pc [5]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b50  (
    .i0(new_pc[50]),
    .i1(\cu_ru/vec_pc [50]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b51  (
    .i0(new_pc[51]),
    .i1(\cu_ru/vec_pc [51]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b52  (
    .i0(new_pc[52]),
    .i1(\cu_ru/vec_pc [52]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b53  (
    .i0(new_pc[53]),
    .i1(\cu_ru/vec_pc [53]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b54  (
    .i0(new_pc[54]),
    .i1(\cu_ru/vec_pc [54]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b55  (
    .i0(new_pc[55]),
    .i1(\cu_ru/vec_pc [55]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b56  (
    .i0(new_pc[56]),
    .i1(\cu_ru/vec_pc [56]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b57  (
    .i0(new_pc[57]),
    .i1(\cu_ru/vec_pc [57]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b58  (
    .i0(new_pc[58]),
    .i1(\cu_ru/vec_pc [58]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b59  (
    .i0(new_pc[59]),
    .i1(\cu_ru/vec_pc [59]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b6  (
    .i0(new_pc[6]),
    .i1(\cu_ru/vec_pc [6]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b60  (
    .i0(new_pc[60]),
    .i1(\cu_ru/vec_pc [60]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b61  (
    .i0(new_pc[61]),
    .i1(\cu_ru/vec_pc [61]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b62  (
    .i0(new_pc[62]),
    .i1(\cu_ru/vec_pc [62]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b63  (
    .i0(new_pc[63]),
    .i1(1'b0),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b7  (
    .i0(new_pc[7]),
    .i1(\cu_ru/vec_pc [7]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b8  (
    .i0(new_pc[8]),
    .i1(\cu_ru/vec_pc [8]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux4_b9  (
    .i0(new_pc[9]),
    .i1(\cu_ru/vec_pc [9]),
    .sel(\cu_ru/n56 ),
    .o(\cu_ru/n57 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b0  (
    .i0(\cu_ru/n57 [0]),
    .i1(\cu_ru/sepc [0]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b1  (
    .i0(\cu_ru/n57 [1]),
    .i1(\cu_ru/sepc [1]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b10  (
    .i0(\cu_ru/n57 [10]),
    .i1(\cu_ru/sepc [10]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b11  (
    .i0(\cu_ru/n57 [11]),
    .i1(\cu_ru/sepc [11]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b12  (
    .i0(\cu_ru/n57 [12]),
    .i1(\cu_ru/sepc [12]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b13  (
    .i0(\cu_ru/n57 [13]),
    .i1(\cu_ru/sepc [13]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b14  (
    .i0(\cu_ru/n57 [14]),
    .i1(\cu_ru/sepc [14]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b15  (
    .i0(\cu_ru/n57 [15]),
    .i1(\cu_ru/sepc [15]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b16  (
    .i0(\cu_ru/n57 [16]),
    .i1(\cu_ru/sepc [16]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b17  (
    .i0(\cu_ru/n57 [17]),
    .i1(\cu_ru/sepc [17]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b18  (
    .i0(\cu_ru/n57 [18]),
    .i1(\cu_ru/sepc [18]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b19  (
    .i0(\cu_ru/n57 [19]),
    .i1(\cu_ru/sepc [19]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b2  (
    .i0(\cu_ru/n57 [2]),
    .i1(\cu_ru/sepc [2]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b20  (
    .i0(\cu_ru/n57 [20]),
    .i1(\cu_ru/sepc [20]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b21  (
    .i0(\cu_ru/n57 [21]),
    .i1(\cu_ru/sepc [21]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b22  (
    .i0(\cu_ru/n57 [22]),
    .i1(\cu_ru/sepc [22]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b23  (
    .i0(\cu_ru/n57 [23]),
    .i1(\cu_ru/sepc [23]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b24  (
    .i0(\cu_ru/n57 [24]),
    .i1(\cu_ru/sepc [24]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b25  (
    .i0(\cu_ru/n57 [25]),
    .i1(\cu_ru/sepc [25]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b26  (
    .i0(\cu_ru/n57 [26]),
    .i1(\cu_ru/sepc [26]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b27  (
    .i0(\cu_ru/n57 [27]),
    .i1(\cu_ru/sepc [27]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b28  (
    .i0(\cu_ru/n57 [28]),
    .i1(\cu_ru/sepc [28]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b29  (
    .i0(\cu_ru/n57 [29]),
    .i1(\cu_ru/sepc [29]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b3  (
    .i0(\cu_ru/n57 [3]),
    .i1(\cu_ru/sepc [3]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b30  (
    .i0(\cu_ru/n57 [30]),
    .i1(\cu_ru/sepc [30]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b31  (
    .i0(\cu_ru/n57 [31]),
    .i1(\cu_ru/sepc [31]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b32  (
    .i0(\cu_ru/n57 [32]),
    .i1(\cu_ru/sepc [32]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b33  (
    .i0(\cu_ru/n57 [33]),
    .i1(\cu_ru/sepc [33]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b34  (
    .i0(\cu_ru/n57 [34]),
    .i1(\cu_ru/sepc [34]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b35  (
    .i0(\cu_ru/n57 [35]),
    .i1(\cu_ru/sepc [35]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b36  (
    .i0(\cu_ru/n57 [36]),
    .i1(\cu_ru/sepc [36]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b37  (
    .i0(\cu_ru/n57 [37]),
    .i1(\cu_ru/sepc [37]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b38  (
    .i0(\cu_ru/n57 [38]),
    .i1(\cu_ru/sepc [38]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b39  (
    .i0(\cu_ru/n57 [39]),
    .i1(\cu_ru/sepc [39]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b4  (
    .i0(\cu_ru/n57 [4]),
    .i1(\cu_ru/sepc [4]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b40  (
    .i0(\cu_ru/n57 [40]),
    .i1(\cu_ru/sepc [40]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b41  (
    .i0(\cu_ru/n57 [41]),
    .i1(\cu_ru/sepc [41]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b42  (
    .i0(\cu_ru/n57 [42]),
    .i1(\cu_ru/sepc [42]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b43  (
    .i0(\cu_ru/n57 [43]),
    .i1(\cu_ru/sepc [43]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b44  (
    .i0(\cu_ru/n57 [44]),
    .i1(\cu_ru/sepc [44]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b45  (
    .i0(\cu_ru/n57 [45]),
    .i1(\cu_ru/sepc [45]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b46  (
    .i0(\cu_ru/n57 [46]),
    .i1(\cu_ru/sepc [46]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b47  (
    .i0(\cu_ru/n57 [47]),
    .i1(\cu_ru/sepc [47]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b48  (
    .i0(\cu_ru/n57 [48]),
    .i1(\cu_ru/sepc [48]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b49  (
    .i0(\cu_ru/n57 [49]),
    .i1(\cu_ru/sepc [49]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b5  (
    .i0(\cu_ru/n57 [5]),
    .i1(\cu_ru/sepc [5]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b50  (
    .i0(\cu_ru/n57 [50]),
    .i1(\cu_ru/sepc [50]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b51  (
    .i0(\cu_ru/n57 [51]),
    .i1(\cu_ru/sepc [51]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b52  (
    .i0(\cu_ru/n57 [52]),
    .i1(\cu_ru/sepc [52]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b53  (
    .i0(\cu_ru/n57 [53]),
    .i1(\cu_ru/sepc [53]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b54  (
    .i0(\cu_ru/n57 [54]),
    .i1(\cu_ru/sepc [54]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b55  (
    .i0(\cu_ru/n57 [55]),
    .i1(\cu_ru/sepc [55]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b56  (
    .i0(\cu_ru/n57 [56]),
    .i1(\cu_ru/sepc [56]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b57  (
    .i0(\cu_ru/n57 [57]),
    .i1(\cu_ru/sepc [57]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b58  (
    .i0(\cu_ru/n57 [58]),
    .i1(\cu_ru/sepc [58]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b59  (
    .i0(\cu_ru/n57 [59]),
    .i1(\cu_ru/sepc [59]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b6  (
    .i0(\cu_ru/n57 [6]),
    .i1(\cu_ru/sepc [6]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b60  (
    .i0(\cu_ru/n57 [60]),
    .i1(\cu_ru/sepc [60]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b61  (
    .i0(\cu_ru/n57 [61]),
    .i1(\cu_ru/sepc [61]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b62  (
    .i0(\cu_ru/n57 [62]),
    .i1(\cu_ru/sepc [62]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b63  (
    .i0(\cu_ru/n57 [63]),
    .i1(\cu_ru/sepc [63]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b7  (
    .i0(\cu_ru/n57 [7]),
    .i1(\cu_ru/sepc [7]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b8  (
    .i0(\cu_ru/n57 [8]),
    .i1(\cu_ru/sepc [8]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux5_b9  (
    .i0(\cu_ru/n57 [9]),
    .i1(\cu_ru/sepc [9]),
    .sel(\cu_ru/m_s_status/n3 ),
    .o(\cu_ru/n58 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b0  (
    .i0(\cu_ru/n58 [0]),
    .i1(\cu_ru/mepc [0]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b1  (
    .i0(\cu_ru/n58 [1]),
    .i1(\cu_ru/mepc [1]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b10  (
    .i0(\cu_ru/n58 [10]),
    .i1(\cu_ru/mepc [10]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b11  (
    .i0(\cu_ru/n58 [11]),
    .i1(\cu_ru/mepc [11]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b12  (
    .i0(\cu_ru/n58 [12]),
    .i1(\cu_ru/mepc [12]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b13  (
    .i0(\cu_ru/n58 [13]),
    .i1(\cu_ru/mepc [13]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b14  (
    .i0(\cu_ru/n58 [14]),
    .i1(\cu_ru/mepc [14]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b15  (
    .i0(\cu_ru/n58 [15]),
    .i1(\cu_ru/mepc [15]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b16  (
    .i0(\cu_ru/n58 [16]),
    .i1(\cu_ru/mepc [16]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b17  (
    .i0(\cu_ru/n58 [17]),
    .i1(\cu_ru/mepc [17]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b18  (
    .i0(\cu_ru/n58 [18]),
    .i1(\cu_ru/mepc [18]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b19  (
    .i0(\cu_ru/n58 [19]),
    .i1(\cu_ru/mepc [19]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b2  (
    .i0(\cu_ru/n58 [2]),
    .i1(\cu_ru/mepc [2]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b20  (
    .i0(\cu_ru/n58 [20]),
    .i1(\cu_ru/mepc [20]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b21  (
    .i0(\cu_ru/n58 [21]),
    .i1(\cu_ru/mepc [21]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b22  (
    .i0(\cu_ru/n58 [22]),
    .i1(\cu_ru/mepc [22]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b23  (
    .i0(\cu_ru/n58 [23]),
    .i1(\cu_ru/mepc [23]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b24  (
    .i0(\cu_ru/n58 [24]),
    .i1(\cu_ru/mepc [24]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b25  (
    .i0(\cu_ru/n58 [25]),
    .i1(\cu_ru/mepc [25]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b26  (
    .i0(\cu_ru/n58 [26]),
    .i1(\cu_ru/mepc [26]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b27  (
    .i0(\cu_ru/n58 [27]),
    .i1(\cu_ru/mepc [27]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b28  (
    .i0(\cu_ru/n58 [28]),
    .i1(\cu_ru/mepc [28]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b29  (
    .i0(\cu_ru/n58 [29]),
    .i1(\cu_ru/mepc [29]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b3  (
    .i0(\cu_ru/n58 [3]),
    .i1(\cu_ru/mepc [3]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b30  (
    .i0(\cu_ru/n58 [30]),
    .i1(\cu_ru/mepc [30]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b31  (
    .i0(\cu_ru/n58 [31]),
    .i1(\cu_ru/mepc [31]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b32  (
    .i0(\cu_ru/n58 [32]),
    .i1(\cu_ru/mepc [32]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b33  (
    .i0(\cu_ru/n58 [33]),
    .i1(\cu_ru/mepc [33]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b34  (
    .i0(\cu_ru/n58 [34]),
    .i1(\cu_ru/mepc [34]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b35  (
    .i0(\cu_ru/n58 [35]),
    .i1(\cu_ru/mepc [35]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b36  (
    .i0(\cu_ru/n58 [36]),
    .i1(\cu_ru/mepc [36]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b37  (
    .i0(\cu_ru/n58 [37]),
    .i1(\cu_ru/mepc [37]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b38  (
    .i0(\cu_ru/n58 [38]),
    .i1(\cu_ru/mepc [38]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b39  (
    .i0(\cu_ru/n58 [39]),
    .i1(\cu_ru/mepc [39]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b4  (
    .i0(\cu_ru/n58 [4]),
    .i1(\cu_ru/mepc [4]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b40  (
    .i0(\cu_ru/n58 [40]),
    .i1(\cu_ru/mepc [40]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b41  (
    .i0(\cu_ru/n58 [41]),
    .i1(\cu_ru/mepc [41]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b42  (
    .i0(\cu_ru/n58 [42]),
    .i1(\cu_ru/mepc [42]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b43  (
    .i0(\cu_ru/n58 [43]),
    .i1(\cu_ru/mepc [43]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b44  (
    .i0(\cu_ru/n58 [44]),
    .i1(\cu_ru/mepc [44]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b45  (
    .i0(\cu_ru/n58 [45]),
    .i1(\cu_ru/mepc [45]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b46  (
    .i0(\cu_ru/n58 [46]),
    .i1(\cu_ru/mepc [46]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b47  (
    .i0(\cu_ru/n58 [47]),
    .i1(\cu_ru/mepc [47]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b48  (
    .i0(\cu_ru/n58 [48]),
    .i1(\cu_ru/mepc [48]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b49  (
    .i0(\cu_ru/n58 [49]),
    .i1(\cu_ru/mepc [49]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b5  (
    .i0(\cu_ru/n58 [5]),
    .i1(\cu_ru/mepc [5]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b50  (
    .i0(\cu_ru/n58 [50]),
    .i1(\cu_ru/mepc [50]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b51  (
    .i0(\cu_ru/n58 [51]),
    .i1(\cu_ru/mepc [51]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b52  (
    .i0(\cu_ru/n58 [52]),
    .i1(\cu_ru/mepc [52]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b53  (
    .i0(\cu_ru/n58 [53]),
    .i1(\cu_ru/mepc [53]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b54  (
    .i0(\cu_ru/n58 [54]),
    .i1(\cu_ru/mepc [54]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b55  (
    .i0(\cu_ru/n58 [55]),
    .i1(\cu_ru/mepc [55]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b56  (
    .i0(\cu_ru/n58 [56]),
    .i1(\cu_ru/mepc [56]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b57  (
    .i0(\cu_ru/n58 [57]),
    .i1(\cu_ru/mepc [57]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b58  (
    .i0(\cu_ru/n58 [58]),
    .i1(\cu_ru/mepc [58]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b59  (
    .i0(\cu_ru/n58 [59]),
    .i1(\cu_ru/mepc [59]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b6  (
    .i0(\cu_ru/n58 [6]),
    .i1(\cu_ru/mepc [6]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b60  (
    .i0(\cu_ru/n58 [60]),
    .i1(\cu_ru/mepc [60]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b61  (
    .i0(\cu_ru/n58 [61]),
    .i1(\cu_ru/mepc [61]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b62  (
    .i0(\cu_ru/n58 [62]),
    .i1(\cu_ru/mepc [62]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b63  (
    .i0(\cu_ru/n58 [63]),
    .i1(\cu_ru/mepc [63]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b7  (
    .i0(\cu_ru/n58 [7]),
    .i1(\cu_ru/mepc [7]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b8  (
    .i0(\cu_ru/n58 [8]),
    .i1(\cu_ru/mepc [8]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux6_b9  (
    .i0(\cu_ru/n58 [9]),
    .i1(\cu_ru/mepc [9]),
    .sel(\cu_ru/m_s_status/n2 ),
    .o(flush_pc[9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  binary_mux_s1_w1 \cu_ru/mux7_b0  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [0]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b1  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [1]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b10  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [10]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b11  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [11]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b12  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [12]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b13  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [13]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b14  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [14]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b15  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [15]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b16  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [16]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b17  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [17]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b18  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [18]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b19  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [19]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b2  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [2]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b20  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [20]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b21  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [21]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b22  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [22]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b23  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [23]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b24  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [24]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b25  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [25]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b26  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [26]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b27  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [27]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b28  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [28]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b29  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [29]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b3  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [3]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b30  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [30]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b31  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [31]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b32  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [32]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b33  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [33]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b34  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [34]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b35  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [35]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b36  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [36]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b37  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [37]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b38  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [38]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b39  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [39]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b4  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [4]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b40  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [40]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b41  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [41]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b42  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [42]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b43  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [43]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b44  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [44]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b45  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [45]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b46  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [46]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b47  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [47]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b48  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [48]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b49  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [49]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b5  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [5]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b50  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [50]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b51  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [51]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b52  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [52]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b53  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [53]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b54  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [54]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b55  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [55]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b56  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [56]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b57  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [57]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b58  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [58]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b59  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [59]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b6  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [6]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b60  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [60]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b61  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [61]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b62  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [62]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b63  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [63]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b7  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [7]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b8  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [8]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux7_b9  (
    .i0(1'b0),
    .i1(\cu_ru/mcycle [9]),
    .sel(\cu_ru/read_cycle_sel ),
    .o(\cu_ru/n59 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(672)
  binary_mux_s1_w1 \cu_ru/mux8_b0  (
    .i0(1'b0),
    .i1(mtime[0]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b1  (
    .i0(1'b0),
    .i1(mtime[1]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b10  (
    .i0(1'b0),
    .i1(mtime[10]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b11  (
    .i0(1'b0),
    .i1(mtime[11]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b12  (
    .i0(1'b0),
    .i1(mtime[12]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b13  (
    .i0(1'b0),
    .i1(mtime[13]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b14  (
    .i0(1'b0),
    .i1(mtime[14]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b15  (
    .i0(1'b0),
    .i1(mtime[15]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b16  (
    .i0(1'b0),
    .i1(mtime[16]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b17  (
    .i0(1'b0),
    .i1(mtime[17]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b18  (
    .i0(1'b0),
    .i1(mtime[18]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b19  (
    .i0(1'b0),
    .i1(mtime[19]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b2  (
    .i0(1'b0),
    .i1(mtime[2]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b20  (
    .i0(1'b0),
    .i1(mtime[20]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b21  (
    .i0(1'b0),
    .i1(mtime[21]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b22  (
    .i0(1'b0),
    .i1(mtime[22]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b23  (
    .i0(1'b0),
    .i1(mtime[23]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b24  (
    .i0(1'b0),
    .i1(mtime[24]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b25  (
    .i0(1'b0),
    .i1(mtime[25]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b26  (
    .i0(1'b0),
    .i1(mtime[26]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b27  (
    .i0(1'b0),
    .i1(mtime[27]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b28  (
    .i0(1'b0),
    .i1(mtime[28]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b29  (
    .i0(1'b0),
    .i1(mtime[29]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b3  (
    .i0(1'b0),
    .i1(mtime[3]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b30  (
    .i0(1'b0),
    .i1(mtime[30]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b31  (
    .i0(1'b0),
    .i1(mtime[31]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b32  (
    .i0(1'b0),
    .i1(mtime[32]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b33  (
    .i0(1'b0),
    .i1(mtime[33]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b34  (
    .i0(1'b0),
    .i1(mtime[34]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b35  (
    .i0(1'b0),
    .i1(mtime[35]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b36  (
    .i0(1'b0),
    .i1(mtime[36]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b37  (
    .i0(1'b0),
    .i1(mtime[37]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b38  (
    .i0(1'b0),
    .i1(mtime[38]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b39  (
    .i0(1'b0),
    .i1(mtime[39]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b4  (
    .i0(1'b0),
    .i1(mtime[4]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b40  (
    .i0(1'b0),
    .i1(mtime[40]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b41  (
    .i0(1'b0),
    .i1(mtime[41]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b42  (
    .i0(1'b0),
    .i1(mtime[42]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b43  (
    .i0(1'b0),
    .i1(mtime[43]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b44  (
    .i0(1'b0),
    .i1(mtime[44]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b45  (
    .i0(1'b0),
    .i1(mtime[45]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b46  (
    .i0(1'b0),
    .i1(mtime[46]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b47  (
    .i0(1'b0),
    .i1(mtime[47]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b48  (
    .i0(1'b0),
    .i1(mtime[48]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b49  (
    .i0(1'b0),
    .i1(mtime[49]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b5  (
    .i0(1'b0),
    .i1(mtime[5]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b50  (
    .i0(1'b0),
    .i1(mtime[50]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b51  (
    .i0(1'b0),
    .i1(mtime[51]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b52  (
    .i0(1'b0),
    .i1(mtime[52]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b53  (
    .i0(1'b0),
    .i1(mtime[53]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b54  (
    .i0(1'b0),
    .i1(mtime[54]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b55  (
    .i0(1'b0),
    .i1(mtime[55]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b56  (
    .i0(1'b0),
    .i1(mtime[56]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b57  (
    .i0(1'b0),
    .i1(mtime[57]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b58  (
    .i0(1'b0),
    .i1(mtime[58]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b59  (
    .i0(1'b0),
    .i1(mtime[59]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b6  (
    .i0(1'b0),
    .i1(mtime[6]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b60  (
    .i0(1'b0),
    .i1(mtime[60]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b61  (
    .i0(1'b0),
    .i1(mtime[61]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b62  (
    .i0(1'b0),
    .i1(mtime[62]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b63  (
    .i0(1'b0),
    .i1(mtime[63]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b7  (
    .i0(1'b0),
    .i1(mtime[7]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b8  (
    .i0(1'b0),
    .i1(mtime[8]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux8_b9  (
    .i0(1'b0),
    .i1(mtime[9]),
    .sel(\cu_ru/read_time_sel ),
    .o(\cu_ru/n60 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  binary_mux_s1_w1 \cu_ru/mux9_b0  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [0]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [0]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b1  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [1]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [1]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b10  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [10]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [10]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b11  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [11]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [11]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b12  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [12]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [12]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b13  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [13]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [13]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b14  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [14]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [14]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b15  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [15]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [15]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b16  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [16]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [16]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b17  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [17]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [17]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b18  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [18]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [18]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b19  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [19]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [19]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b2  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [2]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [2]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b20  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [20]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [20]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b21  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [21]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [21]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b22  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [22]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [22]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b23  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [23]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [23]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b24  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [24]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [24]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b25  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [25]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [25]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b26  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [26]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [26]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b27  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [27]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [27]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b28  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [28]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [28]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b29  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [29]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [29]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b3  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [3]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [3]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b30  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [30]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [30]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b31  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [31]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [31]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b32  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [32]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [32]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b33  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [33]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [33]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b34  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [34]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [34]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b35  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [35]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [35]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b36  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [36]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [36]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b37  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [37]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [37]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b38  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [38]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [38]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b39  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [39]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [39]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b4  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [4]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [4]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b40  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [40]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [40]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b41  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [41]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [41]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b42  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [42]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [42]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b43  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [43]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [43]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b44  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [44]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [44]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b45  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [45]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [45]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b46  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [46]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [46]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b47  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [47]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [47]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b48  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [48]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [48]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b49  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [49]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [49]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b5  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [5]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [5]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b50  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [50]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [50]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b51  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [51]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [51]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b52  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [52]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [52]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b53  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [53]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [53]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b54  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [54]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [54]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b55  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [55]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [55]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b56  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [56]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [56]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b57  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [57]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [57]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b58  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [58]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [58]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b59  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [59]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [59]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b6  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [6]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [6]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b60  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [60]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [60]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b61  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [61]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [61]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b62  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [62]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [62]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b63  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [63]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [63]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b7  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [7]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [7]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b8  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [8]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [8]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  binary_mux_s1_w1 \cu_ru/mux9_b9  (
    .i0(1'b0),
    .i1(\cu_ru/minstret [9]),
    .sel(\cu_ru/read_instret_sel ),
    .o(\cu_ru/n62 [9]));  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  ne_w5 \cu_ru/neq0  (
    .i0(wb_rd_index),
    .i1(5'b00000),
    .o(\cu_ru/n51 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(368)
  add_pu5_mu5_o5 \cu_ru/sub0  (
    .i0(id_rs1_index),
    .i1(5'b00001),
    .o(\cu_ru/n46 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(363)
  add_pu5_mu5_o5 \cu_ru/sub1  (
    .i0(id_rs2_index),
    .i1(5'b00001),
    .o(\cu_ru/n49 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(364)
  add_pu5_mu5_o5 \cu_ru/sub2  (
    .i0(wb_rd_index),
    .i1(5'b00001),
    .o(\cu_ru/n52 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(369)
  not \cu_ru/trap_target_m_inv  (\cu_ru/trap_target_m_neg , \cu_ru/trap_target_m );
  not \cu_ru/trap_target_s_inv  (\cu_ru/trap_target_s_neg , \cu_ru/trap_target_s );
  and \cu_ru/u10  (\cu_ru/srw_satp_sel , wb_valid, \cu_ru/n8 );  // ../../RTL/CPU/CU&RU/cu_ru.v(273)
  or \cu_ru/u100  (csr_data[52], \cu_ru/n113 [52], \cu_ru/n114 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u101  (csr_data[53], \cu_ru/n113 [53], \cu_ru/n114 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u102  (csr_data[54], \cu_ru/n113 [54], \cu_ru/n114 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u103  (csr_data[55], \cu_ru/n113 [55], \cu_ru/n114 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u1033  (\cu_ru/n83 [2], \cu_ru/n81 [2], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u1035  (\cu_ru/n83 [4], \cu_ru/n81 [4], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u1037  (\cu_ru/n83 [6], \cu_ru/n81 [6], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u1039  (\cu_ru/n83 [8], \cu_ru/n81 [8], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u104  (csr_data[56], \cu_ru/n113 [56], \cu_ru/n114 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u1045  (\cu_ru/n83 [14], \cu_ru/n81 [14], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u1048  (\cu_ru/n83 [17], \cu_ru/n81 [17], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u1049  (\cu_ru/n83 [18], \cu_ru/n81 [18], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u105  (csr_data[57], \cu_ru/n113 [57], \cu_ru/n114 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u1051  (\cu_ru/n83 [20], \cu_ru/n81 [20], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u1053  (\cu_ru/n83 [22], \cu_ru/n81 [22], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u1056  (\cu_ru/n83 [25], \cu_ru/n81 [25], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u1059  (\cu_ru/n83 [28], \cu_ru/n81 [28], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u106  (csr_data[58], \cu_ru/n113 [58], \cu_ru/n114 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u1061  (\cu_ru/n83 [30], \cu_ru/n81 [30], \cu_ru/n82 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(686)
  or \cu_ru/u107  (csr_data[59], \cu_ru/n113 [59], \cu_ru/n114 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u108  (csr_data[60], \cu_ru/n113 [60], \cu_ru/n114 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u109  (csr_data[61], \cu_ru/n113 [61], \cu_ru/n114 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u1095  (\cu_ru/n81 [1], \cu_ru/n79 [1], \cu_ru/n80 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1096  (\cu_ru/n81 [2], \cu_ru/n77 [2], \cu_ru/n80 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1097  (\cu_ru/n81 [3], \cu_ru/n77 [3], \cu_ru/n80 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1098  (\cu_ru/n81 [4], \cu_ru/n77 [4], \cu_ru/n80 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1099  (\cu_ru/n81 [5], \cu_ru/n79 [5], \cu_ru/n80 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  and \cu_ru/u11  (\cu_ru/mrw_mstatus_sel , wb_valid, \cu_ru/n9 );  // ../../RTL/CPU/CU&RU/cu_ru.v(278)
  or \cu_ru/u110  (csr_data[62], \cu_ru/n113 [62], \cu_ru/n114 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u1100  (\cu_ru/n81 [6], \cu_ru/n77 [6], \cu_ru/n80 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1101  (\cu_ru/n81 [7], \cu_ru/n77 [7], \cu_ru/n80 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1102  (\cu_ru/n81 [8], \cu_ru/n77 [8], \cu_ru/n80 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1103  (\cu_ru/n81 [9], \cu_ru/n79 [9], \cu_ru/n80 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1104  (\cu_ru/n81 [10], \cu_ru/n77 [10], \cu_ru/n80 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1105  (\cu_ru/n81 [11], \cu_ru/n77 [11], \cu_ru/n80 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1106  (\cu_ru/n81 [12], \cu_ru/n77 [12], \cu_ru/n80 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1107  (\cu_ru/n81 [13], \cu_ru/n77 [13], \cu_ru/n80 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1108  (\cu_ru/n81 [14], \cu_ru/n77 [14], \cu_ru/n80 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1109  (\cu_ru/n81 [15], \cu_ru/n77 [15], \cu_ru/n80 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u111  (csr_data[63], \cu_ru/n113 [63], \cu_ru/n114 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u1110  (\cu_ru/n81 [16], \cu_ru/n77 [16], \cu_ru/n80 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1111  (\cu_ru/n81 [17], \cu_ru/n77 [17], \cu_ru/n80 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1112  (\cu_ru/n81 [18], \cu_ru/n77 [18], \cu_ru/n80 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1113  (\cu_ru/n81 [19], \cu_ru/n77 [19], \cu_ru/n80 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1114  (\cu_ru/n81 [20], \cu_ru/n77 [20], \cu_ru/n80 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1115  (\cu_ru/n81 [21], \cu_ru/n77 [21], \cu_ru/n80 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1116  (\cu_ru/n81 [22], \cu_ru/n77 [22], \cu_ru/n80 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1117  (\cu_ru/n81 [23], \cu_ru/n77 [23], \cu_ru/n80 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1118  (\cu_ru/n81 [24], \cu_ru/n77 [24], \cu_ru/n80 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1119  (\cu_ru/n81 [25], \cu_ru/n77 [25], \cu_ru/n80 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u112  (\cu_ru/n113 [1], \cu_ru/n111 [1], \cu_ru/n112 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1120  (\cu_ru/n81 [26], \cu_ru/n77 [26], \cu_ru/n80 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1121  (\cu_ru/n81 [27], \cu_ru/n77 [27], \cu_ru/n80 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1122  (\cu_ru/n81 [28], \cu_ru/n77 [28], \cu_ru/n80 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1123  (\cu_ru/n81 [29], \cu_ru/n77 [29], \cu_ru/n80 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1124  (\cu_ru/n81 [30], \cu_ru/n77 [30], \cu_ru/n80 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1125  (\cu_ru/n81 [31], \cu_ru/n77 [31], \cu_ru/n80 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1126  (\cu_ru/n81 [32], \cu_ru/n77 [32], \cu_ru/n80 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1127  (\cu_ru/n81 [33], \cu_ru/n77 [33], \cu_ru/n80 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1128  (\cu_ru/n81 [34], \cu_ru/n77 [34], \cu_ru/n80 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1129  (\cu_ru/n81 [35], \cu_ru/n77 [35], \cu_ru/n80 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u113  (\cu_ru/n113 [2], \cu_ru/n109 [2], \cu_ru/n112 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1130  (\cu_ru/n81 [36], \cu_ru/n77 [36], \cu_ru/n80 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1131  (\cu_ru/n81 [37], \cu_ru/n77 [37], \cu_ru/n80 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1132  (\cu_ru/n81 [38], \cu_ru/n77 [38], \cu_ru/n80 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1133  (\cu_ru/n81 [39], \cu_ru/n77 [39], \cu_ru/n80 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1134  (\cu_ru/n81 [40], \cu_ru/n77 [40], \cu_ru/n80 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1135  (\cu_ru/n81 [41], \cu_ru/n77 [41], \cu_ru/n80 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1136  (\cu_ru/n81 [42], \cu_ru/n77 [42], \cu_ru/n80 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1137  (\cu_ru/n81 [43], \cu_ru/n77 [43], \cu_ru/n80 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u114  (\cu_ru/n113 [3], \cu_ru/n111 [3], \cu_ru/n112 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u115  (\cu_ru/n113 [4], \cu_ru/n109 [4], \cu_ru/n112 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1154  (\cu_ru/n81 [60], \cu_ru/n77 [60], \cu_ru/n80 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1155  (\cu_ru/n81 [61], \cu_ru/n77 [61], \cu_ru/n80 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1156  (\cu_ru/n81 [62], \cu_ru/n77 [62], \cu_ru/n80 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1157  (\cu_ru/n81 [63], \cu_ru/n77 [63], \cu_ru/n80 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  or \cu_ru/u1158  (\cu_ru/n79 [1], \cu_ru/n77 [1], \cu_ru/n78 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(684)
  or \cu_ru/u116  (\cu_ru/n113 [5], \cu_ru/n111 [5], \cu_ru/n112 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1162  (\cu_ru/n79 [5], \cu_ru/n77 [5], \cu_ru/n78 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(684)
  or \cu_ru/u1166  (\cu_ru/n79 [9], \cu_ru/n77 [9], \cu_ru/n78 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(684)
  or \cu_ru/u117  (\cu_ru/n113 [6], \cu_ru/n109 [6], \cu_ru/n112 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u118  (\cu_ru/n113 [7], \cu_ru/n111 [7], \cu_ru/n112 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u119  (\cu_ru/n113 [8], \cu_ru/n109 [8], \cu_ru/n112 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  and \cu_ru/u12  (\cu_ru/mrw_medeleg_sel , wb_valid, \cu_ru/n10 );  // ../../RTL/CPU/CU&RU/cu_ru.v(280)
  or \cu_ru/u120  (\cu_ru/n113 [9], \cu_ru/n111 [9], \cu_ru/n112 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u121  (\cu_ru/n113 [10], \cu_ru/n109 [10], \cu_ru/n112 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u122  (\cu_ru/n113 [11], \cu_ru/n111 [11], \cu_ru/n112 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1221  (\cu_ru/n77 [1], \cu_ru/n75 [1], \cu_ru/n76 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1222  (\cu_ru/n77 [2], \cu_ru/n75 [2], \cu_ru/n76 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1223  (\cu_ru/n77 [3], \cu_ru/n75 [3], \cu_ru/n76 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1224  (\cu_ru/n77 [4], \cu_ru/n75 [4], \cu_ru/n76 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1225  (\cu_ru/n77 [5], \cu_ru/n75 [5], \cu_ru/n76 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1226  (\cu_ru/n77 [6], \cu_ru/n75 [6], \cu_ru/n76 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1227  (\cu_ru/n77 [7], \cu_ru/n75 [7], \cu_ru/n76 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1228  (\cu_ru/n77 [8], \cu_ru/n75 [8], \cu_ru/n76 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1229  (\cu_ru/n77 [9], \cu_ru/n75 [9], \cu_ru/n76 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u123  (\cu_ru/n113 [12], \cu_ru/n109 [12], \cu_ru/n112 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1230  (\cu_ru/n77 [10], \cu_ru/n75 [10], \cu_ru/n76 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1231  (\cu_ru/n77 [11], \cu_ru/n75 [11], \cu_ru/n76 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1232  (\cu_ru/n77 [12], \cu_ru/n75 [12], \cu_ru/n76 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1233  (\cu_ru/n77 [13], \cu_ru/n75 [13], \cu_ru/n76 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1234  (\cu_ru/n77 [14], \cu_ru/n75 [14], \cu_ru/n76 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1235  (\cu_ru/n77 [15], \cu_ru/n75 [15], \cu_ru/n76 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1236  (\cu_ru/n77 [16], \cu_ru/n75 [16], \cu_ru/n76 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1237  (\cu_ru/n77 [17], \cu_ru/n75 [17], \cu_ru/n76 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1238  (\cu_ru/n77 [18], \cu_ru/n75 [18], \cu_ru/n76 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1239  (\cu_ru/n77 [19], \cu_ru/n75 [19], \cu_ru/n76 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u124  (\cu_ru/n113 [13], \cu_ru/n109 [13], \cu_ru/n112 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1240  (\cu_ru/n77 [20], \cu_ru/n75 [20], \cu_ru/n76 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1241  (\cu_ru/n77 [21], \cu_ru/n75 [21], \cu_ru/n76 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1242  (\cu_ru/n77 [22], \cu_ru/n75 [22], \cu_ru/n76 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1243  (\cu_ru/n77 [23], \cu_ru/n75 [23], \cu_ru/n76 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1244  (\cu_ru/n77 [24], \cu_ru/n75 [24], \cu_ru/n76 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1245  (\cu_ru/n77 [25], \cu_ru/n75 [25], \cu_ru/n76 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1246  (\cu_ru/n77 [26], \cu_ru/n75 [26], \cu_ru/n76 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1247  (\cu_ru/n77 [27], \cu_ru/n75 [27], \cu_ru/n76 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1248  (\cu_ru/n77 [28], \cu_ru/n75 [28], \cu_ru/n76 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1249  (\cu_ru/n77 [29], \cu_ru/n75 [29], \cu_ru/n76 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u125  (\cu_ru/n113 [14], \cu_ru/n109 [14], \cu_ru/n112 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1250  (\cu_ru/n77 [30], \cu_ru/n75 [30], \cu_ru/n76 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1251  (\cu_ru/n77 [31], \cu_ru/n75 [31], \cu_ru/n76 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1252  (\cu_ru/n77 [32], \cu_ru/n75 [32], \cu_ru/n76 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1253  (\cu_ru/n77 [33], \cu_ru/n75 [33], \cu_ru/n76 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1254  (\cu_ru/n77 [34], \cu_ru/n75 [34], \cu_ru/n76 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1255  (\cu_ru/n77 [35], \cu_ru/n75 [35], \cu_ru/n76 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1256  (\cu_ru/n77 [36], \cu_ru/n75 [36], \cu_ru/n76 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1257  (\cu_ru/n77 [37], \cu_ru/n75 [37], \cu_ru/n76 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1258  (\cu_ru/n77 [38], \cu_ru/n75 [38], \cu_ru/n76 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1259  (\cu_ru/n77 [39], \cu_ru/n75 [39], \cu_ru/n76 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u126  (\cu_ru/n113 [15], \cu_ru/n109 [15], \cu_ru/n112 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1260  (\cu_ru/n77 [40], \cu_ru/n75 [40], \cu_ru/n76 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1261  (\cu_ru/n77 [41], \cu_ru/n75 [41], \cu_ru/n76 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1262  (\cu_ru/n77 [42], \cu_ru/n75 [42], \cu_ru/n76 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1263  (\cu_ru/n77 [43], \cu_ru/n75 [43], \cu_ru/n76 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1264  (\cu_ru/n77 [44], \cu_ru/n75 [44], \cu_ru/n76 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1265  (\cu_ru/n77 [45], \cu_ru/n75 [45], \cu_ru/n76 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1266  (\cu_ru/n77 [46], \cu_ru/n75 [46], \cu_ru/n76 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1267  (\cu_ru/n77 [47], \cu_ru/n75 [47], \cu_ru/n76 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1268  (\cu_ru/n77 [48], \cu_ru/n75 [48], \cu_ru/n76 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1269  (\cu_ru/n77 [49], \cu_ru/n75 [49], \cu_ru/n76 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u127  (\cu_ru/n113 [16], \cu_ru/n109 [16], \cu_ru/n112 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1270  (\cu_ru/n77 [50], \cu_ru/n75 [50], \cu_ru/n76 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1271  (\cu_ru/n77 [51], \cu_ru/n75 [51], \cu_ru/n76 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1272  (\cu_ru/n77 [52], \cu_ru/n75 [52], \cu_ru/n76 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1273  (\cu_ru/n77 [53], \cu_ru/n75 [53], \cu_ru/n76 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1274  (\cu_ru/n77 [54], \cu_ru/n75 [54], \cu_ru/n76 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1275  (\cu_ru/n77 [55], \cu_ru/n75 [55], \cu_ru/n76 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1276  (\cu_ru/n77 [56], \cu_ru/n75 [56], \cu_ru/n76 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1277  (\cu_ru/n77 [57], \cu_ru/n75 [57], \cu_ru/n76 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1278  (\cu_ru/n77 [58], \cu_ru/n75 [58], \cu_ru/n76 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1279  (\cu_ru/n77 [59], \cu_ru/n75 [59], \cu_ru/n76 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u128  (\cu_ru/n113 [17], \cu_ru/n109 [17], \cu_ru/n112 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1280  (\cu_ru/n77 [60], \cu_ru/n75 [60], \cu_ru/n76 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1281  (\cu_ru/n77 [61], \cu_ru/n75 [61], \cu_ru/n76 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1282  (\cu_ru/n77 [62], \cu_ru/n75 [62], \cu_ru/n76 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1283  (\cu_ru/n77 [63], \cu_ru/n75 [63], \cu_ru/n76 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1284  (\cu_ru/n75 [1], \cu_ru/n73 [1], \cu_ru/n74 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1285  (\cu_ru/n75 [2], \cu_ru/n73 [2], \cu_ru/n74 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1286  (\cu_ru/n75 [3], \cu_ru/n73 [3], \cu_ru/n74 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1287  (\cu_ru/n75 [4], \cu_ru/n73 [4], \cu_ru/n74 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1288  (\cu_ru/n75 [5], \cu_ru/n73 [5], \cu_ru/n74 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1289  (\cu_ru/n75 [6], \cu_ru/n73 [6], \cu_ru/n74 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u129  (\cu_ru/n113 [18], \cu_ru/n109 [18], \cu_ru/n112 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1290  (\cu_ru/n75 [7], \cu_ru/n73 [7], \cu_ru/n74 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1291  (\cu_ru/n75 [8], \cu_ru/n73 [8], \cu_ru/n74 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1292  (\cu_ru/n75 [9], \cu_ru/n73 [9], \cu_ru/n74 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1293  (\cu_ru/n75 [10], \cu_ru/n73 [10], \cu_ru/n74 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1294  (\cu_ru/n75 [11], \cu_ru/n73 [11], \cu_ru/n74 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1295  (\cu_ru/n75 [12], \cu_ru/n73 [12], \cu_ru/n74 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1296  (\cu_ru/n75 [13], \cu_ru/n73 [13], \cu_ru/n74 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1297  (\cu_ru/n75 [14], \cu_ru/n73 [14], \cu_ru/n74 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1298  (\cu_ru/n75 [15], \cu_ru/n73 [15], \cu_ru/n74 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1299  (\cu_ru/n75 [16], \cu_ru/n73 [16], \cu_ru/n74 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  and \cu_ru/u13  (\cu_ru/mrw_mideleg_sel , wb_valid, \cu_ru/n11 );  // ../../RTL/CPU/CU&RU/cu_ru.v(281)
  or \cu_ru/u130  (\cu_ru/n113 [19], \cu_ru/n109 [19], \cu_ru/n112 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1300  (\cu_ru/n75 [17], \cu_ru/n73 [17], \cu_ru/n74 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1301  (\cu_ru/n75 [18], \cu_ru/n73 [18], \cu_ru/n74 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1302  (\cu_ru/n75 [19], \cu_ru/n73 [19], \cu_ru/n74 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1303  (\cu_ru/n75 [20], \cu_ru/n73 [20], \cu_ru/n74 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1304  (\cu_ru/n75 [21], \cu_ru/n73 [21], \cu_ru/n74 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1305  (\cu_ru/n75 [22], \cu_ru/n73 [22], \cu_ru/n74 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1306  (\cu_ru/n75 [23], \cu_ru/n73 [23], \cu_ru/n74 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1307  (\cu_ru/n75 [24], \cu_ru/n73 [24], \cu_ru/n74 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1308  (\cu_ru/n75 [25], \cu_ru/n73 [25], \cu_ru/n74 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1309  (\cu_ru/n75 [26], \cu_ru/n73 [26], \cu_ru/n74 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u131  (\cu_ru/n113 [20], \cu_ru/n109 [20], \cu_ru/n112 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1310  (\cu_ru/n75 [27], \cu_ru/n73 [27], \cu_ru/n74 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1311  (\cu_ru/n75 [28], \cu_ru/n73 [28], \cu_ru/n74 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1312  (\cu_ru/n75 [29], \cu_ru/n73 [29], \cu_ru/n74 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1313  (\cu_ru/n75 [30], \cu_ru/n73 [30], \cu_ru/n74 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1314  (\cu_ru/n75 [31], \cu_ru/n73 [31], \cu_ru/n74 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1315  (\cu_ru/n75 [32], \cu_ru/n73 [32], \cu_ru/n74 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1316  (\cu_ru/n75 [33], \cu_ru/n73 [33], \cu_ru/n74 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1317  (\cu_ru/n75 [34], \cu_ru/n73 [34], \cu_ru/n74 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1318  (\cu_ru/n75 [35], \cu_ru/n73 [35], \cu_ru/n74 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1319  (\cu_ru/n75 [36], \cu_ru/n73 [36], \cu_ru/n74 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u132  (\cu_ru/n113 [21], \cu_ru/n109 [21], \cu_ru/n112 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1320  (\cu_ru/n75 [37], \cu_ru/n73 [37], \cu_ru/n74 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1321  (\cu_ru/n75 [38], \cu_ru/n73 [38], \cu_ru/n74 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1322  (\cu_ru/n75 [39], \cu_ru/n73 [39], \cu_ru/n74 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1323  (\cu_ru/n75 [40], \cu_ru/n73 [40], \cu_ru/n74 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1324  (\cu_ru/n75 [41], \cu_ru/n73 [41], \cu_ru/n74 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1325  (\cu_ru/n75 [42], \cu_ru/n73 [42], \cu_ru/n74 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1326  (\cu_ru/n75 [43], \cu_ru/n73 [43], \cu_ru/n74 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1327  (\cu_ru/n75 [44], \cu_ru/n73 [44], \cu_ru/n74 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1328  (\cu_ru/n75 [45], \cu_ru/n73 [45], \cu_ru/n74 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1329  (\cu_ru/n75 [46], \cu_ru/n73 [46], \cu_ru/n74 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u133  (\cu_ru/n113 [22], \cu_ru/n109 [22], \cu_ru/n112 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1330  (\cu_ru/n75 [47], \cu_ru/n73 [47], \cu_ru/n74 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1331  (\cu_ru/n75 [48], \cu_ru/n73 [48], \cu_ru/n74 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1332  (\cu_ru/n75 [49], \cu_ru/n73 [49], \cu_ru/n74 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1333  (\cu_ru/n75 [50], \cu_ru/n73 [50], \cu_ru/n74 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1334  (\cu_ru/n75 [51], \cu_ru/n73 [51], \cu_ru/n74 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1335  (\cu_ru/n75 [52], \cu_ru/n73 [52], \cu_ru/n74 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1336  (\cu_ru/n75 [53], \cu_ru/n73 [53], \cu_ru/n74 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1337  (\cu_ru/n75 [54], \cu_ru/n73 [54], \cu_ru/n74 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1338  (\cu_ru/n75 [55], \cu_ru/n73 [55], \cu_ru/n74 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1339  (\cu_ru/n75 [56], \cu_ru/n73 [56], \cu_ru/n74 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u134  (\cu_ru/n113 [23], \cu_ru/n109 [23], \cu_ru/n112 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1340  (\cu_ru/n75 [57], \cu_ru/n73 [57], \cu_ru/n74 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1341  (\cu_ru/n75 [58], \cu_ru/n73 [58], \cu_ru/n74 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1342  (\cu_ru/n75 [59], \cu_ru/n73 [59], \cu_ru/n74 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1343  (\cu_ru/n75 [60], \cu_ru/n73 [60], \cu_ru/n74 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1344  (\cu_ru/n75 [61], \cu_ru/n73 [61], \cu_ru/n74 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1345  (\cu_ru/n75 [62], \cu_ru/n73 [62], \cu_ru/n74 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1346  (\cu_ru/n75 [63], \cu_ru/n73 [63], \cu_ru/n74 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1347  (\cu_ru/n73 [1], \cu_ru/n71 [1], \cu_ru/n72 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1348  (\cu_ru/n73 [2], \cu_ru/n71 [2], \cu_ru/n72 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1349  (\cu_ru/n73 [3], \cu_ru/n71 [3], \cu_ru/n72 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u135  (\cu_ru/n113 [24], \cu_ru/n109 [24], \cu_ru/n112 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1350  (\cu_ru/n73 [4], \cu_ru/n71 [4], \cu_ru/n72 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1351  (\cu_ru/n73 [5], \cu_ru/n71 [5], \cu_ru/n72 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1352  (\cu_ru/n73 [6], \cu_ru/n71 [6], \cu_ru/n72 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1353  (\cu_ru/n73 [7], \cu_ru/n71 [7], \cu_ru/n72 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1354  (\cu_ru/n73 [8], \cu_ru/n71 [8], \cu_ru/n72 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1355  (\cu_ru/n73 [9], \cu_ru/n71 [9], \cu_ru/n72 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1356  (\cu_ru/n73 [10], \cu_ru/n71 [10], \cu_ru/n72 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1357  (\cu_ru/n73 [11], \cu_ru/n71 [11], \cu_ru/n72 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1358  (\cu_ru/n73 [12], \cu_ru/n71 [12], \cu_ru/n72 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1359  (\cu_ru/n73 [13], \cu_ru/n71 [13], \cu_ru/n72 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u136  (\cu_ru/n113 [25], \cu_ru/n109 [25], \cu_ru/n112 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1360  (\cu_ru/n73 [14], \cu_ru/n71 [14], \cu_ru/n72 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1361  (\cu_ru/n73 [15], \cu_ru/n71 [15], \cu_ru/n72 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1362  (\cu_ru/n73 [16], \cu_ru/n71 [16], \cu_ru/n72 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1363  (\cu_ru/n73 [17], \cu_ru/n71 [17], \cu_ru/n72 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1364  (\cu_ru/n73 [18], \cu_ru/n71 [18], \cu_ru/n72 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1365  (\cu_ru/n73 [19], \cu_ru/n71 [19], \cu_ru/n72 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1366  (\cu_ru/n73 [20], \cu_ru/n71 [20], \cu_ru/n72 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1367  (\cu_ru/n73 [21], \cu_ru/n71 [21], \cu_ru/n72 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1368  (\cu_ru/n73 [22], \cu_ru/n71 [22], \cu_ru/n72 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1369  (\cu_ru/n73 [23], \cu_ru/n71 [23], \cu_ru/n72 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u137  (\cu_ru/n113 [26], \cu_ru/n109 [26], \cu_ru/n112 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1370  (\cu_ru/n73 [24], \cu_ru/n71 [24], \cu_ru/n72 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1371  (\cu_ru/n73 [25], \cu_ru/n71 [25], \cu_ru/n72 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1372  (\cu_ru/n73 [26], \cu_ru/n71 [26], \cu_ru/n72 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1373  (\cu_ru/n73 [27], \cu_ru/n71 [27], \cu_ru/n72 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1374  (\cu_ru/n73 [28], \cu_ru/n71 [28], \cu_ru/n72 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1375  (\cu_ru/n73 [29], \cu_ru/n71 [29], \cu_ru/n72 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1376  (\cu_ru/n73 [30], \cu_ru/n71 [30], \cu_ru/n72 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1377  (\cu_ru/n73 [31], \cu_ru/n71 [31], \cu_ru/n72 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1378  (\cu_ru/n73 [32], \cu_ru/n71 [32], \cu_ru/n72 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1379  (\cu_ru/n73 [33], \cu_ru/n71 [33], \cu_ru/n72 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u138  (\cu_ru/n113 [27], \cu_ru/n109 [27], \cu_ru/n112 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1380  (\cu_ru/n73 [34], \cu_ru/n71 [34], \cu_ru/n72 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1381  (\cu_ru/n73 [35], \cu_ru/n71 [35], \cu_ru/n72 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1382  (\cu_ru/n73 [36], \cu_ru/n71 [36], \cu_ru/n72 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1383  (\cu_ru/n73 [37], \cu_ru/n71 [37], \cu_ru/n72 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1384  (\cu_ru/n73 [38], \cu_ru/n71 [38], \cu_ru/n72 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1385  (\cu_ru/n73 [39], \cu_ru/n71 [39], \cu_ru/n72 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1386  (\cu_ru/n73 [40], \cu_ru/n71 [40], \cu_ru/n72 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1387  (\cu_ru/n73 [41], \cu_ru/n71 [41], \cu_ru/n72 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1388  (\cu_ru/n73 [42], \cu_ru/n71 [42], \cu_ru/n72 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1389  (\cu_ru/n73 [43], \cu_ru/n71 [43], \cu_ru/n72 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u139  (\cu_ru/n113 [28], \cu_ru/n109 [28], \cu_ru/n112 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1390  (\cu_ru/n73 [44], \cu_ru/n71 [44], \cu_ru/n72 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1391  (\cu_ru/n73 [45], \cu_ru/n71 [45], \cu_ru/n72 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1392  (\cu_ru/n73 [46], \cu_ru/n71 [46], \cu_ru/n72 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1393  (\cu_ru/n73 [47], \cu_ru/n71 [47], \cu_ru/n72 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1394  (\cu_ru/n73 [48], \cu_ru/n71 [48], \cu_ru/n72 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1395  (\cu_ru/n73 [49], \cu_ru/n71 [49], \cu_ru/n72 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1396  (\cu_ru/n73 [50], \cu_ru/n71 [50], \cu_ru/n72 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1397  (\cu_ru/n73 [51], \cu_ru/n71 [51], \cu_ru/n72 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1398  (\cu_ru/n73 [52], \cu_ru/n71 [52], \cu_ru/n72 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1399  (\cu_ru/n73 [53], \cu_ru/n71 [53], \cu_ru/n72 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  and \cu_ru/u14  (\cu_ru/mrw_mie_sel , wb_valid, \cu_ru/n12 );  // ../../RTL/CPU/CU&RU/cu_ru.v(282)
  or \cu_ru/u140  (\cu_ru/n113 [29], \cu_ru/n109 [29], \cu_ru/n112 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1400  (\cu_ru/n73 [54], \cu_ru/n71 [54], \cu_ru/n72 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1401  (\cu_ru/n73 [55], \cu_ru/n71 [55], \cu_ru/n72 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1402  (\cu_ru/n73 [56], \cu_ru/n71 [56], \cu_ru/n72 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1403  (\cu_ru/n73 [57], \cu_ru/n71 [57], \cu_ru/n72 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1404  (\cu_ru/n73 [58], \cu_ru/n71 [58], \cu_ru/n72 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1405  (\cu_ru/n73 [59], \cu_ru/n71 [59], \cu_ru/n72 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1406  (\cu_ru/n73 [60], \cu_ru/n71 [60], \cu_ru/n72 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1407  (\cu_ru/n73 [61], \cu_ru/n71 [61], \cu_ru/n72 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1408  (\cu_ru/n73 [62], \cu_ru/n71 [62], \cu_ru/n72 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1409  (\cu_ru/n73 [63], \cu_ru/n71 [63], \cu_ru/n72 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u141  (\cu_ru/n113 [30], \cu_ru/n109 [30], \cu_ru/n112 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1410  (\cu_ru/n71 [1], \cu_ru/n69 [1], \cu_ru/n70 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1411  (\cu_ru/n71 [2], \cu_ru/n69 [2], \cu_ru/n70 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1412  (\cu_ru/n71 [3], \cu_ru/n69 [3], \cu_ru/n70 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1413  (\cu_ru/n71 [4], \cu_ru/n69 [4], \cu_ru/n70 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1414  (\cu_ru/n71 [5], \cu_ru/n69 [5], \cu_ru/n70 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1415  (\cu_ru/n71 [6], \cu_ru/n69 [6], \cu_ru/n70 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1416  (\cu_ru/n71 [7], \cu_ru/n69 [7], \cu_ru/n70 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1417  (\cu_ru/n71 [8], \cu_ru/n69 [8], \cu_ru/n70 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1418  (\cu_ru/n71 [9], \cu_ru/n69 [9], \cu_ru/n70 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1419  (\cu_ru/n71 [10], \cu_ru/n69 [10], \cu_ru/n70 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u142  (\cu_ru/n113 [31], \cu_ru/n109 [31], \cu_ru/n112 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1420  (\cu_ru/n71 [11], \cu_ru/n69 [11], \cu_ru/n70 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1421  (\cu_ru/n71 [12], \cu_ru/n69 [12], \cu_ru/n70 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1422  (\cu_ru/n71 [13], \cu_ru/n69 [13], \cu_ru/n70 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1423  (\cu_ru/n71 [14], \cu_ru/n69 [14], \cu_ru/n70 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1424  (\cu_ru/n71 [15], \cu_ru/n69 [15], \cu_ru/n70 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1425  (\cu_ru/n71 [16], \cu_ru/n69 [16], \cu_ru/n70 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1426  (\cu_ru/n71 [17], \cu_ru/n69 [17], \cu_ru/n70 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1427  (\cu_ru/n71 [18], \cu_ru/n69 [18], \cu_ru/n70 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1428  (\cu_ru/n71 [19], \cu_ru/n69 [19], \cu_ru/n70 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1429  (\cu_ru/n71 [20], \cu_ru/n69 [20], \cu_ru/n70 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u143  (\cu_ru/n113 [32], \cu_ru/n109 [32], \cu_ru/n112 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1430  (\cu_ru/n71 [21], \cu_ru/n69 [21], \cu_ru/n70 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1431  (\cu_ru/n71 [22], \cu_ru/n69 [22], \cu_ru/n70 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1432  (\cu_ru/n71 [23], \cu_ru/n69 [23], \cu_ru/n70 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1433  (\cu_ru/n71 [24], \cu_ru/n69 [24], \cu_ru/n70 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1434  (\cu_ru/n71 [25], \cu_ru/n69 [25], \cu_ru/n70 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1435  (\cu_ru/n71 [26], \cu_ru/n69 [26], \cu_ru/n70 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1436  (\cu_ru/n71 [27], \cu_ru/n69 [27], \cu_ru/n70 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1437  (\cu_ru/n71 [28], \cu_ru/n69 [28], \cu_ru/n70 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1438  (\cu_ru/n71 [29], \cu_ru/n69 [29], \cu_ru/n70 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1439  (\cu_ru/n71 [30], \cu_ru/n69 [30], \cu_ru/n70 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u144  (\cu_ru/n113 [33], \cu_ru/n109 [33], \cu_ru/n112 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1440  (\cu_ru/n71 [31], \cu_ru/n69 [31], \cu_ru/n70 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1441  (\cu_ru/n71 [32], \cu_ru/n69 [32], \cu_ru/n70 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1442  (\cu_ru/n71 [33], \cu_ru/n69 [33], \cu_ru/n70 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1443  (\cu_ru/n71 [34], \cu_ru/n69 [34], \cu_ru/n70 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1444  (\cu_ru/n71 [35], \cu_ru/n69 [35], \cu_ru/n70 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1445  (\cu_ru/n71 [36], \cu_ru/n69 [36], \cu_ru/n70 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1446  (\cu_ru/n71 [37], \cu_ru/n69 [37], \cu_ru/n70 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1447  (\cu_ru/n71 [38], \cu_ru/n69 [38], \cu_ru/n70 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1448  (\cu_ru/n71 [39], \cu_ru/n69 [39], \cu_ru/n70 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1449  (\cu_ru/n71 [40], \cu_ru/n69 [40], \cu_ru/n70 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u145  (\cu_ru/n113 [34], \cu_ru/n109 [34], \cu_ru/n112 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1450  (\cu_ru/n71 [41], \cu_ru/n69 [41], \cu_ru/n70 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1451  (\cu_ru/n71 [42], \cu_ru/n69 [42], \cu_ru/n70 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1452  (\cu_ru/n71 [43], \cu_ru/n69 [43], \cu_ru/n70 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1453  (\cu_ru/n71 [44], \cu_ru/n69 [44], \cu_ru/n70 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1454  (\cu_ru/n71 [45], \cu_ru/n69 [45], \cu_ru/n70 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1455  (\cu_ru/n71 [46], \cu_ru/n69 [46], \cu_ru/n70 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1456  (\cu_ru/n71 [47], \cu_ru/n69 [47], \cu_ru/n70 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1457  (\cu_ru/n71 [48], \cu_ru/n69 [48], \cu_ru/n70 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1458  (\cu_ru/n71 [49], \cu_ru/n69 [49], \cu_ru/n70 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1459  (\cu_ru/n71 [50], \cu_ru/n69 [50], \cu_ru/n70 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u146  (\cu_ru/n113 [35], \cu_ru/n109 [35], \cu_ru/n112 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1460  (\cu_ru/n71 [51], \cu_ru/n69 [51], \cu_ru/n70 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1461  (\cu_ru/n71 [52], \cu_ru/n69 [52], \cu_ru/n70 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1462  (\cu_ru/n71 [53], \cu_ru/n69 [53], \cu_ru/n70 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1463  (\cu_ru/n71 [54], \cu_ru/n69 [54], \cu_ru/n70 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1464  (\cu_ru/n71 [55], \cu_ru/n69 [55], \cu_ru/n70 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1465  (\cu_ru/n71 [56], \cu_ru/n69 [56], \cu_ru/n70 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1466  (\cu_ru/n71 [57], \cu_ru/n69 [57], \cu_ru/n70 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1467  (\cu_ru/n71 [58], \cu_ru/n69 [58], \cu_ru/n70 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1468  (\cu_ru/n71 [59], \cu_ru/n69 [59], \cu_ru/n70 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1469  (\cu_ru/n71 [60], \cu_ru/n69 [60], \cu_ru/n70 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u147  (\cu_ru/n113 [36], \cu_ru/n109 [36], \cu_ru/n112 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1470  (\cu_ru/n71 [61], \cu_ru/n69 [61], \cu_ru/n70 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1471  (\cu_ru/n71 [62], \cu_ru/n69 [62], \cu_ru/n70 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1472  (\cu_ru/n71 [63], \cu_ru/n69 [63], \cu_ru/n70 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1473  (\cu_ru/n69 [1], \cu_ru/n65 [1], \cu_ru/n68 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1474  (\cu_ru/n69 [2], \cu_ru/n63 [2], \cu_ru/n68 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1475  (\cu_ru/n69 [3], \cu_ru/n63 [3], \cu_ru/n68 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1476  (\cu_ru/n69 [4], \cu_ru/n63 [4], \cu_ru/n68 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1477  (\cu_ru/n69 [5], \cu_ru/n65 [5], \cu_ru/n68 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1478  (\cu_ru/n69 [6], \cu_ru/n63 [6], \cu_ru/n68 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1479  (\cu_ru/n69 [7], \cu_ru/n63 [7], \cu_ru/n68 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u148  (\cu_ru/n113 [37], \cu_ru/n109 [37], \cu_ru/n112 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1480  (\cu_ru/n69 [8], \cu_ru/n65 [8], \cu_ru/n68 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1481  (\cu_ru/n69 [9], \cu_ru/n63 [9], \cu_ru/n68 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1482  (\cu_ru/n69 [10], \cu_ru/n63 [10], \cu_ru/n68 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1483  (\cu_ru/n69 [11], \cu_ru/n63 [11], \cu_ru/n68 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1484  (\cu_ru/n69 [12], \cu_ru/n63 [12], \cu_ru/n68 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1485  (\cu_ru/n69 [13], \cu_ru/n63 [13], \cu_ru/n68 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1486  (\cu_ru/n69 [14], \cu_ru/n63 [14], \cu_ru/n68 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1487  (\cu_ru/n69 [15], \cu_ru/n63 [15], \cu_ru/n68 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1488  (\cu_ru/n69 [16], \cu_ru/n63 [16], \cu_ru/n68 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1489  (\cu_ru/n69 [17], \cu_ru/n63 [17], \cu_ru/n68 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u149  (\cu_ru/n113 [38], \cu_ru/n109 [38], \cu_ru/n112 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1490  (\cu_ru/n69 [18], \cu_ru/n65 [18], \cu_ru/n68 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1491  (\cu_ru/n69 [19], \cu_ru/n65 [19], \cu_ru/n68 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1492  (\cu_ru/n69 [20], \cu_ru/n63 [20], \cu_ru/n68 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1493  (\cu_ru/n69 [21], \cu_ru/n63 [21], \cu_ru/n68 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1494  (\cu_ru/n69 [22], \cu_ru/n63 [22], \cu_ru/n68 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1495  (\cu_ru/n69 [23], \cu_ru/n63 [23], \cu_ru/n68 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1496  (\cu_ru/n69 [24], \cu_ru/n63 [24], \cu_ru/n68 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1497  (\cu_ru/n69 [25], \cu_ru/n63 [25], \cu_ru/n68 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1498  (\cu_ru/n69 [26], \cu_ru/n63 [26], \cu_ru/n68 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1499  (\cu_ru/n69 [27], \cu_ru/n63 [27], \cu_ru/n68 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  and \cu_ru/u15  (\cu_ru/mrw_mtvec_sel , wb_valid, \cu_ru/n13 );  // ../../RTL/CPU/CU&RU/cu_ru.v(283)
  or \cu_ru/u150  (\cu_ru/n113 [39], \cu_ru/n109 [39], \cu_ru/n112 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1500  (\cu_ru/n69 [28], \cu_ru/n63 [28], \cu_ru/n68 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1501  (\cu_ru/n69 [29], \cu_ru/n63 [29], \cu_ru/n68 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1502  (\cu_ru/n69 [30], \cu_ru/n63 [30], \cu_ru/n68 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1503  (\cu_ru/n69 [31], \cu_ru/n63 [31], \cu_ru/n68 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1504  (\cu_ru/n69 [32], \cu_ru/n65 [32], \cu_ru/n68 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1505  (\cu_ru/n69 [33], \cu_ru/n65 [33], \cu_ru/n68 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1506  (\cu_ru/n69 [34], \cu_ru/n63 [34], \cu_ru/n68 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1507  (\cu_ru/n69 [35], \cu_ru/n63 [35], \cu_ru/n68 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1508  (\cu_ru/n69 [36], \cu_ru/n63 [36], \cu_ru/n68 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1509  (\cu_ru/n69 [37], \cu_ru/n63 [37], \cu_ru/n68 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u151  (\cu_ru/n113 [40], \cu_ru/n109 [40], \cu_ru/n112 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1510  (\cu_ru/n69 [38], \cu_ru/n63 [38], \cu_ru/n68 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1511  (\cu_ru/n69 [39], \cu_ru/n63 [39], \cu_ru/n68 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1512  (\cu_ru/n69 [40], \cu_ru/n63 [40], \cu_ru/n68 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1513  (\cu_ru/n69 [41], \cu_ru/n63 [41], \cu_ru/n68 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1514  (\cu_ru/n69 [42], \cu_ru/n63 [42], \cu_ru/n68 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1515  (\cu_ru/n69 [43], \cu_ru/n63 [43], \cu_ru/n68 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1516  (\cu_ru/n69 [44], \cu_ru/n63 [44], \cu_ru/n68 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1517  (\cu_ru/n69 [45], \cu_ru/n63 [45], \cu_ru/n68 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1518  (\cu_ru/n69 [46], \cu_ru/n63 [46], \cu_ru/n68 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1519  (\cu_ru/n69 [47], \cu_ru/n63 [47], \cu_ru/n68 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u152  (\cu_ru/n113 [41], \cu_ru/n109 [41], \cu_ru/n112 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1520  (\cu_ru/n69 [48], \cu_ru/n63 [48], \cu_ru/n68 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1521  (\cu_ru/n69 [49], \cu_ru/n63 [49], \cu_ru/n68 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1522  (\cu_ru/n69 [50], \cu_ru/n63 [50], \cu_ru/n68 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1523  (\cu_ru/n69 [51], \cu_ru/n63 [51], \cu_ru/n68 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1524  (\cu_ru/n69 [52], \cu_ru/n63 [52], \cu_ru/n68 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1525  (\cu_ru/n69 [53], \cu_ru/n63 [53], \cu_ru/n68 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1526  (\cu_ru/n69 [54], \cu_ru/n63 [54], \cu_ru/n68 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1527  (\cu_ru/n69 [55], \cu_ru/n63 [55], \cu_ru/n68 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1528  (\cu_ru/n69 [56], \cu_ru/n63 [56], \cu_ru/n68 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1529  (\cu_ru/n69 [57], \cu_ru/n63 [57], \cu_ru/n68 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u153  (\cu_ru/n113 [42], \cu_ru/n109 [42], \cu_ru/n112 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1530  (\cu_ru/n69 [58], \cu_ru/n63 [58], \cu_ru/n68 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1531  (\cu_ru/n69 [59], \cu_ru/n63 [59], \cu_ru/n68 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1532  (\cu_ru/n69 [60], \cu_ru/n63 [60], \cu_ru/n68 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1533  (\cu_ru/n69 [61], \cu_ru/n63 [61], \cu_ru/n68 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1534  (\cu_ru/n69 [62], \cu_ru/n63 [62], \cu_ru/n68 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1535  (\cu_ru/n69 [63], \cu_ru/n63 [63], \cu_ru/n68 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1536  (\cu_ru/n65 [1], \cu_ru/n63 [1], \cu_ru/n64 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  or \cu_ru/u154  (\cu_ru/n113 [43], \cu_ru/n109 [43], \cu_ru/n112 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u1540  (\cu_ru/n65 [5], \cu_ru/n63 [5], \cu_ru/n64 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  or \cu_ru/u1543  (\cu_ru/n65 [8], \cu_ru/n63 [8], \cu_ru/n64 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  AL_MUX \cu_ru/u155  (
    .i0(1'b0),
    .i1(\cu_ru/n51 ),
    .sel(wb_gpr_write),
    .o(\cu_ru/n53 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(371)
  or \cu_ru/u1553  (\cu_ru/n65 [18], \cu_ru/n63 [18], \cu_ru/n64 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  or \cu_ru/u1554  (\cu_ru/n65 [19], \cu_ru/n63 [19], \cu_ru/n64 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  or \cu_ru/u1567  (\cu_ru/n65 [32], \cu_ru/n63 [32], \cu_ru/n64 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  or \cu_ru/u1568  (\cu_ru/n65 [33], \cu_ru/n63 [33], \cu_ru/n64 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(676)
  or \cu_ru/u158  (\cu_ru/n56 , \cu_ru/trap_target_m , \cu_ru/trap_target_s );  // ../../RTL/CPU/CU&RU/cu_ru.v(667)
  or \cu_ru/u159  (csr_data[0], \cu_ru/n115 [0], \cu_ru/n116 );  // ../../RTL/CPU/CU&RU/cu_ru.v(706)
  or \cu_ru/u1599  (\cu_ru/n63 [1], \cu_ru/n61 [1], \cu_ru/n62 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  and \cu_ru/u16  (\cu_ru/mrw_mscratch_sel , wb_valid, \cu_ru/n14 );  // ../../RTL/CPU/CU&RU/cu_ru.v(285)
  or \cu_ru/u160  (pip_flush, \cu_ru/n56 , pc_jmp);  // ../../RTL/CPU/CU&RU/cu_ru.v(668)
  or \cu_ru/u1600  (\cu_ru/n63 [2], \cu_ru/n61 [2], \cu_ru/n62 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1601  (\cu_ru/n63 [3], \cu_ru/n61 [3], \cu_ru/n62 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1602  (\cu_ru/n63 [4], \cu_ru/n61 [4], \cu_ru/n62 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1603  (\cu_ru/n63 [5], \cu_ru/n61 [5], \cu_ru/n62 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1604  (\cu_ru/n63 [6], \cu_ru/n61 [6], \cu_ru/n62 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1605  (\cu_ru/n63 [7], \cu_ru/n61 [7], \cu_ru/n62 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1606  (\cu_ru/n63 [8], \cu_ru/n61 [8], \cu_ru/n62 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1607  (\cu_ru/n63 [9], \cu_ru/n61 [9], \cu_ru/n62 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1608  (\cu_ru/n63 [10], \cu_ru/n61 [10], \cu_ru/n62 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1609  (\cu_ru/n63 [11], \cu_ru/n61 [11], \cu_ru/n62 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1610  (\cu_ru/n63 [12], \cu_ru/n61 [12], \cu_ru/n62 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1611  (\cu_ru/n63 [13], \cu_ru/n61 [13], \cu_ru/n62 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1612  (\cu_ru/n63 [14], \cu_ru/n61 [14], \cu_ru/n62 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1613  (\cu_ru/n63 [15], \cu_ru/n61 [15], \cu_ru/n62 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1614  (\cu_ru/n63 [16], \cu_ru/n61 [16], \cu_ru/n62 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1615  (\cu_ru/n63 [17], \cu_ru/n61 [17], \cu_ru/n62 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1616  (\cu_ru/n63 [18], \cu_ru/n61 [18], \cu_ru/n62 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1617  (\cu_ru/n63 [19], \cu_ru/n61 [19], \cu_ru/n62 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1618  (\cu_ru/n63 [20], \cu_ru/n61 [20], \cu_ru/n62 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1619  (\cu_ru/n63 [21], \cu_ru/n61 [21], \cu_ru/n62 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u162  (\cu_ru/n61 [0], \cu_ru/n59 [0], \cu_ru/n60 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1620  (\cu_ru/n63 [22], \cu_ru/n61 [22], \cu_ru/n62 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1621  (\cu_ru/n63 [23], \cu_ru/n61 [23], \cu_ru/n62 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1622  (\cu_ru/n63 [24], \cu_ru/n61 [24], \cu_ru/n62 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1623  (\cu_ru/n63 [25], \cu_ru/n61 [25], \cu_ru/n62 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1624  (\cu_ru/n63 [26], \cu_ru/n61 [26], \cu_ru/n62 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1625  (\cu_ru/n63 [27], \cu_ru/n61 [27], \cu_ru/n62 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1626  (\cu_ru/n63 [28], \cu_ru/n61 [28], \cu_ru/n62 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1627  (\cu_ru/n63 [29], \cu_ru/n61 [29], \cu_ru/n62 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1628  (\cu_ru/n63 [30], \cu_ru/n61 [30], \cu_ru/n62 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1629  (\cu_ru/n63 [31], \cu_ru/n61 [31], \cu_ru/n62 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u163  (\cu_ru/n63 [0], \cu_ru/n61 [0], \cu_ru/n62 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1630  (\cu_ru/n63 [32], \cu_ru/n61 [32], \cu_ru/n62 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1631  (\cu_ru/n63 [33], \cu_ru/n61 [33], \cu_ru/n62 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1632  (\cu_ru/n63 [34], \cu_ru/n61 [34], \cu_ru/n62 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1633  (\cu_ru/n63 [35], \cu_ru/n61 [35], \cu_ru/n62 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1634  (\cu_ru/n63 [36], \cu_ru/n61 [36], \cu_ru/n62 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1635  (\cu_ru/n63 [37], \cu_ru/n61 [37], \cu_ru/n62 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1636  (\cu_ru/n63 [38], \cu_ru/n61 [38], \cu_ru/n62 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1637  (\cu_ru/n63 [39], \cu_ru/n61 [39], \cu_ru/n62 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1638  (\cu_ru/n63 [40], \cu_ru/n61 [40], \cu_ru/n62 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1639  (\cu_ru/n63 [41], \cu_ru/n61 [41], \cu_ru/n62 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  AL_MUX \cu_ru/u164  (
    .i0(1'b0),
    .i1(\cu_ru/mstatus [1]),
    .sel(\cu_ru/read_sie_sel ),
    .o(\cu_ru/n66 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(677)
  or \cu_ru/u1640  (\cu_ru/n63 [42], \cu_ru/n61 [42], \cu_ru/n62 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1641  (\cu_ru/n63 [43], \cu_ru/n61 [43], \cu_ru/n62 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1642  (\cu_ru/n63 [44], \cu_ru/n61 [44], \cu_ru/n62 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1643  (\cu_ru/n63 [45], \cu_ru/n61 [45], \cu_ru/n62 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1644  (\cu_ru/n63 [46], \cu_ru/n61 [46], \cu_ru/n62 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1645  (\cu_ru/n63 [47], \cu_ru/n61 [47], \cu_ru/n62 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1646  (\cu_ru/n63 [48], \cu_ru/n61 [48], \cu_ru/n62 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1647  (\cu_ru/n63 [49], \cu_ru/n61 [49], \cu_ru/n62 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1648  (\cu_ru/n63 [50], \cu_ru/n61 [50], \cu_ru/n62 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1649  (\cu_ru/n63 [51], \cu_ru/n61 [51], \cu_ru/n62 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1650  (\cu_ru/n63 [52], \cu_ru/n61 [52], \cu_ru/n62 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1651  (\cu_ru/n63 [53], \cu_ru/n61 [53], \cu_ru/n62 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1652  (\cu_ru/n63 [54], \cu_ru/n61 [54], \cu_ru/n62 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1653  (\cu_ru/n63 [55], \cu_ru/n61 [55], \cu_ru/n62 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1654  (\cu_ru/n63 [56], \cu_ru/n61 [56], \cu_ru/n62 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1655  (\cu_ru/n63 [57], \cu_ru/n61 [57], \cu_ru/n62 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1656  (\cu_ru/n63 [58], \cu_ru/n61 [58], \cu_ru/n62 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1657  (\cu_ru/n63 [59], \cu_ru/n61 [59], \cu_ru/n62 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1658  (\cu_ru/n63 [60], \cu_ru/n61 [60], \cu_ru/n62 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1659  (\cu_ru/n63 [61], \cu_ru/n61 [61], \cu_ru/n62 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u166  (\cu_ru/n67 [0], \cu_ru/n63 [0], \cu_ru/n66 );  // ../../RTL/CPU/CU&RU/cu_ru.v(677)
  or \cu_ru/u1660  (\cu_ru/n63 [62], \cu_ru/n61 [62], \cu_ru/n62 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1661  (\cu_ru/n63 [63], \cu_ru/n61 [63], \cu_ru/n62 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(674)
  or \cu_ru/u1662  (\cu_ru/n61 [1], \cu_ru/n59 [1], \cu_ru/n60 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1663  (\cu_ru/n61 [2], \cu_ru/n59 [2], \cu_ru/n60 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1664  (\cu_ru/n61 [3], \cu_ru/n59 [3], \cu_ru/n60 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1665  (\cu_ru/n61 [4], \cu_ru/n59 [4], \cu_ru/n60 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1666  (\cu_ru/n61 [5], \cu_ru/n59 [5], \cu_ru/n60 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1667  (\cu_ru/n61 [6], \cu_ru/n59 [6], \cu_ru/n60 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1668  (\cu_ru/n61 [7], \cu_ru/n59 [7], \cu_ru/n60 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1669  (\cu_ru/n61 [8], \cu_ru/n59 [8], \cu_ru/n60 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u167  (\cu_ru/n69 [0], \cu_ru/n67 [0], \cu_ru/n68 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(678)
  or \cu_ru/u1670  (\cu_ru/n61 [9], \cu_ru/n59 [9], \cu_ru/n60 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1671  (\cu_ru/n61 [10], \cu_ru/n59 [10], \cu_ru/n60 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1672  (\cu_ru/n61 [11], \cu_ru/n59 [11], \cu_ru/n60 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1673  (\cu_ru/n61 [12], \cu_ru/n59 [12], \cu_ru/n60 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1674  (\cu_ru/n61 [13], \cu_ru/n59 [13], \cu_ru/n60 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1675  (\cu_ru/n61 [14], \cu_ru/n59 [14], \cu_ru/n60 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1676  (\cu_ru/n61 [15], \cu_ru/n59 [15], \cu_ru/n60 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1677  (\cu_ru/n61 [16], \cu_ru/n59 [16], \cu_ru/n60 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1678  (\cu_ru/n61 [17], \cu_ru/n59 [17], \cu_ru/n60 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1679  (\cu_ru/n61 [18], \cu_ru/n59 [18], \cu_ru/n60 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u168  (\cu_ru/n71 [0], \cu_ru/n69 [0], \cu_ru/n70 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(680)
  or \cu_ru/u1680  (\cu_ru/n61 [19], \cu_ru/n59 [19], \cu_ru/n60 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1681  (\cu_ru/n61 [20], \cu_ru/n59 [20], \cu_ru/n60 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1682  (\cu_ru/n61 [21], \cu_ru/n59 [21], \cu_ru/n60 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1683  (\cu_ru/n61 [22], \cu_ru/n59 [22], \cu_ru/n60 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1684  (\cu_ru/n61 [23], \cu_ru/n59 [23], \cu_ru/n60 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1685  (\cu_ru/n61 [24], \cu_ru/n59 [24], \cu_ru/n60 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1686  (\cu_ru/n61 [25], \cu_ru/n59 [25], \cu_ru/n60 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1687  (\cu_ru/n61 [26], \cu_ru/n59 [26], \cu_ru/n60 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1688  (\cu_ru/n61 [27], \cu_ru/n59 [27], \cu_ru/n60 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1689  (\cu_ru/n61 [28], \cu_ru/n59 [28], \cu_ru/n60 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u169  (\cu_ru/n73 [0], \cu_ru/n71 [0], \cu_ru/n72 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(681)
  or \cu_ru/u1690  (\cu_ru/n61 [29], \cu_ru/n59 [29], \cu_ru/n60 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1691  (\cu_ru/n61 [30], \cu_ru/n59 [30], \cu_ru/n60 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1692  (\cu_ru/n61 [31], \cu_ru/n59 [31], \cu_ru/n60 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1693  (\cu_ru/n61 [32], \cu_ru/n59 [32], \cu_ru/n60 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1694  (\cu_ru/n61 [33], \cu_ru/n59 [33], \cu_ru/n60 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1695  (\cu_ru/n61 [34], \cu_ru/n59 [34], \cu_ru/n60 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1696  (\cu_ru/n61 [35], \cu_ru/n59 [35], \cu_ru/n60 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1697  (\cu_ru/n61 [36], \cu_ru/n59 [36], \cu_ru/n60 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1698  (\cu_ru/n61 [37], \cu_ru/n59 [37], \cu_ru/n60 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1699  (\cu_ru/n61 [38], \cu_ru/n59 [38], \cu_ru/n60 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  and \cu_ru/u17  (\cu_ru/mrw_mepc_sel , wb_valid, \cu_ru/n15 );  // ../../RTL/CPU/CU&RU/cu_ru.v(286)
  or \cu_ru/u170  (\cu_ru/n75 [0], \cu_ru/n73 [0], \cu_ru/n74 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(682)
  or \cu_ru/u1700  (\cu_ru/n61 [39], \cu_ru/n59 [39], \cu_ru/n60 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1701  (\cu_ru/n61 [40], \cu_ru/n59 [40], \cu_ru/n60 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1702  (\cu_ru/n61 [41], \cu_ru/n59 [41], \cu_ru/n60 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1703  (\cu_ru/n61 [42], \cu_ru/n59 [42], \cu_ru/n60 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1704  (\cu_ru/n61 [43], \cu_ru/n59 [43], \cu_ru/n60 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1705  (\cu_ru/n61 [44], \cu_ru/n59 [44], \cu_ru/n60 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1706  (\cu_ru/n61 [45], \cu_ru/n59 [45], \cu_ru/n60 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1707  (\cu_ru/n61 [46], \cu_ru/n59 [46], \cu_ru/n60 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1708  (\cu_ru/n61 [47], \cu_ru/n59 [47], \cu_ru/n60 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1709  (\cu_ru/n61 [48], \cu_ru/n59 [48], \cu_ru/n60 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u171  (\cu_ru/n77 [0], \cu_ru/n75 [0], \cu_ru/n76 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(683)
  or \cu_ru/u1710  (\cu_ru/n61 [49], \cu_ru/n59 [49], \cu_ru/n60 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1711  (\cu_ru/n61 [50], \cu_ru/n59 [50], \cu_ru/n60 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1712  (\cu_ru/n61 [51], \cu_ru/n59 [51], \cu_ru/n60 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1713  (\cu_ru/n61 [52], \cu_ru/n59 [52], \cu_ru/n60 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1714  (\cu_ru/n61 [53], \cu_ru/n59 [53], \cu_ru/n60 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1715  (\cu_ru/n61 [54], \cu_ru/n59 [54], \cu_ru/n60 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1716  (\cu_ru/n61 [55], \cu_ru/n59 [55], \cu_ru/n60 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1717  (\cu_ru/n61 [56], \cu_ru/n59 [56], \cu_ru/n60 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1718  (\cu_ru/n61 [57], \cu_ru/n59 [57], \cu_ru/n60 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1719  (\cu_ru/n61 [58], \cu_ru/n59 [58], \cu_ru/n60 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1720  (\cu_ru/n61 [59], \cu_ru/n59 [59], \cu_ru/n60 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1721  (\cu_ru/n61 [60], \cu_ru/n59 [60], \cu_ru/n60 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1722  (\cu_ru/n61 [61], \cu_ru/n59 [61], \cu_ru/n60 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1723  (\cu_ru/n61 [62], \cu_ru/n59 [62], \cu_ru/n60 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u1724  (\cu_ru/n61 [63], \cu_ru/n59 [63], \cu_ru/n60 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(673)
  or \cu_ru/u173  (\cu_ru/n81 [0], \cu_ru/n77 [0], \cu_ru/n80 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(685)
  and \cu_ru/u18  (\cu_ru/mrw_mcause_sel , wb_valid, \cu_ru/n16 );  // ../../RTL/CPU/CU&RU/cu_ru.v(287)
  or \cu_ru/u180  (\cu_ru/n95 [0], \cu_ru/n81 [0], \cu_ru/n94 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  AL_MUX \cu_ru/u181  (
    .i0(1'b0),
    .i1(\cu_ru/mie ),
    .sel(\cu_ru/read_mie_sel ),
    .o(\cu_ru/n98 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(694)
  or \cu_ru/u183  (\cu_ru/n99 [0], \cu_ru/n95 [0], \cu_ru/n98 );  // ../../RTL/CPU/CU&RU/cu_ru.v(694)
  or \cu_ru/u184  (\cu_ru/n101 [0], \cu_ru/n99 [0], \cu_ru/n100 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u185  (\cu_ru/n103 [0], \cu_ru/n101 [0], \cu_ru/n102 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u186  (\cu_ru/n105 [0], \cu_ru/n103 [0], \cu_ru/n104 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u187  (\cu_ru/n107 [0], \cu_ru/n105 [0], \cu_ru/n106 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u188  (\cu_ru/n109 [0], \cu_ru/n107 [0], \cu_ru/n108 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  and \cu_ru/u19  (\cu_ru/mrw_mtval_sel , wb_valid, \cu_ru/n17 );  // ../../RTL/CPU/CU&RU/cu_ru.v(288)
  or \cu_ru/u190  (\cu_ru/n113 [0], \cu_ru/n109 [0], \cu_ru/n112 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  AL_MUX \cu_ru/u191  (
    .i0(1'b0),
    .i1(\cu_ru/mcountinhibit ),
    .sel(\cu_ru/read_mcounterinhibit_sel ),
    .o(\cu_ru/n116 ));  // ../../RTL/CPU/CU&RU/cu_ru.v(706)
  or \cu_ru/u192  (\cu_ru/n115 [0], \cu_ru/n113 [0], \cu_ru/n114 [0]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u193  (\cu_ru/n113 [44], \cu_ru/n109 [44], \cu_ru/n112 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u194  (\cu_ru/n113 [45], \cu_ru/n109 [45], \cu_ru/n112 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u195  (\cu_ru/n113 [46], \cu_ru/n109 [46], \cu_ru/n112 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u196  (\cu_ru/n113 [47], \cu_ru/n109 [47], \cu_ru/n112 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u197  (\cu_ru/n113 [48], \cu_ru/n109 [48], \cu_ru/n112 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u198  (\cu_ru/n113 [49], \cu_ru/n109 [49], \cu_ru/n112 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u199  (\cu_ru/n113 [50], \cu_ru/n109 [50], \cu_ru/n112 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  and \cu_ru/u2  (\cu_ru/srw_sstatus_sel , wb_valid, \cu_ru/n0 );  // ../../RTL/CPU/CU&RU/cu_ru.v(264)
  and \cu_ru/u20  (\cu_ru/mrw_mip_sel , wb_valid, \cu_ru/n18 );  // ../../RTL/CPU/CU&RU/cu_ru.v(289)
  or \cu_ru/u200  (\cu_ru/n113 [51], \cu_ru/n109 [51], \cu_ru/n112 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u201  (\cu_ru/n113 [52], \cu_ru/n109 [52], \cu_ru/n112 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u202  (\cu_ru/n113 [53], \cu_ru/n109 [53], \cu_ru/n112 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u203  (\cu_ru/n113 [54], \cu_ru/n109 [54], \cu_ru/n112 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u204  (\cu_ru/n113 [55], \cu_ru/n109 [55], \cu_ru/n112 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u205  (\cu_ru/n113 [56], \cu_ru/n109 [56], \cu_ru/n112 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u206  (\cu_ru/n113 [57], \cu_ru/n109 [57], \cu_ru/n112 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u207  (\cu_ru/n113 [58], \cu_ru/n109 [58], \cu_ru/n112 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u208  (\cu_ru/n113 [59], \cu_ru/n109 [59], \cu_ru/n112 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u209  (\cu_ru/n113 [60], \cu_ru/n109 [60], \cu_ru/n112 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  and \cu_ru/u21  (\cu_ru/mrw_mcycle_sel , wb_valid, \cu_ru/n19 );  // ../../RTL/CPU/CU&RU/cu_ru.v(293)
  or \cu_ru/u210  (\cu_ru/n113 [61], \cu_ru/n109 [61], \cu_ru/n112 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u211  (\cu_ru/n113 [62], \cu_ru/n109 [62], \cu_ru/n112 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u212  (\cu_ru/n113 [63], \cu_ru/n109 [63], \cu_ru/n112 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(703)
  or \cu_ru/u213  (\cu_ru/n111 [1], \cu_ru/n109 [1], \cu_ru/n110 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  or \cu_ru/u215  (\cu_ru/n111 [3], \cu_ru/n109 [3], \cu_ru/n110 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  or \cu_ru/u217  (\cu_ru/n111 [5], \cu_ru/n109 [5], \cu_ru/n110 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  or \cu_ru/u219  (\cu_ru/n111 [7], \cu_ru/n109 [7], \cu_ru/n110 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  and \cu_ru/u22  (\cu_ru/mrw_mcounterinhibit_sel , wb_valid, \cu_ru/n20 );  // ../../RTL/CPU/CU&RU/cu_ru.v(297)
  or \cu_ru/u221  (\cu_ru/n111 [9], \cu_ru/n109 [9], \cu_ru/n110 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  or \cu_ru/u223  (\cu_ru/n111 [11], \cu_ru/n109 [11], \cu_ru/n110 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(701)
  or \cu_ru/u25  (\cu_ru/n23 , \cu_ru/m_s_tval/n1 , wb_ill_ins);  // ../../RTL/CPU/CU&RU/cu_ru.v(341)
  or \cu_ru/u26  (\cu_ru/n24 , \cu_ru/n23 , wb_ld_acc_fault);  // ../../RTL/CPU/CU&RU/cu_ru.v(341)
  or \cu_ru/u27  (\cu_ru/n25 , \cu_ru/n24 , wb_ld_page_fault);  // ../../RTL/CPU/CU&RU/cu_ru.v(341)
  or \cu_ru/u276  (\cu_ru/n109 [1], \cu_ru/n107 [1], \cu_ru/n108 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u277  (\cu_ru/n109 [2], \cu_ru/n107 [2], \cu_ru/n108 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u278  (\cu_ru/n109 [3], \cu_ru/n107 [3], \cu_ru/n108 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u279  (\cu_ru/n109 [4], \cu_ru/n107 [4], \cu_ru/n108 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u28  (\cu_ru/n26 , \cu_ru/n25 , wb_st_acc_fault);  // ../../RTL/CPU/CU&RU/cu_ru.v(341)
  or \cu_ru/u280  (\cu_ru/n109 [5], \cu_ru/n107 [5], \cu_ru/n108 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u281  (\cu_ru/n109 [6], \cu_ru/n107 [6], \cu_ru/n108 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u282  (\cu_ru/n109 [7], \cu_ru/n107 [7], \cu_ru/n108 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u283  (\cu_ru/n109 [8], \cu_ru/n107 [8], \cu_ru/n108 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u284  (\cu_ru/n109 [9], \cu_ru/n107 [9], \cu_ru/n108 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u285  (\cu_ru/n109 [10], \cu_ru/n107 [10], \cu_ru/n108 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u286  (\cu_ru/n109 [11], \cu_ru/n107 [11], \cu_ru/n108 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u287  (\cu_ru/n109 [12], \cu_ru/n107 [12], \cu_ru/n108 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u288  (\cu_ru/n109 [13], \cu_ru/n107 [13], \cu_ru/n108 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u289  (\cu_ru/n109 [14], \cu_ru/n107 [14], \cu_ru/n108 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u29  (\cu_ru/n27 , \cu_ru/n26 , wb_st_page_fault);  // ../../RTL/CPU/CU&RU/cu_ru.v(341)
  or \cu_ru/u290  (\cu_ru/n109 [15], \cu_ru/n107 [15], \cu_ru/n108 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u291  (\cu_ru/n109 [16], \cu_ru/n107 [16], \cu_ru/n108 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u292  (\cu_ru/n109 [17], \cu_ru/n107 [17], \cu_ru/n108 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u293  (\cu_ru/n109 [18], \cu_ru/n107 [18], \cu_ru/n108 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u294  (\cu_ru/n109 [19], \cu_ru/n107 [19], \cu_ru/n108 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u295  (\cu_ru/n109 [20], \cu_ru/n107 [20], \cu_ru/n108 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u296  (\cu_ru/n109 [21], \cu_ru/n107 [21], \cu_ru/n108 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u297  (\cu_ru/n109 [22], \cu_ru/n107 [22], \cu_ru/n108 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u298  (\cu_ru/n109 [23], \cu_ru/n107 [23], \cu_ru/n108 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u299  (\cu_ru/n109 [24], \cu_ru/n107 [24], \cu_ru/n108 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  and \cu_ru/u3  (\cu_ru/srw_sie_sel , wb_valid, \cu_ru/n1 );  // ../../RTL/CPU/CU&RU/cu_ru.v(265)
  or \cu_ru/u30  (\cu_ru/n28 , \cu_ru/n27 , wb_ld_addr_mis);  // ../../RTL/CPU/CU&RU/cu_ru.v(341)
  or \cu_ru/u300  (\cu_ru/n109 [25], \cu_ru/n107 [25], \cu_ru/n108 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u301  (\cu_ru/n109 [26], \cu_ru/n107 [26], \cu_ru/n108 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u302  (\cu_ru/n109 [27], \cu_ru/n107 [27], \cu_ru/n108 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u303  (\cu_ru/n109 [28], \cu_ru/n107 [28], \cu_ru/n108 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u304  (\cu_ru/n109 [29], \cu_ru/n107 [29], \cu_ru/n108 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u305  (\cu_ru/n109 [30], \cu_ru/n107 [30], \cu_ru/n108 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u306  (\cu_ru/n109 [31], \cu_ru/n107 [31], \cu_ru/n108 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u307  (\cu_ru/n109 [32], \cu_ru/n107 [32], \cu_ru/n108 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u308  (\cu_ru/n109 [33], \cu_ru/n107 [33], \cu_ru/n108 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u309  (\cu_ru/n109 [34], \cu_ru/n107 [34], \cu_ru/n108 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u31  (\cu_ru/n29 , \cu_ru/n28 , wb_st_addr_mis);  // ../../RTL/CPU/CU&RU/cu_ru.v(341)
  or \cu_ru/u310  (\cu_ru/n109 [35], \cu_ru/n107 [35], \cu_ru/n108 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u311  (\cu_ru/n109 [36], \cu_ru/n107 [36], \cu_ru/n108 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u312  (\cu_ru/n109 [37], \cu_ru/n107 [37], \cu_ru/n108 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u313  (\cu_ru/n109 [38], \cu_ru/n107 [38], \cu_ru/n108 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u314  (\cu_ru/n109 [39], \cu_ru/n107 [39], \cu_ru/n108 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u315  (\cu_ru/n109 [40], \cu_ru/n107 [40], \cu_ru/n108 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u316  (\cu_ru/n109 [41], \cu_ru/n107 [41], \cu_ru/n108 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u317  (\cu_ru/n109 [42], \cu_ru/n107 [42], \cu_ru/n108 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u318  (\cu_ru/n109 [43], \cu_ru/n107 [43], \cu_ru/n108 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u319  (\cu_ru/n109 [44], \cu_ru/n107 [44], \cu_ru/n108 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u32  (\cu_ru/n30 , \cu_ru/n29 , wb_ecall);  // ../../RTL/CPU/CU&RU/cu_ru.v(341)
  or \cu_ru/u320  (\cu_ru/n109 [45], \cu_ru/n107 [45], \cu_ru/n108 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u321  (\cu_ru/n109 [46], \cu_ru/n107 [46], \cu_ru/n108 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u322  (\cu_ru/n109 [47], \cu_ru/n107 [47], \cu_ru/n108 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u323  (\cu_ru/n109 [48], \cu_ru/n107 [48], \cu_ru/n108 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u324  (\cu_ru/n109 [49], \cu_ru/n107 [49], \cu_ru/n108 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u325  (\cu_ru/n109 [50], \cu_ru/n107 [50], \cu_ru/n108 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u326  (\cu_ru/n109 [51], \cu_ru/n107 [51], \cu_ru/n108 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u327  (\cu_ru/n109 [52], \cu_ru/n107 [52], \cu_ru/n108 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u328  (\cu_ru/n109 [53], \cu_ru/n107 [53], \cu_ru/n108 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u329  (\cu_ru/n109 [54], \cu_ru/n107 [54], \cu_ru/n108 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u33  (\cu_ru/n31 , \cu_ru/n30 , wb_ebreak);  // ../../RTL/CPU/CU&RU/cu_ru.v(341)
  or \cu_ru/u330  (\cu_ru/n109 [55], \cu_ru/n107 [55], \cu_ru/n108 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u331  (\cu_ru/n109 [56], \cu_ru/n107 [56], \cu_ru/n108 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u332  (\cu_ru/n109 [57], \cu_ru/n107 [57], \cu_ru/n108 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u333  (\cu_ru/n109 [58], \cu_ru/n107 [58], \cu_ru/n108 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u334  (\cu_ru/n109 [59], \cu_ru/n107 [59], \cu_ru/n108 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u335  (\cu_ru/n109 [60], \cu_ru/n107 [60], \cu_ru/n108 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u336  (\cu_ru/n109 [61], \cu_ru/n107 [61], \cu_ru/n108 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u337  (\cu_ru/n109 [62], \cu_ru/n107 [62], \cu_ru/n108 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u338  (\cu_ru/n109 [63], \cu_ru/n107 [63], \cu_ru/n108 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(700)
  or \cu_ru/u339  (\cu_ru/n107 [1], \cu_ru/n105 [1], \cu_ru/n106 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  and \cu_ru/u34  (\cu_ru/exception , wb_valid, \cu_ru/n31 );  // ../../RTL/CPU/CU&RU/cu_ru.v(341)
  or \cu_ru/u340  (\cu_ru/n107 [2], \cu_ru/n105 [2], \cu_ru/n106 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u341  (\cu_ru/n107 [3], \cu_ru/n105 [3], \cu_ru/n106 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u342  (\cu_ru/n107 [4], \cu_ru/n105 [4], \cu_ru/n106 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u343  (\cu_ru/n107 [5], \cu_ru/n105 [5], \cu_ru/n106 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u344  (\cu_ru/n107 [6], \cu_ru/n105 [6], \cu_ru/n106 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u345  (\cu_ru/n107 [7], \cu_ru/n105 [7], \cu_ru/n106 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u346  (\cu_ru/n107 [8], \cu_ru/n105 [8], \cu_ru/n106 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u347  (\cu_ru/n107 [9], \cu_ru/n105 [9], \cu_ru/n106 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u348  (\cu_ru/n107 [10], \cu_ru/n105 [10], \cu_ru/n106 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u349  (\cu_ru/n107 [11], \cu_ru/n105 [11], \cu_ru/n106 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u350  (\cu_ru/n107 [12], \cu_ru/n105 [12], \cu_ru/n106 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u351  (\cu_ru/n107 [13], \cu_ru/n105 [13], \cu_ru/n106 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u352  (\cu_ru/n107 [14], \cu_ru/n105 [14], \cu_ru/n106 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u353  (\cu_ru/n107 [15], \cu_ru/n105 [15], \cu_ru/n106 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u354  (\cu_ru/n107 [16], \cu_ru/n105 [16], \cu_ru/n106 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u355  (\cu_ru/n107 [17], \cu_ru/n105 [17], \cu_ru/n106 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u356  (\cu_ru/n107 [18], \cu_ru/n105 [18], \cu_ru/n106 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u357  (\cu_ru/n107 [19], \cu_ru/n105 [19], \cu_ru/n106 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u358  (\cu_ru/n107 [20], \cu_ru/n105 [20], \cu_ru/n106 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u359  (\cu_ru/n107 [21], \cu_ru/n105 [21], \cu_ru/n106 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  and \cu_ru/u36  (\cu_ru/n33 , \cu_ru/exception_neg , wb_valid);  // ../../RTL/CPU/CU&RU/cu_ru.v(344)
  or \cu_ru/u360  (\cu_ru/n107 [22], \cu_ru/n105 [22], \cu_ru/n106 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u361  (\cu_ru/n107 [23], \cu_ru/n105 [23], \cu_ru/n106 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u362  (\cu_ru/n107 [24], \cu_ru/n105 [24], \cu_ru/n106 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u363  (\cu_ru/n107 [25], \cu_ru/n105 [25], \cu_ru/n106 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u364  (\cu_ru/n107 [26], \cu_ru/n105 [26], \cu_ru/n106 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u365  (\cu_ru/n107 [27], \cu_ru/n105 [27], \cu_ru/n106 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u366  (\cu_ru/n107 [28], \cu_ru/n105 [28], \cu_ru/n106 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u367  (\cu_ru/n107 [29], \cu_ru/n105 [29], \cu_ru/n106 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u368  (\cu_ru/n107 [30], \cu_ru/n105 [30], \cu_ru/n106 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u369  (\cu_ru/n107 [31], \cu_ru/n105 [31], \cu_ru/n106 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  and \cu_ru/u37  (\cu_ru/n34 , \cu_ru/n33 , \cu_ru/int_target_m );  // ../../RTL/CPU/CU&RU/cu_ru.v(344)
  or \cu_ru/u370  (\cu_ru/n107 [32], \cu_ru/n105 [32], \cu_ru/n106 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u371  (\cu_ru/n107 [33], \cu_ru/n105 [33], \cu_ru/n106 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u372  (\cu_ru/n107 [34], \cu_ru/n105 [34], \cu_ru/n106 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u373  (\cu_ru/n107 [35], \cu_ru/n105 [35], \cu_ru/n106 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u374  (\cu_ru/n107 [36], \cu_ru/n105 [36], \cu_ru/n106 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u375  (\cu_ru/n107 [37], \cu_ru/n105 [37], \cu_ru/n106 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u376  (\cu_ru/n107 [38], \cu_ru/n105 [38], \cu_ru/n106 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u377  (\cu_ru/n107 [39], \cu_ru/n105 [39], \cu_ru/n106 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u378  (\cu_ru/n107 [40], \cu_ru/n105 [40], \cu_ru/n106 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u379  (\cu_ru/n107 [41], \cu_ru/n105 [41], \cu_ru/n106 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  and \cu_ru/u38  (\cu_ru/n35 , \cu_ru/n34 , int_req);  // ../../RTL/CPU/CU&RU/cu_ru.v(344)
  or \cu_ru/u380  (\cu_ru/n107 [42], \cu_ru/n105 [42], \cu_ru/n106 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u381  (\cu_ru/n107 [43], \cu_ru/n105 [43], \cu_ru/n106 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u382  (\cu_ru/n107 [44], \cu_ru/n105 [44], \cu_ru/n106 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u383  (\cu_ru/n107 [45], \cu_ru/n105 [45], \cu_ru/n106 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u384  (\cu_ru/n107 [46], \cu_ru/n105 [46], \cu_ru/n106 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u385  (\cu_ru/n107 [47], \cu_ru/n105 [47], \cu_ru/n106 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u386  (\cu_ru/n107 [48], \cu_ru/n105 [48], \cu_ru/n106 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u387  (\cu_ru/n107 [49], \cu_ru/n105 [49], \cu_ru/n106 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u388  (\cu_ru/n107 [50], \cu_ru/n105 [50], \cu_ru/n106 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u389  (\cu_ru/n107 [51], \cu_ru/n105 [51], \cu_ru/n106 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  and \cu_ru/u39  (\cu_ru/n36 , \cu_ru/n35 , wb_int_acc);  // ../../RTL/CPU/CU&RU/cu_ru.v(344)
  or \cu_ru/u390  (\cu_ru/n107 [52], \cu_ru/n105 [52], \cu_ru/n106 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u391  (\cu_ru/n107 [53], \cu_ru/n105 [53], \cu_ru/n106 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u392  (\cu_ru/n107 [54], \cu_ru/n105 [54], \cu_ru/n106 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u393  (\cu_ru/n107 [55], \cu_ru/n105 [55], \cu_ru/n106 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u394  (\cu_ru/n107 [56], \cu_ru/n105 [56], \cu_ru/n106 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u395  (\cu_ru/n107 [57], \cu_ru/n105 [57], \cu_ru/n106 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u396  (\cu_ru/n107 [58], \cu_ru/n105 [58], \cu_ru/n106 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u397  (\cu_ru/n107 [59], \cu_ru/n105 [59], \cu_ru/n106 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u398  (\cu_ru/n107 [60], \cu_ru/n105 [60], \cu_ru/n106 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u399  (\cu_ru/n107 [61], \cu_ru/n105 [61], \cu_ru/n106 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  and \cu_ru/u4  (\cu_ru/srw_stvec_sel , wb_valid, \cu_ru/n2 );  // ../../RTL/CPU/CU&RU/cu_ru.v(266)
  and \cu_ru/u40  (\cu_ru/n37 , wb_valid, \cu_ru/exc_target_m );  // ../../RTL/CPU/CU&RU/cu_ru.v(344)
  or \cu_ru/u400  (\cu_ru/n107 [62], \cu_ru/n105 [62], \cu_ru/n106 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u401  (\cu_ru/n107 [63], \cu_ru/n105 [63], \cu_ru/n106 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(699)
  or \cu_ru/u402  (\cu_ru/n105 [1], \cu_ru/n103 [1], \cu_ru/n104 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u403  (\cu_ru/n105 [2], \cu_ru/n103 [2], \cu_ru/n104 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u404  (\cu_ru/n105 [3], \cu_ru/n103 [3], \cu_ru/n104 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u405  (\cu_ru/n105 [4], \cu_ru/n103 [4], \cu_ru/n104 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u406  (\cu_ru/n105 [5], \cu_ru/n103 [5], \cu_ru/n104 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u407  (\cu_ru/n105 [6], \cu_ru/n103 [6], \cu_ru/n104 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u408  (\cu_ru/n105 [7], \cu_ru/n103 [7], \cu_ru/n104 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u409  (\cu_ru/n105 [8], \cu_ru/n103 [8], \cu_ru/n104 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u41  (\cu_ru/trap_target_m , \cu_ru/n36 , \cu_ru/n37 );  // ../../RTL/CPU/CU&RU/cu_ru.v(344)
  or \cu_ru/u410  (\cu_ru/n105 [9], \cu_ru/n103 [9], \cu_ru/n104 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u411  (\cu_ru/n105 [10], \cu_ru/n103 [10], \cu_ru/n104 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u412  (\cu_ru/n105 [11], \cu_ru/n103 [11], \cu_ru/n104 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u413  (\cu_ru/n105 [12], \cu_ru/n103 [12], \cu_ru/n104 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u414  (\cu_ru/n105 [13], \cu_ru/n103 [13], \cu_ru/n104 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u415  (\cu_ru/n105 [14], \cu_ru/n103 [14], \cu_ru/n104 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u416  (\cu_ru/n105 [15], \cu_ru/n103 [15], \cu_ru/n104 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u417  (\cu_ru/n105 [16], \cu_ru/n103 [16], \cu_ru/n104 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u418  (\cu_ru/n105 [17], \cu_ru/n103 [17], \cu_ru/n104 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u419  (\cu_ru/n105 [18], \cu_ru/n103 [18], \cu_ru/n104 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  and \cu_ru/u42  (\cu_ru/n38 , \cu_ru/n33 , \cu_ru/int_target_s );  // ../../RTL/CPU/CU&RU/cu_ru.v(345)
  or \cu_ru/u420  (\cu_ru/n105 [19], \cu_ru/n103 [19], \cu_ru/n104 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u421  (\cu_ru/n105 [20], \cu_ru/n103 [20], \cu_ru/n104 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u422  (\cu_ru/n105 [21], \cu_ru/n103 [21], \cu_ru/n104 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u423  (\cu_ru/n105 [22], \cu_ru/n103 [22], \cu_ru/n104 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u424  (\cu_ru/n105 [23], \cu_ru/n103 [23], \cu_ru/n104 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u425  (\cu_ru/n105 [24], \cu_ru/n103 [24], \cu_ru/n104 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u426  (\cu_ru/n105 [25], \cu_ru/n103 [25], \cu_ru/n104 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u427  (\cu_ru/n105 [26], \cu_ru/n103 [26], \cu_ru/n104 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u428  (\cu_ru/n105 [27], \cu_ru/n103 [27], \cu_ru/n104 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u429  (\cu_ru/n105 [28], \cu_ru/n103 [28], \cu_ru/n104 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  and \cu_ru/u43  (\cu_ru/n39 , \cu_ru/n38 , int_req);  // ../../RTL/CPU/CU&RU/cu_ru.v(345)
  or \cu_ru/u430  (\cu_ru/n105 [29], \cu_ru/n103 [29], \cu_ru/n104 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u431  (\cu_ru/n105 [30], \cu_ru/n103 [30], \cu_ru/n104 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u432  (\cu_ru/n105 [31], \cu_ru/n103 [31], \cu_ru/n104 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u433  (\cu_ru/n105 [32], \cu_ru/n103 [32], \cu_ru/n104 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u434  (\cu_ru/n105 [33], \cu_ru/n103 [33], \cu_ru/n104 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u435  (\cu_ru/n105 [34], \cu_ru/n103 [34], \cu_ru/n104 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u436  (\cu_ru/n105 [35], \cu_ru/n103 [35], \cu_ru/n104 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u437  (\cu_ru/n105 [36], \cu_ru/n103 [36], \cu_ru/n104 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u438  (\cu_ru/n105 [37], \cu_ru/n103 [37], \cu_ru/n104 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u439  (\cu_ru/n105 [38], \cu_ru/n103 [38], \cu_ru/n104 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  and \cu_ru/u44  (\cu_ru/n40 , \cu_ru/n39 , wb_int_acc);  // ../../RTL/CPU/CU&RU/cu_ru.v(345)
  or \cu_ru/u440  (\cu_ru/n105 [39], \cu_ru/n103 [39], \cu_ru/n104 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u441  (\cu_ru/n105 [40], \cu_ru/n103 [40], \cu_ru/n104 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u442  (\cu_ru/n105 [41], \cu_ru/n103 [41], \cu_ru/n104 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u443  (\cu_ru/n105 [42], \cu_ru/n103 [42], \cu_ru/n104 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u444  (\cu_ru/n105 [43], \cu_ru/n103 [43], \cu_ru/n104 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u445  (\cu_ru/n105 [44], \cu_ru/n103 [44], \cu_ru/n104 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u446  (\cu_ru/n105 [45], \cu_ru/n103 [45], \cu_ru/n104 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u447  (\cu_ru/n105 [46], \cu_ru/n103 [46], \cu_ru/n104 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u448  (\cu_ru/n105 [47], \cu_ru/n103 [47], \cu_ru/n104 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u449  (\cu_ru/n105 [48], \cu_ru/n103 [48], \cu_ru/n104 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  and \cu_ru/u45  (\cu_ru/n41 , wb_valid, \cu_ru/exc_target_s );  // ../../RTL/CPU/CU&RU/cu_ru.v(345)
  or \cu_ru/u450  (\cu_ru/n105 [49], \cu_ru/n103 [49], \cu_ru/n104 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u451  (\cu_ru/n105 [50], \cu_ru/n103 [50], \cu_ru/n104 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u452  (\cu_ru/n105 [51], \cu_ru/n103 [51], \cu_ru/n104 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u453  (\cu_ru/n105 [52], \cu_ru/n103 [52], \cu_ru/n104 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u454  (\cu_ru/n105 [53], \cu_ru/n103 [53], \cu_ru/n104 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u455  (\cu_ru/n105 [54], \cu_ru/n103 [54], \cu_ru/n104 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u456  (\cu_ru/n105 [55], \cu_ru/n103 [55], \cu_ru/n104 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u457  (\cu_ru/n105 [56], \cu_ru/n103 [56], \cu_ru/n104 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u458  (\cu_ru/n105 [57], \cu_ru/n103 [57], \cu_ru/n104 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u459  (\cu_ru/n105 [58], \cu_ru/n103 [58], \cu_ru/n104 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u46  (\cu_ru/trap_target_s , \cu_ru/n40 , \cu_ru/n41 );  // ../../RTL/CPU/CU&RU/cu_ru.v(345)
  or \cu_ru/u460  (\cu_ru/n105 [59], \cu_ru/n103 [59], \cu_ru/n104 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u461  (\cu_ru/n105 [60], \cu_ru/n103 [60], \cu_ru/n104 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u462  (\cu_ru/n105 [61], \cu_ru/n103 [61], \cu_ru/n104 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u463  (\cu_ru/n105 [62], \cu_ru/n103 [62], \cu_ru/n104 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u464  (\cu_ru/n105 [63], \cu_ru/n103 [63], \cu_ru/n104 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(698)
  or \cu_ru/u465  (\cu_ru/n103 [1], \cu_ru/n101 [1], \cu_ru/n102 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u466  (\cu_ru/n103 [2], \cu_ru/n101 [2], \cu_ru/n102 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u467  (\cu_ru/n103 [3], \cu_ru/n101 [3], \cu_ru/n102 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u468  (\cu_ru/n103 [4], \cu_ru/n101 [4], \cu_ru/n102 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u469  (\cu_ru/n103 [5], \cu_ru/n101 [5], \cu_ru/n102 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u47  (\cu_ru/n42 , wb_ebreak, \cu_ru/int_target_m );  // ../../RTL/CPU/CU&RU/cu_ru.v(349)
  or \cu_ru/u470  (\cu_ru/n103 [6], \cu_ru/n101 [6], \cu_ru/n102 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u471  (\cu_ru/n103 [7], \cu_ru/n101 [7], \cu_ru/n102 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u472  (\cu_ru/n103 [8], \cu_ru/n101 [8], \cu_ru/n102 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u473  (\cu_ru/n103 [9], \cu_ru/n101 [9], \cu_ru/n102 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u474  (\cu_ru/n103 [10], \cu_ru/n101 [10], \cu_ru/n102 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u475  (\cu_ru/n103 [11], \cu_ru/n101 [11], \cu_ru/n102 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u476  (\cu_ru/n103 [12], \cu_ru/n101 [12], \cu_ru/n102 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u477  (\cu_ru/n103 [13], \cu_ru/n101 [13], \cu_ru/n102 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u478  (\cu_ru/n103 [14], \cu_ru/n101 [14], \cu_ru/n102 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u479  (\cu_ru/n103 [15], \cu_ru/n101 [15], \cu_ru/n102 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u48  (\cu_ru/next_pc , \cu_ru/n42 , \cu_ru/int_target_s );  // ../../RTL/CPU/CU&RU/cu_ru.v(349)
  or \cu_ru/u480  (\cu_ru/n103 [16], \cu_ru/n101 [16], \cu_ru/n102 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u481  (\cu_ru/n103 [17], \cu_ru/n101 [17], \cu_ru/n102 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u482  (\cu_ru/n103 [18], \cu_ru/n101 [18], \cu_ru/n102 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u483  (\cu_ru/n103 [19], \cu_ru/n101 [19], \cu_ru/n102 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u484  (\cu_ru/n103 [20], \cu_ru/n101 [20], \cu_ru/n102 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u485  (\cu_ru/n103 [21], \cu_ru/n101 [21], \cu_ru/n102 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u486  (\cu_ru/n103 [22], \cu_ru/n101 [22], \cu_ru/n102 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u487  (\cu_ru/n103 [23], \cu_ru/n101 [23], \cu_ru/n102 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u488  (\cu_ru/n103 [24], \cu_ru/n101 [24], \cu_ru/n102 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u489  (\cu_ru/n103 [25], \cu_ru/n101 [25], \cu_ru/n102 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u49  (csr_data[1], \cu_ru/n113 [1], \cu_ru/n114 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u490  (\cu_ru/n103 [26], \cu_ru/n101 [26], \cu_ru/n102 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u491  (\cu_ru/n103 [27], \cu_ru/n101 [27], \cu_ru/n102 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u492  (\cu_ru/n103 [28], \cu_ru/n101 [28], \cu_ru/n102 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u493  (\cu_ru/n103 [29], \cu_ru/n101 [29], \cu_ru/n102 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u494  (\cu_ru/n103 [30], \cu_ru/n101 [30], \cu_ru/n102 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u495  (\cu_ru/n103 [31], \cu_ru/n101 [31], \cu_ru/n102 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u496  (\cu_ru/n103 [32], \cu_ru/n101 [32], \cu_ru/n102 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u497  (\cu_ru/n103 [33], \cu_ru/n101 [33], \cu_ru/n102 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u498  (\cu_ru/n103 [34], \cu_ru/n101 [34], \cu_ru/n102 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u499  (\cu_ru/n103 [35], \cu_ru/n101 [35], \cu_ru/n102 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  and \cu_ru/u5  (\cu_ru/srw_sscratch_sel , wb_valid, \cu_ru/n3 );  // ../../RTL/CPU/CU&RU/cu_ru.v(268)
  or \cu_ru/u50  (csr_data[2], \cu_ru/n113 [2], \cu_ru/n114 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u500  (\cu_ru/n103 [36], \cu_ru/n101 [36], \cu_ru/n102 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u501  (\cu_ru/n103 [37], \cu_ru/n101 [37], \cu_ru/n102 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u502  (\cu_ru/n103 [38], \cu_ru/n101 [38], \cu_ru/n102 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u503  (\cu_ru/n103 [39], \cu_ru/n101 [39], \cu_ru/n102 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u504  (\cu_ru/n103 [40], \cu_ru/n101 [40], \cu_ru/n102 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u505  (\cu_ru/n103 [41], \cu_ru/n101 [41], \cu_ru/n102 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u506  (\cu_ru/n103 [42], \cu_ru/n101 [42], \cu_ru/n102 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u507  (\cu_ru/n103 [43], \cu_ru/n101 [43], \cu_ru/n102 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u508  (\cu_ru/n103 [44], \cu_ru/n101 [44], \cu_ru/n102 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u509  (\cu_ru/n103 [45], \cu_ru/n101 [45], \cu_ru/n102 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u51  (csr_data[3], \cu_ru/n113 [3], \cu_ru/n114 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u510  (\cu_ru/n103 [46], \cu_ru/n101 [46], \cu_ru/n102 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u511  (\cu_ru/n103 [47], \cu_ru/n101 [47], \cu_ru/n102 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u512  (\cu_ru/n103 [48], \cu_ru/n101 [48], \cu_ru/n102 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u513  (\cu_ru/n103 [49], \cu_ru/n101 [49], \cu_ru/n102 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u514  (\cu_ru/n103 [50], \cu_ru/n101 [50], \cu_ru/n102 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u515  (\cu_ru/n103 [51], \cu_ru/n101 [51], \cu_ru/n102 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u516  (\cu_ru/n103 [52], \cu_ru/n101 [52], \cu_ru/n102 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u517  (\cu_ru/n103 [53], \cu_ru/n101 [53], \cu_ru/n102 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u518  (\cu_ru/n103 [54], \cu_ru/n101 [54], \cu_ru/n102 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u519  (\cu_ru/n103 [55], \cu_ru/n101 [55], \cu_ru/n102 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u52  (csr_data[4], \cu_ru/n113 [4], \cu_ru/n114 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u520  (\cu_ru/n103 [56], \cu_ru/n101 [56], \cu_ru/n102 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u521  (\cu_ru/n103 [57], \cu_ru/n101 [57], \cu_ru/n102 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u522  (\cu_ru/n103 [58], \cu_ru/n101 [58], \cu_ru/n102 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u523  (\cu_ru/n103 [59], \cu_ru/n101 [59], \cu_ru/n102 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u524  (\cu_ru/n103 [60], \cu_ru/n101 [60], \cu_ru/n102 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u525  (\cu_ru/n103 [61], \cu_ru/n101 [61], \cu_ru/n102 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u526  (\cu_ru/n103 [62], \cu_ru/n101 [62], \cu_ru/n102 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u527  (\cu_ru/n103 [63], \cu_ru/n101 [63], \cu_ru/n102 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(697)
  or \cu_ru/u528  (\cu_ru/n101 [1], \cu_ru/n97 [1], \cu_ru/n100 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u529  (\cu_ru/n101 [2], \cu_ru/n95 [2], \cu_ru/n100 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u53  (csr_data[5], \cu_ru/n113 [5], \cu_ru/n114 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u530  (\cu_ru/n101 [3], \cu_ru/n95 [3], \cu_ru/n100 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u531  (\cu_ru/n101 [4], \cu_ru/n95 [4], \cu_ru/n100 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u532  (\cu_ru/n101 [5], \cu_ru/n97 [5], \cu_ru/n100 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u533  (\cu_ru/n101 [6], \cu_ru/n95 [6], \cu_ru/n100 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u534  (\cu_ru/n101 [7], \cu_ru/n95 [7], \cu_ru/n100 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u535  (\cu_ru/n101 [8], \cu_ru/n95 [8], \cu_ru/n100 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u536  (\cu_ru/n101 [9], \cu_ru/n97 [9], \cu_ru/n100 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u537  (\cu_ru/n101 [10], \cu_ru/n85 [10], \cu_ru/n100 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u538  (\cu_ru/n101 [11], \cu_ru/n91 [11], \cu_ru/n100 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u539  (\cu_ru/n101 [12], \cu_ru/n95 [12], \cu_ru/n100 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u54  (csr_data[6], \cu_ru/n113 [6], \cu_ru/n114 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u540  (\cu_ru/n101 [13], \cu_ru/n95 [13], \cu_ru/n100 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u541  (\cu_ru/n101 [14], \cu_ru/n85 [14], \cu_ru/n100 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u542  (\cu_ru/n101 [15], \cu_ru/n95 [15], \cu_ru/n100 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u543  (\cu_ru/n101 [16], \cu_ru/n81 [16], \cu_ru/n100 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u544  (\cu_ru/n101 [17], \cu_ru/n91 [17], \cu_ru/n100 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u545  (\cu_ru/n101 [18], \cu_ru/n91 [18], \cu_ru/n100 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u546  (\cu_ru/n101 [19], \cu_ru/n91 [19], \cu_ru/n100 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u547  (\cu_ru/n101 [20], \cu_ru/n91 [20], \cu_ru/n100 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u548  (\cu_ru/n101 [21], \cu_ru/n91 [21], \cu_ru/n100 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u549  (\cu_ru/n101 [22], \cu_ru/n91 [22], \cu_ru/n100 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u55  (csr_data[7], \cu_ru/n113 [7], \cu_ru/n114 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u550  (\cu_ru/n101 [23], \cu_ru/n81 [23], \cu_ru/n100 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u551  (\cu_ru/n101 [24], \cu_ru/n81 [24], \cu_ru/n100 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u552  (\cu_ru/n101 [25], \cu_ru/n83 [25], \cu_ru/n100 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u553  (\cu_ru/n101 [26], \cu_ru/n81 [26], \cu_ru/n100 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u554  (\cu_ru/n101 [27], \cu_ru/n81 [27], \cu_ru/n100 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u555  (\cu_ru/n101 [28], \cu_ru/n85 [28], \cu_ru/n100 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u556  (\cu_ru/n101 [29], \cu_ru/n81 [29], \cu_ru/n100 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u557  (\cu_ru/n101 [30], \cu_ru/n85 [30], \cu_ru/n100 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u558  (\cu_ru/n101 [31], \cu_ru/n81 [31], \cu_ru/n100 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u559  (\cu_ru/n101 [32], \cu_ru/n91 [32], \cu_ru/n100 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u56  (csr_data[8], \cu_ru/n113 [8], \cu_ru/n114 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u560  (\cu_ru/n101 [33], \cu_ru/n91 [33], \cu_ru/n100 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u561  (\cu_ru/n101 [34], \cu_ru/n91 [34], \cu_ru/n100 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u562  (\cu_ru/n101 [35], \cu_ru/n91 [35], \cu_ru/n100 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u563  (\cu_ru/n101 [36], \cu_ru/n81 [36], \cu_ru/n100 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u564  (\cu_ru/n101 [37], \cu_ru/n81 [37], \cu_ru/n100 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u565  (\cu_ru/n101 [38], \cu_ru/n81 [38], \cu_ru/n100 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u566  (\cu_ru/n101 [39], \cu_ru/n81 [39], \cu_ru/n100 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u567  (\cu_ru/n101 [40], \cu_ru/n81 [40], \cu_ru/n100 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u568  (\cu_ru/n101 [41], \cu_ru/n81 [41], \cu_ru/n100 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u569  (\cu_ru/n101 [42], \cu_ru/n81 [42], \cu_ru/n100 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u57  (csr_data[9], \cu_ru/n113 [9], \cu_ru/n114 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u570  (\cu_ru/n101 [43], \cu_ru/n81 [43], \cu_ru/n100 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u571  (\cu_ru/n101 [44], \cu_ru/n77 [44], \cu_ru/n100 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u572  (\cu_ru/n101 [45], \cu_ru/n77 [45], \cu_ru/n100 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u573  (\cu_ru/n101 [46], \cu_ru/n77 [46], \cu_ru/n100 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u574  (\cu_ru/n101 [47], \cu_ru/n77 [47], \cu_ru/n100 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u575  (\cu_ru/n101 [48], \cu_ru/n77 [48], \cu_ru/n100 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u576  (\cu_ru/n101 [49], \cu_ru/n77 [49], \cu_ru/n100 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u577  (\cu_ru/n101 [50], \cu_ru/n77 [50], \cu_ru/n100 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u578  (\cu_ru/n101 [51], \cu_ru/n77 [51], \cu_ru/n100 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u579  (\cu_ru/n101 [52], \cu_ru/n77 [52], \cu_ru/n100 [52]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u58  (csr_data[10], \cu_ru/n113 [10], \cu_ru/n114 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u580  (\cu_ru/n101 [53], \cu_ru/n77 [53], \cu_ru/n100 [53]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u581  (\cu_ru/n101 [54], \cu_ru/n77 [54], \cu_ru/n100 [54]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u582  (\cu_ru/n101 [55], \cu_ru/n77 [55], \cu_ru/n100 [55]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u583  (\cu_ru/n101 [56], \cu_ru/n77 [56], \cu_ru/n100 [56]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u584  (\cu_ru/n101 [57], \cu_ru/n77 [57], \cu_ru/n100 [57]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u585  (\cu_ru/n101 [58], \cu_ru/n77 [58], \cu_ru/n100 [58]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u586  (\cu_ru/n101 [59], \cu_ru/n77 [59], \cu_ru/n100 [59]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u587  (\cu_ru/n101 [60], \cu_ru/n81 [60], \cu_ru/n100 [60]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u588  (\cu_ru/n101 [61], \cu_ru/n81 [61], \cu_ru/n100 [61]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u589  (\cu_ru/n101 [62], \cu_ru/n81 [62], \cu_ru/n100 [62]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u59  (csr_data[11], \cu_ru/n113 [11], \cu_ru/n114 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u590  (\cu_ru/n101 [63], \cu_ru/n81 [63], \cu_ru/n100 [63]);  // ../../RTL/CPU/CU&RU/cu_ru.v(695)
  or \cu_ru/u591  (\cu_ru/n97 [1], \cu_ru/n95 [1], \cu_ru/n96 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(693)
  or \cu_ru/u595  (\cu_ru/n97 [5], \cu_ru/n95 [5], \cu_ru/n96 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(693)
  or \cu_ru/u599  (\cu_ru/n97 [9], \cu_ru/n95 [9], \cu_ru/n96 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(693)
  and \cu_ru/u6  (\cu_ru/srw_sepc_sel , wb_valid, \cu_ru/n4 );  // ../../RTL/CPU/CU&RU/cu_ru.v(269)
  or \cu_ru/u60  (csr_data[12], \cu_ru/n113 [12], \cu_ru/n114 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u61  (csr_data[13], \cu_ru/n113 [13], \cu_ru/n114 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u62  (csr_data[14], \cu_ru/n113 [14], \cu_ru/n114 [14]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u63  (csr_data[15], \cu_ru/n113 [15], \cu_ru/n114 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u64  (csr_data[16], \cu_ru/n113 [16], \cu_ru/n114 [16]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u65  (csr_data[17], \cu_ru/n113 [17], \cu_ru/n114 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u654  (\cu_ru/n95 [1], \cu_ru/n91 [1], \cu_ru/n94 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u655  (\cu_ru/n95 [2], \cu_ru/n87 [2], \cu_ru/n94 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u656  (\cu_ru/n95 [3], \cu_ru/n91 [3], \cu_ru/n94 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u657  (\cu_ru/n95 [4], \cu_ru/n85 [4], \cu_ru/n94 [4]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u658  (\cu_ru/n95 [5], \cu_ru/n91 [5], \cu_ru/n94 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u659  (\cu_ru/n95 [6], \cu_ru/n83 [6], \cu_ru/n94 [6]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u66  (csr_data[18], \cu_ru/n113 [18], \cu_ru/n114 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u660  (\cu_ru/n95 [7], \cu_ru/n91 [7], \cu_ru/n94 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u661  (\cu_ru/n95 [8], \cu_ru/n91 [8], \cu_ru/n94 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u662  (\cu_ru/n95 [9], \cu_ru/n85 [9], \cu_ru/n94 [9]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u665  (\cu_ru/n95 [12], \cu_ru/n91 [12], \cu_ru/n94 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u666  (\cu_ru/n95 [13], \cu_ru/n81 [13], \cu_ru/n94 [13]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u668  (\cu_ru/n95 [15], \cu_ru/n81 [15], \cu_ru/n94 [15]);  // ../../RTL/CPU/CU&RU/cu_ru.v(692)
  or \cu_ru/u67  (csr_data[19], \cu_ru/n113 [19], \cu_ru/n114 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u68  (csr_data[20], \cu_ru/n113 [20], \cu_ru/n114 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u69  (csr_data[21], \cu_ru/n113 [21], \cu_ru/n114 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  and \cu_ru/u7  (\cu_ru/srw_scause_sel , wb_valid, \cu_ru/n5 );  // ../../RTL/CPU/CU&RU/cu_ru.v(270)
  or \cu_ru/u70  (csr_data[22], \cu_ru/n113 [22], \cu_ru/n114 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u71  (csr_data[23], \cu_ru/n113 [23], \cu_ru/n114 [23]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u72  (csr_data[24], \cu_ru/n113 [24], \cu_ru/n114 [24]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u73  (csr_data[25], \cu_ru/n113 [25], \cu_ru/n114 [25]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u74  (csr_data[26], \cu_ru/n113 [26], \cu_ru/n114 [26]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u75  (csr_data[27], \cu_ru/n113 [27], \cu_ru/n114 [27]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u76  (csr_data[28], \cu_ru/n113 [28], \cu_ru/n114 [28]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u77  (csr_data[29], \cu_ru/n113 [29], \cu_ru/n114 [29]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u78  (csr_data[30], \cu_ru/n113 [30], \cu_ru/n114 [30]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u780  (\cu_ru/n91 [1], \cu_ru/n81 [1], \cu_ru/n90 [1]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u782  (\cu_ru/n91 [3], \cu_ru/n81 [3], \cu_ru/n90 [3]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u784  (\cu_ru/n91 [5], \cu_ru/n85 [5], \cu_ru/n90 [5]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u786  (\cu_ru/n91 [7], \cu_ru/n81 [7], \cu_ru/n90 [7]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u787  (\cu_ru/n91 [8], \cu_ru/n83 [8], \cu_ru/n90 [8]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u79  (csr_data[31], \cu_ru/n113 [31], \cu_ru/n114 [31]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u790  (\cu_ru/n91 [11], \cu_ru/n81 [11], \cu_ru/n90 [11]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u791  (\cu_ru/n91 [12], \cu_ru/n85 [12], \cu_ru/n90 [12]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u796  (\cu_ru/n91 [17], \cu_ru/n85 [17], \cu_ru/n90 [17]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u797  (\cu_ru/n91 [18], \cu_ru/n83 [18], \cu_ru/n90 [18]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u798  (\cu_ru/n91 [19], \cu_ru/n81 [19], \cu_ru/n90 [19]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u799  (\cu_ru/n91 [20], \cu_ru/n85 [20], \cu_ru/n90 [20]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  and \cu_ru/u8  (\cu_ru/srw_stval_sel , wb_valid, \cu_ru/n6 );  // ../../RTL/CPU/CU&RU/cu_ru.v(271)
  or \cu_ru/u80  (csr_data[32], \cu_ru/n113 [32], \cu_ru/n114 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u800  (\cu_ru/n91 [21], \cu_ru/n81 [21], \cu_ru/n90 [21]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u801  (\cu_ru/n91 [22], \cu_ru/n85 [22], \cu_ru/n90 [22]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u81  (csr_data[33], \cu_ru/n113 [33], \cu_ru/n114 [33]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u811  (\cu_ru/n91 [32], \cu_ru/n81 [32], \cu_ru/n90 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u812  (\cu_ru/n91 [33], \cu_ru/n81 [33], \cu_ru/n90 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u813  (\cu_ru/n91 [34], \cu_ru/n81 [34], \cu_ru/n90 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u814  (\cu_ru/n91 [35], \cu_ru/n81 [35], \cu_ru/n90 [32]);  // ../../RTL/CPU/CU&RU/cu_ru.v(690)
  or \cu_ru/u82  (csr_data[34], \cu_ru/n113 [34], \cu_ru/n114 [34]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u83  (csr_data[35], \cu_ru/n113 [35], \cu_ru/n114 [35]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u84  (csr_data[36], \cu_ru/n113 [36], \cu_ru/n114 [36]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u85  (csr_data[37], \cu_ru/n113 [37], \cu_ru/n114 [37]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u86  (csr_data[38], \cu_ru/n113 [38], \cu_ru/n114 [38]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u87  (csr_data[39], \cu_ru/n113 [39], \cu_ru/n114 [39]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u88  (csr_data[40], \cu_ru/n113 [40], \cu_ru/n114 [40]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u89  (csr_data[41], \cu_ru/n113 [41], \cu_ru/n114 [41]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  and \cu_ru/u9  (\cu_ru/srw_sip_sel , wb_valid, \cu_ru/n7 );  // ../../RTL/CPU/CU&RU/cu_ru.v(272)
  or \cu_ru/u90  (csr_data[42], \cu_ru/n113 [42], \cu_ru/n114 [42]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u907  (\cu_ru/n87 [2], \cu_ru/n85 [2], \cu_ru/n86 [2]);  // ../../RTL/CPU/CU&RU/cu_ru.v(688)
  or \cu_ru/u91  (csr_data[43], \cu_ru/n113 [43], \cu_ru/n114 [43]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u92  (csr_data[44], \cu_ru/n113 [44], \cu_ru/n114 [44]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u93  (csr_data[45], \cu_ru/n113 [45], \cu_ru/n114 [45]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u94  (csr_data[46], \cu_ru/n113 [46], \cu_ru/n114 [46]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u95  (csr_data[47], \cu_ru/n113 [47], \cu_ru/n114 [47]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u96  (csr_data[48], \cu_ru/n113 [48], \cu_ru/n114 [48]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u97  (csr_data[49], \cu_ru/n113 [49], \cu_ru/n114 [49]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u970  (\cu_ru/n85 [2], \cu_ru/n83 [2], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u972  (\cu_ru/n85 [4], \cu_ru/n83 [4], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u973  (\cu_ru/n85 [5], \cu_ru/n81 [5], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u977  (\cu_ru/n85 [9], \cu_ru/n81 [9], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u978  (\cu_ru/n85 [10], \cu_ru/n81 [10], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u98  (csr_data[50], \cu_ru/n113 [50], \cu_ru/n114 [50]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u980  (\cu_ru/n85 [12], \cu_ru/n81 [12], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u982  (\cu_ru/n85 [14], \cu_ru/n83 [14], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u985  (\cu_ru/n85 [17], \cu_ru/n83 [17], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u988  (\cu_ru/n85 [20], \cu_ru/n83 [20], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u99  (csr_data[51], \cu_ru/n113 [51], \cu_ru/n114 [51]);  // ../../RTL/CPU/CU&RU/cu_ru.v(704)
  or \cu_ru/u990  (\cu_ru/n85 [22], \cu_ru/n83 [22], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u996  (\cu_ru/n85 [28], \cu_ru/n83 [28], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  or \cu_ru/u998  (\cu_ru/n85 [30], \cu_ru/n83 [30], \cu_ru/n84 [10]);  // ../../RTL/CPU/CU&RU/cu_ru.v(687)
  not ex_more_exception_inv (ex_more_exception_neg, ex_more_exception);
  not \ex_size[2]_inv  (\ex_size[2]_neg , ex_size[2]);
  add_pu64_pu64_o64 \exu/alu_au/add0  (
    .i0(ds1),
    .i1(\exu/alu_au/n17 ),
    .o(\exu/alu_au/add_64 ));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  add_pu32_pu32_o32 \exu/alu_au/add1  (
    .i0(\exu/alu_au/add_64 [31:0]),
    .i1(32'b00000000000000000000000000000001),
    .o(\exu/alu_au/sub_64 [31:0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(80)
  add_pu64_pu64_o64 \exu/alu_au/add2  (
    .i0(as1),
    .i1({as2[56],as2[56],as2[56],as2[56],as2[56],as2[56],as2[56],as2[56],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20],as2[20:0]}),
    .o(addr_ex));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(118)
  lt_u64_u64 \exu/alu_au/lt0  (
    .ci(1'b0),
    .i0(ds1),
    .i1(ds2),
    .o(\exu/alu_au/n5 ));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(72)
  lt_u64_u64 \exu/alu_au/lt1  (
    .ci(1'b0),
    .i0(ds2),
    .i1(ds1),
    .o(\exu/alu_au/n12 ));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(75)
  binary_mux_s1_w1 \exu/alu_au/mux0_b0  (
    .i0(ds2[0]),
    .i1(\exu/alu_au/n16 [0]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b1  (
    .i0(ds2[1]),
    .i1(\exu/alu_au/n16 [1]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b10  (
    .i0(ds2[10]),
    .i1(\exu/alu_au/n16 [10]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b11  (
    .i0(ds2[11]),
    .i1(\exu/alu_au/n16 [11]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b12  (
    .i0(ds2[12]),
    .i1(\exu/alu_au/n16 [12]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b13  (
    .i0(ds2[13]),
    .i1(\exu/alu_au/n16 [13]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b14  (
    .i0(ds2[14]),
    .i1(\exu/alu_au/n16 [14]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b15  (
    .i0(ds2[15]),
    .i1(\exu/alu_au/n16 [15]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b16  (
    .i0(ds2[16]),
    .i1(\exu/alu_au/n16 [16]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b17  (
    .i0(ds2[17]),
    .i1(\exu/alu_au/n16 [17]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b18  (
    .i0(ds2[18]),
    .i1(\exu/alu_au/n16 [18]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b19  (
    .i0(ds2[19]),
    .i1(\exu/alu_au/n16 [19]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b2  (
    .i0(ds2[2]),
    .i1(\exu/alu_au/n16 [2]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b20  (
    .i0(ds2[20]),
    .i1(\exu/alu_au/n16 [20]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b21  (
    .i0(ds2[21]),
    .i1(\exu/alu_au/n16 [21]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b22  (
    .i0(ds2[22]),
    .i1(\exu/alu_au/n16 [22]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b23  (
    .i0(ds2[23]),
    .i1(\exu/alu_au/n16 [23]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b24  (
    .i0(ds2[24]),
    .i1(\exu/alu_au/n16 [24]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b25  (
    .i0(ds2[25]),
    .i1(\exu/alu_au/n16 [25]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b26  (
    .i0(ds2[26]),
    .i1(\exu/alu_au/n16 [26]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b27  (
    .i0(ds2[27]),
    .i1(\exu/alu_au/n16 [27]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b28  (
    .i0(ds2[28]),
    .i1(\exu/alu_au/n16 [28]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b29  (
    .i0(ds2[29]),
    .i1(\exu/alu_au/n16 [29]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b3  (
    .i0(ds2[3]),
    .i1(\exu/alu_au/n16 [3]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b30  (
    .i0(ds2[30]),
    .i1(\exu/alu_au/n16 [30]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b31  (
    .i0(ds2[31]),
    .i1(\exu/alu_au/n16 [31]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b32  (
    .i0(ds2[32]),
    .i1(\exu/alu_au/n16 [32]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b33  (
    .i0(ds2[33]),
    .i1(\exu/alu_au/n16 [33]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b34  (
    .i0(ds2[34]),
    .i1(\exu/alu_au/n16 [34]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b35  (
    .i0(ds2[35]),
    .i1(\exu/alu_au/n16 [35]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b36  (
    .i0(ds2[36]),
    .i1(\exu/alu_au/n16 [36]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b37  (
    .i0(ds2[37]),
    .i1(\exu/alu_au/n16 [37]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b38  (
    .i0(ds2[38]),
    .i1(\exu/alu_au/n16 [38]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b39  (
    .i0(ds2[39]),
    .i1(\exu/alu_au/n16 [39]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b4  (
    .i0(ds2[4]),
    .i1(\exu/alu_au/n16 [4]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b40  (
    .i0(ds2[40]),
    .i1(\exu/alu_au/n16 [40]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b41  (
    .i0(ds2[41]),
    .i1(\exu/alu_au/n16 [41]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b42  (
    .i0(ds2[42]),
    .i1(\exu/alu_au/n16 [42]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b43  (
    .i0(ds2[43]),
    .i1(\exu/alu_au/n16 [43]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b44  (
    .i0(ds2[44]),
    .i1(\exu/alu_au/n16 [44]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b45  (
    .i0(ds2[45]),
    .i1(\exu/alu_au/n16 [45]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b46  (
    .i0(ds2[46]),
    .i1(\exu/alu_au/n16 [46]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b47  (
    .i0(ds2[47]),
    .i1(\exu/alu_au/n16 [47]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b48  (
    .i0(ds2[48]),
    .i1(\exu/alu_au/n16 [48]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b49  (
    .i0(ds2[49]),
    .i1(\exu/alu_au/n16 [49]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b5  (
    .i0(ds2[5]),
    .i1(\exu/alu_au/n16 [5]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b50  (
    .i0(ds2[50]),
    .i1(\exu/alu_au/n16 [50]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b51  (
    .i0(ds2[51]),
    .i1(\exu/alu_au/n16 [51]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b52  (
    .i0(ds2[52]),
    .i1(\exu/alu_au/n16 [52]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b53  (
    .i0(ds2[53]),
    .i1(\exu/alu_au/n16 [53]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b54  (
    .i0(ds2[54]),
    .i1(\exu/alu_au/n16 [54]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b55  (
    .i0(ds2[55]),
    .i1(\exu/alu_au/n16 [55]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b56  (
    .i0(ds2[56]),
    .i1(\exu/alu_au/n16 [56]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b57  (
    .i0(ds2[57]),
    .i1(\exu/alu_au/n16 [57]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b58  (
    .i0(ds2[58]),
    .i1(\exu/alu_au/n16 [58]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b59  (
    .i0(ds2[59]),
    .i1(\exu/alu_au/n16 [59]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b6  (
    .i0(ds2[6]),
    .i1(\exu/alu_au/n16 [6]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b60  (
    .i0(ds2[60]),
    .i1(\exu/alu_au/n16 [60]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b61  (
    .i0(ds2[61]),
    .i1(\exu/alu_au/n16 [61]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b62  (
    .i0(ds2[62]),
    .i1(\exu/alu_au/n16 [62]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b63  (
    .i0(ds2[63]),
    .i1(\exu/alu_au/n16 [63]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b7  (
    .i0(ds2[7]),
    .i1(\exu/alu_au/n16 [7]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b8  (
    .i0(ds2[8]),
    .i1(\exu/alu_au/n16 [8]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux0_b9  (
    .i0(ds2[9]),
    .i1(\exu/alu_au/n16 [9]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n17 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  binary_mux_s1_w1 \exu/alu_au/mux10_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [0]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [1]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [10]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [11]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [12]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [13]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [14]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [15]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [16]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [17]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [18]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [19]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [2]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [20]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [21]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [22]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [23]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [24]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [25]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [26]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [27]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [28]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [29]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [3]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [30]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [31]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [32]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [33]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [34]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [35]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [36]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [37]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [38]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [39]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [4]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [40]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [41]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [42]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [43]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [44]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [45]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [46]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [47]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [48]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [49]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [5]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [50]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [51]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [52]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [53]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [54]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [55]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [56]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [57]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [58]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [59]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [6]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [60]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [61]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [62]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [63]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [7]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [8]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux10_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [9]),
    .sel(rd_data_or),
    .o(\exu/alu_au/n35 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  binary_mux_s1_w1 \exu/alu_au/mux11_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [0]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [1]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [10]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [11]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [12]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [13]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [14]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [15]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [16]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [17]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [18]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [19]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [2]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [20]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [21]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [22]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [23]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [24]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [25]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [26]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [27]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [28]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [29]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [3]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [30]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [31]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [32]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [33]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [34]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [35]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [36]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [37]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [38]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [39]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [4]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [40]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [41]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [42]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [43]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [44]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [45]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [46]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [47]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [48]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [49]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [5]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [50]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [51]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [52]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [53]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [54]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [55]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [56]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [57]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [58]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [59]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [6]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [60]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [61]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [62]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [63]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [7]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [8]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux11_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [9]),
    .sel(rd_data_xor),
    .o(\exu/alu_au/n37 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  binary_mux_s1_w1 \exu/alu_au/mux12_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/ds1_light_than_ds2 ),
    .sel(rd_data_slt),
    .o(\exu/alu_au/n39 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(105)
  binary_mux_s1_w1 \exu/alu_au/mux15_b0  (
    .i0(1'b0),
    .i1(ds2[0]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b1  (
    .i0(1'b0),
    .i1(ds2[1]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b10  (
    .i0(1'b0),
    .i1(ds2[10]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b11  (
    .i0(1'b0),
    .i1(ds2[11]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b12  (
    .i0(1'b0),
    .i1(ds2[12]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b13  (
    .i0(1'b0),
    .i1(ds2[13]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b14  (
    .i0(1'b0),
    .i1(ds2[14]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b15  (
    .i0(1'b0),
    .i1(ds2[15]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b16  (
    .i0(1'b0),
    .i1(ds2[16]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b17  (
    .i0(1'b0),
    .i1(ds2[17]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b18  (
    .i0(1'b0),
    .i1(ds2[18]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b19  (
    .i0(1'b0),
    .i1(ds2[19]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b2  (
    .i0(1'b0),
    .i1(ds2[2]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b20  (
    .i0(1'b0),
    .i1(ds2[20]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b21  (
    .i0(1'b0),
    .i1(ds2[21]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b22  (
    .i0(1'b0),
    .i1(ds2[22]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b23  (
    .i0(1'b0),
    .i1(ds2[23]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b24  (
    .i0(1'b0),
    .i1(ds2[24]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b25  (
    .i0(1'b0),
    .i1(ds2[25]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b26  (
    .i0(1'b0),
    .i1(ds2[26]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b27  (
    .i0(1'b0),
    .i1(ds2[27]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b28  (
    .i0(1'b0),
    .i1(ds2[28]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b29  (
    .i0(1'b0),
    .i1(ds2[29]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b3  (
    .i0(1'b0),
    .i1(ds2[3]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b30  (
    .i0(1'b0),
    .i1(ds2[30]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b31  (
    .i0(1'b0),
    .i1(ds2[31]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b32  (
    .i0(1'b0),
    .i1(ds2[32]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b33  (
    .i0(1'b0),
    .i1(ds2[33]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b34  (
    .i0(1'b0),
    .i1(ds2[34]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b35  (
    .i0(1'b0),
    .i1(ds2[35]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b36  (
    .i0(1'b0),
    .i1(ds2[36]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b37  (
    .i0(1'b0),
    .i1(ds2[37]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b38  (
    .i0(1'b0),
    .i1(ds2[38]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b39  (
    .i0(1'b0),
    .i1(ds2[39]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b4  (
    .i0(1'b0),
    .i1(ds2[4]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b40  (
    .i0(1'b0),
    .i1(ds2[40]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b41  (
    .i0(1'b0),
    .i1(ds2[41]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b42  (
    .i0(1'b0),
    .i1(ds2[42]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b43  (
    .i0(1'b0),
    .i1(ds2[43]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b44  (
    .i0(1'b0),
    .i1(ds2[44]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b45  (
    .i0(1'b0),
    .i1(ds2[45]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b46  (
    .i0(1'b0),
    .i1(ds2[46]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b47  (
    .i0(1'b0),
    .i1(ds2[47]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b48  (
    .i0(1'b0),
    .i1(ds2[48]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b49  (
    .i0(1'b0),
    .i1(ds2[49]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b5  (
    .i0(1'b0),
    .i1(ds2[5]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b50  (
    .i0(1'b0),
    .i1(ds2[50]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b51  (
    .i0(1'b0),
    .i1(ds2[51]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b52  (
    .i0(1'b0),
    .i1(ds2[52]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b53  (
    .i0(1'b0),
    .i1(ds2[53]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b54  (
    .i0(1'b0),
    .i1(ds2[54]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b55  (
    .i0(1'b0),
    .i1(ds2[55]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b56  (
    .i0(1'b0),
    .i1(ds2[56]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b57  (
    .i0(1'b0),
    .i1(ds2[57]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b58  (
    .i0(1'b0),
    .i1(ds2[58]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b59  (
    .i0(1'b0),
    .i1(ds2[59]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b6  (
    .i0(1'b0),
    .i1(ds2[6]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b60  (
    .i0(1'b0),
    .i1(ds2[60]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b61  (
    .i0(1'b0),
    .i1(ds2[61]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b62  (
    .i0(1'b0),
    .i1(ds2[62]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b63  (
    .i0(1'b0),
    .i1(ds2[63]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b7  (
    .i0(1'b0),
    .i1(ds2[7]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b8  (
    .i0(1'b0),
    .i1(ds2[8]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux15_b9  (
    .i0(1'b0),
    .i1(ds2[9]),
    .sel(mem_csr_data_ds2),
    .o(\exu/alu_au/n43 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(110)
  binary_mux_s1_w1 \exu/alu_au/mux16_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [0]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [1]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [10]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [11]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [12]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [13]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [14]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [15]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [16]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [17]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [18]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [19]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [2]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [20]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [21]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [22]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [23]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [24]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [25]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [26]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [27]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [28]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [29]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [3]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [30]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [32]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [33]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [34]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [35]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [36]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [37]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [38]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [39]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [4]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [40]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [41]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [42]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [43]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [44]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [45]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [46]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [47]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [48]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [49]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [5]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [50]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [51]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [52]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [53]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [54]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [55]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [56]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [57]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [58]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [59]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [6]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [60]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [61]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [62]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [63]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [7]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [8]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux16_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [9]),
    .sel(mem_csr_data_add),
    .o(\exu/alu_au/n45 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  binary_mux_s1_w1 \exu/alu_au/mux17_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [0]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [1]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [10]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [11]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [12]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [13]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [14]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [15]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [16]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [17]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [18]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [19]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [2]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [20]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [21]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [22]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [23]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [24]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [25]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [26]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [27]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [28]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [29]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [3]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [30]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [31]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [32]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [33]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [34]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [35]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [36]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [37]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [38]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [39]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [4]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [40]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [41]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [42]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [43]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [44]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [45]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [46]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [47]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [48]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [49]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [5]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [50]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [51]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [52]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [53]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [54]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [55]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [56]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [57]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [58]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [59]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [6]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [60]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [61]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [62]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [63]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [7]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [8]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux17_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [9]),
    .sel(mem_csr_data_and),
    .o(\exu/alu_au/n47 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  binary_mux_s1_w1 \exu/alu_au/mux18_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [0]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [1]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [10]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [11]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [12]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [13]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [14]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [15]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [16]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [17]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [18]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [19]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [2]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [20]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [21]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [22]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [23]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [24]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [25]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [26]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [27]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [28]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [29]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [3]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [30]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [31]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [32]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [33]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [34]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [35]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [36]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [37]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [38]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [39]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [4]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [40]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [41]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [42]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [43]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [44]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [45]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [46]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [47]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [48]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [49]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [5]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [50]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [51]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [52]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [53]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [54]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [55]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [56]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [57]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [58]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [59]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [6]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [60]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [61]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [62]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [63]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [7]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [8]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux18_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_or [9]),
    .sel(mem_csr_data_or),
    .o(\exu/alu_au/n49 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  binary_mux_s1_w1 \exu/alu_au/mux19_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [0]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [1]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [10]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [11]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [12]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [13]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [14]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [15]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [16]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [17]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [18]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [19]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [2]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [20]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [21]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [22]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [23]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [24]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [25]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [26]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [27]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [28]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [29]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [3]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [30]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [31]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [32]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [33]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [34]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [35]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [36]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [37]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [38]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [39]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [4]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [40]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [41]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [42]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [43]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [44]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [45]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [46]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [47]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [48]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [49]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [5]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [50]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [51]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [52]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [53]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [54]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [55]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [56]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [57]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [58]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [59]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [6]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [60]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [61]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [62]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [63]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [7]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [8]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux19_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_xor [9]),
    .sel(mem_csr_data_xor),
    .o(\exu/alu_au/n51 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  binary_mux_s1_w1 \exu/alu_au/mux1_b0  (
    .i0(\exu/alu_au/add_64 [32]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b1  (
    .i0(\exu/alu_au/add_64 [33]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b10  (
    .i0(\exu/alu_au/add_64 [42]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b11  (
    .i0(\exu/alu_au/add_64 [43]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b12  (
    .i0(\exu/alu_au/add_64 [44]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b13  (
    .i0(\exu/alu_au/add_64 [45]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b14  (
    .i0(\exu/alu_au/add_64 [46]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b15  (
    .i0(\exu/alu_au/add_64 [47]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b16  (
    .i0(\exu/alu_au/add_64 [48]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b17  (
    .i0(\exu/alu_au/add_64 [49]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b18  (
    .i0(\exu/alu_au/add_64 [50]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b19  (
    .i0(\exu/alu_au/add_64 [51]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b2  (
    .i0(\exu/alu_au/add_64 [34]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b20  (
    .i0(\exu/alu_au/add_64 [52]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b21  (
    .i0(\exu/alu_au/add_64 [53]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b22  (
    .i0(\exu/alu_au/add_64 [54]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b23  (
    .i0(\exu/alu_au/add_64 [55]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b24  (
    .i0(\exu/alu_au/add_64 [56]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b25  (
    .i0(\exu/alu_au/add_64 [57]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b26  (
    .i0(\exu/alu_au/add_64 [58]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b27  (
    .i0(\exu/alu_au/add_64 [59]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b28  (
    .i0(\exu/alu_au/add_64 [60]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b29  (
    .i0(\exu/alu_au/add_64 [61]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b3  (
    .i0(\exu/alu_au/add_64 [35]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b30  (
    .i0(\exu/alu_au/add_64 [62]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b31  (
    .i0(\exu/alu_au/add_64 [63]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b4  (
    .i0(\exu/alu_au/add_64 [36]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b5  (
    .i0(\exu/alu_au/add_64 [37]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b6  (
    .i0(\exu/alu_au/add_64 [38]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b7  (
    .i0(\exu/alu_au/add_64 [39]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b8  (
    .i0(\exu/alu_au/add_64 [40]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux1_b9  (
    .i0(\exu/alu_au/add_64 [41]),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_add [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(81)
  binary_mux_s1_w1 \exu/alu_au/mux20_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [0]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [1]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [10]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [11]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [12]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [13]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [14]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [15]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [16]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [17]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [18]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [19]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [2]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [20]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [21]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [22]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [23]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [24]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [25]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [26]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [27]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [28]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [29]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [3]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [30]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [31]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [32]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [33]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [34]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [35]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [36]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [37]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [38]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [39]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [4]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [40]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [41]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [42]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [43]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [44]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [45]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [46]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [47]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [48]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [49]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [5]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [50]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [51]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [52]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [53]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [54]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [55]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [56]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [57]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [58]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [59]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [6]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [60]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [61]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [62]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [63]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [7]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [8]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux20_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_max [9]),
    .sel(mem_csr_data_max),
    .o(\exu/alu_au/n53 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  binary_mux_s1_w1 \exu/alu_au/mux21_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [0]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [1]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [10]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [11]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [12]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [13]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [14]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [15]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [16]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [17]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [18]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [19]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [2]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [20]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [21]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [22]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [23]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [24]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [25]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [26]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [27]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [28]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [29]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [3]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [30]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [31]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [32]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [33]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [34]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [35]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [36]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [37]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [38]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [39]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [4]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [40]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [41]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [42]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [43]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [44]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [45]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [46]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [47]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [48]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [49]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [5]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [50]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [51]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [52]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [53]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [54]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [55]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [56]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [57]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [58]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [59]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [6]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [60]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [61]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [62]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [63]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [7]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [8]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux21_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_min [9]),
    .sel(mem_csr_data_min),
    .o(\exu/alu_au/n55 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  binary_mux_s1_w1 \exu/alu_au/mux2_b0  (
    .i0(\exu/alu_au/add_64 [32]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b1  (
    .i0(\exu/alu_au/add_64 [33]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b10  (
    .i0(\exu/alu_au/add_64 [42]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b11  (
    .i0(\exu/alu_au/add_64 [43]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b12  (
    .i0(\exu/alu_au/add_64 [44]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b13  (
    .i0(\exu/alu_au/add_64 [45]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b14  (
    .i0(\exu/alu_au/add_64 [46]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b15  (
    .i0(\exu/alu_au/add_64 [47]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b16  (
    .i0(\exu/alu_au/add_64 [48]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b17  (
    .i0(\exu/alu_au/add_64 [49]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b18  (
    .i0(\exu/alu_au/add_64 [50]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b19  (
    .i0(\exu/alu_au/add_64 [51]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b2  (
    .i0(\exu/alu_au/add_64 [34]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b20  (
    .i0(\exu/alu_au/add_64 [52]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b21  (
    .i0(\exu/alu_au/add_64 [53]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b22  (
    .i0(\exu/alu_au/add_64 [54]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b23  (
    .i0(\exu/alu_au/add_64 [55]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b24  (
    .i0(\exu/alu_au/add_64 [56]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b25  (
    .i0(\exu/alu_au/add_64 [57]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b26  (
    .i0(\exu/alu_au/add_64 [58]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b27  (
    .i0(\exu/alu_au/add_64 [59]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b28  (
    .i0(\exu/alu_au/add_64 [60]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b29  (
    .i0(\exu/alu_au/add_64 [61]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b3  (
    .i0(\exu/alu_au/add_64 [35]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b30  (
    .i0(\exu/alu_au/add_64 [62]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b31  (
    .i0(\exu/alu_au/add_64 [63]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b4  (
    .i0(\exu/alu_au/add_64 [36]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b5  (
    .i0(\exu/alu_au/add_64 [37]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b6  (
    .i0(\exu/alu_au/add_64 [38]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b7  (
    .i0(\exu/alu_au/add_64 [39]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b8  (
    .i0(\exu/alu_au/add_64 [40]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux2_b9  (
    .i0(\exu/alu_au/add_64 [41]),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(ex_size[2]),
    .o(\exu/alu_au/alu_sub [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(84)
  binary_mux_s1_w1 \exu/alu_au/mux3_b0  (
    .i0(ds2[0]),
    .i1(\exu/alu_au/n16 [0]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b1  (
    .i0(ds2[1]),
    .i1(\exu/alu_au/n16 [1]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b10  (
    .i0(ds2[10]),
    .i1(\exu/alu_au/n16 [10]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b11  (
    .i0(ds2[11]),
    .i1(\exu/alu_au/n16 [11]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b12  (
    .i0(ds2[12]),
    .i1(\exu/alu_au/n16 [12]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b13  (
    .i0(ds2[13]),
    .i1(\exu/alu_au/n16 [13]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b14  (
    .i0(ds2[14]),
    .i1(\exu/alu_au/n16 [14]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b15  (
    .i0(ds2[15]),
    .i1(\exu/alu_au/n16 [15]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b16  (
    .i0(ds2[16]),
    .i1(\exu/alu_au/n16 [16]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b17  (
    .i0(ds2[17]),
    .i1(\exu/alu_au/n16 [17]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b18  (
    .i0(ds2[18]),
    .i1(\exu/alu_au/n16 [18]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b19  (
    .i0(ds2[19]),
    .i1(\exu/alu_au/n16 [19]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b2  (
    .i0(ds2[2]),
    .i1(\exu/alu_au/n16 [2]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b20  (
    .i0(ds2[20]),
    .i1(\exu/alu_au/n16 [20]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b21  (
    .i0(ds2[21]),
    .i1(\exu/alu_au/n16 [21]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b22  (
    .i0(ds2[22]),
    .i1(\exu/alu_au/n16 [22]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b23  (
    .i0(ds2[23]),
    .i1(\exu/alu_au/n16 [23]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b24  (
    .i0(ds2[24]),
    .i1(\exu/alu_au/n16 [24]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b25  (
    .i0(ds2[25]),
    .i1(\exu/alu_au/n16 [25]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b26  (
    .i0(ds2[26]),
    .i1(\exu/alu_au/n16 [26]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b27  (
    .i0(ds2[27]),
    .i1(\exu/alu_au/n16 [27]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b28  (
    .i0(ds2[28]),
    .i1(\exu/alu_au/n16 [28]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b29  (
    .i0(ds2[29]),
    .i1(\exu/alu_au/n16 [29]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b3  (
    .i0(ds2[3]),
    .i1(\exu/alu_au/n16 [3]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b30  (
    .i0(ds2[30]),
    .i1(\exu/alu_au/n16 [30]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b31  (
    .i0(ds2[31]),
    .i1(\exu/alu_au/n16 [31]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b32  (
    .i0(ds2[32]),
    .i1(\exu/alu_au/n16 [32]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b33  (
    .i0(ds2[33]),
    .i1(\exu/alu_au/n16 [33]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b34  (
    .i0(ds2[34]),
    .i1(\exu/alu_au/n16 [34]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b35  (
    .i0(ds2[35]),
    .i1(\exu/alu_au/n16 [35]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b36  (
    .i0(ds2[36]),
    .i1(\exu/alu_au/n16 [36]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b37  (
    .i0(ds2[37]),
    .i1(\exu/alu_au/n16 [37]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b38  (
    .i0(ds2[38]),
    .i1(\exu/alu_au/n16 [38]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b39  (
    .i0(ds2[39]),
    .i1(\exu/alu_au/n16 [39]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b4  (
    .i0(ds2[4]),
    .i1(\exu/alu_au/n16 [4]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b40  (
    .i0(ds2[40]),
    .i1(\exu/alu_au/n16 [40]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b41  (
    .i0(ds2[41]),
    .i1(\exu/alu_au/n16 [41]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b42  (
    .i0(ds2[42]),
    .i1(\exu/alu_au/n16 [42]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b43  (
    .i0(ds2[43]),
    .i1(\exu/alu_au/n16 [43]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b44  (
    .i0(ds2[44]),
    .i1(\exu/alu_au/n16 [44]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b45  (
    .i0(ds2[45]),
    .i1(\exu/alu_au/n16 [45]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b46  (
    .i0(ds2[46]),
    .i1(\exu/alu_au/n16 [46]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b47  (
    .i0(ds2[47]),
    .i1(\exu/alu_au/n16 [47]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b48  (
    .i0(ds2[48]),
    .i1(\exu/alu_au/n16 [48]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b49  (
    .i0(ds2[49]),
    .i1(\exu/alu_au/n16 [49]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b5  (
    .i0(ds2[5]),
    .i1(\exu/alu_au/n16 [5]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b50  (
    .i0(ds2[50]),
    .i1(\exu/alu_au/n16 [50]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b51  (
    .i0(ds2[51]),
    .i1(\exu/alu_au/n16 [51]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b52  (
    .i0(ds2[52]),
    .i1(\exu/alu_au/n16 [52]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b53  (
    .i0(ds2[53]),
    .i1(\exu/alu_au/n16 [53]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b54  (
    .i0(ds2[54]),
    .i1(\exu/alu_au/n16 [54]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b55  (
    .i0(ds2[55]),
    .i1(\exu/alu_au/n16 [55]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b56  (
    .i0(ds2[56]),
    .i1(\exu/alu_au/n16 [56]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b57  (
    .i0(ds2[57]),
    .i1(\exu/alu_au/n16 [57]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b58  (
    .i0(ds2[58]),
    .i1(\exu/alu_au/n16 [58]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b59  (
    .i0(ds2[59]),
    .i1(\exu/alu_au/n16 [59]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b6  (
    .i0(ds2[6]),
    .i1(\exu/alu_au/n16 [6]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b60  (
    .i0(ds2[60]),
    .i1(\exu/alu_au/n16 [60]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b61  (
    .i0(ds2[61]),
    .i1(\exu/alu_au/n16 [61]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b62  (
    .i0(ds2[62]),
    .i1(\exu/alu_au/n16 [62]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b63  (
    .i0(ds2[63]),
    .i1(\exu/alu_au/n16 [63]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b7  (
    .i0(ds2[7]),
    .i1(\exu/alu_au/n16 [7]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b8  (
    .i0(ds2[8]),
    .i1(\exu/alu_au/n16 [8]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux3_b9  (
    .i0(ds2[9]),
    .i1(\exu/alu_au/n16 [9]),
    .sel(and_clr),
    .o(\exu/alu_au/n18 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  binary_mux_s1_w1 \exu/alu_au/mux4_b0  (
    .i0(ds2[0]),
    .i1(ds1[0]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b1  (
    .i0(ds2[1]),
    .i1(ds1[1]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b10  (
    .i0(ds2[10]),
    .i1(ds1[10]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b11  (
    .i0(ds2[11]),
    .i1(ds1[11]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b12  (
    .i0(ds2[12]),
    .i1(ds1[12]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b13  (
    .i0(ds2[13]),
    .i1(ds1[13]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b14  (
    .i0(ds2[14]),
    .i1(ds1[14]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b15  (
    .i0(ds2[15]),
    .i1(ds1[15]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b16  (
    .i0(ds2[16]),
    .i1(ds1[16]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b17  (
    .i0(ds2[17]),
    .i1(ds1[17]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b18  (
    .i0(ds2[18]),
    .i1(ds1[18]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b19  (
    .i0(ds2[19]),
    .i1(ds1[19]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b2  (
    .i0(ds2[2]),
    .i1(ds1[2]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b20  (
    .i0(ds2[20]),
    .i1(ds1[20]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b21  (
    .i0(ds2[21]),
    .i1(ds1[21]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b22  (
    .i0(ds2[22]),
    .i1(ds1[22]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b23  (
    .i0(ds2[23]),
    .i1(ds1[23]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b24  (
    .i0(ds2[24]),
    .i1(ds1[24]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b25  (
    .i0(ds2[25]),
    .i1(ds1[25]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b26  (
    .i0(ds2[26]),
    .i1(ds1[26]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b27  (
    .i0(ds2[27]),
    .i1(ds1[27]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b28  (
    .i0(ds2[28]),
    .i1(ds1[28]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b29  (
    .i0(ds2[29]),
    .i1(ds1[29]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b3  (
    .i0(ds2[3]),
    .i1(ds1[3]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b30  (
    .i0(ds2[30]),
    .i1(ds1[30]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b31  (
    .i0(ds2[31]),
    .i1(ds1[31]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b32  (
    .i0(ds2[32]),
    .i1(ds1[32]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b33  (
    .i0(ds2[33]),
    .i1(ds1[33]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b34  (
    .i0(ds2[34]),
    .i1(ds1[34]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b35  (
    .i0(ds2[35]),
    .i1(ds1[35]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b36  (
    .i0(ds2[36]),
    .i1(ds1[36]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b37  (
    .i0(ds2[37]),
    .i1(ds1[37]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b38  (
    .i0(ds2[38]),
    .i1(ds1[38]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b39  (
    .i0(ds2[39]),
    .i1(ds1[39]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b4  (
    .i0(ds2[4]),
    .i1(ds1[4]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b40  (
    .i0(ds2[40]),
    .i1(ds1[40]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b41  (
    .i0(ds2[41]),
    .i1(ds1[41]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b42  (
    .i0(ds2[42]),
    .i1(ds1[42]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b43  (
    .i0(ds2[43]),
    .i1(ds1[43]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b44  (
    .i0(ds2[44]),
    .i1(ds1[44]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b45  (
    .i0(ds2[45]),
    .i1(ds1[45]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b46  (
    .i0(ds2[46]),
    .i1(ds1[46]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b47  (
    .i0(ds2[47]),
    .i1(ds1[47]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b48  (
    .i0(ds2[48]),
    .i1(ds1[48]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b49  (
    .i0(ds2[49]),
    .i1(ds1[49]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b5  (
    .i0(ds2[5]),
    .i1(ds1[5]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b50  (
    .i0(ds2[50]),
    .i1(ds1[50]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b51  (
    .i0(ds2[51]),
    .i1(ds1[51]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b52  (
    .i0(ds2[52]),
    .i1(ds1[52]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b53  (
    .i0(ds2[53]),
    .i1(ds1[53]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b54  (
    .i0(ds2[54]),
    .i1(ds1[54]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b55  (
    .i0(ds2[55]),
    .i1(ds1[55]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b56  (
    .i0(ds2[56]),
    .i1(ds1[56]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b57  (
    .i0(ds2[57]),
    .i1(ds1[57]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b58  (
    .i0(ds2[58]),
    .i1(ds1[58]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b59  (
    .i0(ds2[59]),
    .i1(ds1[59]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b6  (
    .i0(ds2[6]),
    .i1(ds1[6]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b60  (
    .i0(ds2[60]),
    .i1(ds1[60]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b61  (
    .i0(ds2[61]),
    .i1(ds1[61]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b62  (
    .i0(ds2[62]),
    .i1(ds1[62]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b63  (
    .i0(ds2[63]),
    .i1(ds1[63]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b7  (
    .i0(ds2[7]),
    .i1(ds1[7]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b8  (
    .i0(ds2[8]),
    .i1(ds1[8]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux4_b9  (
    .i0(ds2[9]),
    .i1(ds1[9]),
    .sel(\exu/alu_au/ds1_great_than_ds2 ),
    .o(\exu/alu_au/alu_max [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(95)
  binary_mux_s1_w1 \exu/alu_au/mux5_b0  (
    .i0(ds2[0]),
    .i1(ds1[0]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b1  (
    .i0(ds2[1]),
    .i1(ds1[1]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b10  (
    .i0(ds2[10]),
    .i1(ds1[10]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b11  (
    .i0(ds2[11]),
    .i1(ds1[11]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b12  (
    .i0(ds2[12]),
    .i1(ds1[12]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b13  (
    .i0(ds2[13]),
    .i1(ds1[13]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b14  (
    .i0(ds2[14]),
    .i1(ds1[14]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b15  (
    .i0(ds2[15]),
    .i1(ds1[15]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b16  (
    .i0(ds2[16]),
    .i1(ds1[16]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b17  (
    .i0(ds2[17]),
    .i1(ds1[17]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b18  (
    .i0(ds2[18]),
    .i1(ds1[18]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b19  (
    .i0(ds2[19]),
    .i1(ds1[19]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b2  (
    .i0(ds2[2]),
    .i1(ds1[2]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b20  (
    .i0(ds2[20]),
    .i1(ds1[20]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b21  (
    .i0(ds2[21]),
    .i1(ds1[21]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b22  (
    .i0(ds2[22]),
    .i1(ds1[22]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b23  (
    .i0(ds2[23]),
    .i1(ds1[23]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b24  (
    .i0(ds2[24]),
    .i1(ds1[24]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b25  (
    .i0(ds2[25]),
    .i1(ds1[25]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b26  (
    .i0(ds2[26]),
    .i1(ds1[26]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b27  (
    .i0(ds2[27]),
    .i1(ds1[27]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b28  (
    .i0(ds2[28]),
    .i1(ds1[28]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b29  (
    .i0(ds2[29]),
    .i1(ds1[29]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b3  (
    .i0(ds2[3]),
    .i1(ds1[3]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b30  (
    .i0(ds2[30]),
    .i1(ds1[30]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b31  (
    .i0(ds2[31]),
    .i1(ds1[31]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b32  (
    .i0(ds2[32]),
    .i1(ds1[32]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b33  (
    .i0(ds2[33]),
    .i1(ds1[33]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b34  (
    .i0(ds2[34]),
    .i1(ds1[34]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b35  (
    .i0(ds2[35]),
    .i1(ds1[35]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b36  (
    .i0(ds2[36]),
    .i1(ds1[36]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b37  (
    .i0(ds2[37]),
    .i1(ds1[37]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b38  (
    .i0(ds2[38]),
    .i1(ds1[38]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b39  (
    .i0(ds2[39]),
    .i1(ds1[39]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b4  (
    .i0(ds2[4]),
    .i1(ds1[4]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b40  (
    .i0(ds2[40]),
    .i1(ds1[40]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b41  (
    .i0(ds2[41]),
    .i1(ds1[41]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b42  (
    .i0(ds2[42]),
    .i1(ds1[42]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b43  (
    .i0(ds2[43]),
    .i1(ds1[43]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b44  (
    .i0(ds2[44]),
    .i1(ds1[44]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b45  (
    .i0(ds2[45]),
    .i1(ds1[45]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b46  (
    .i0(ds2[46]),
    .i1(ds1[46]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b47  (
    .i0(ds2[47]),
    .i1(ds1[47]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b48  (
    .i0(ds2[48]),
    .i1(ds1[48]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b49  (
    .i0(ds2[49]),
    .i1(ds1[49]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b5  (
    .i0(ds2[5]),
    .i1(ds1[5]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b50  (
    .i0(ds2[50]),
    .i1(ds1[50]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b51  (
    .i0(ds2[51]),
    .i1(ds1[51]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b52  (
    .i0(ds2[52]),
    .i1(ds1[52]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b53  (
    .i0(ds2[53]),
    .i1(ds1[53]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b54  (
    .i0(ds2[54]),
    .i1(ds1[54]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b55  (
    .i0(ds2[55]),
    .i1(ds1[55]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b56  (
    .i0(ds2[56]),
    .i1(ds1[56]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b57  (
    .i0(ds2[57]),
    .i1(ds1[57]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b58  (
    .i0(ds2[58]),
    .i1(ds1[58]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b59  (
    .i0(ds2[59]),
    .i1(ds1[59]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b6  (
    .i0(ds2[6]),
    .i1(ds1[6]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b60  (
    .i0(ds2[60]),
    .i1(ds1[60]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b61  (
    .i0(ds2[61]),
    .i1(ds1[61]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b62  (
    .i0(ds2[62]),
    .i1(ds1[62]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b63  (
    .i0(ds2[63]),
    .i1(ds1[63]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b7  (
    .i0(ds2[7]),
    .i1(ds1[7]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b8  (
    .i0(ds2[8]),
    .i1(ds1[8]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux5_b9  (
    .i0(ds2[9]),
    .i1(ds1[9]),
    .sel(\exu/alu_au/ds1_light_than_ds2 ),
    .o(\exu/alu_au/alu_min [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(96)
  binary_mux_s1_w1 \exu/alu_au/mux6_b0  (
    .i0(1'b0),
    .i1(ds1[0]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b1  (
    .i0(1'b0),
    .i1(ds1[1]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b10  (
    .i0(1'b0),
    .i1(ds1[10]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b11  (
    .i0(1'b0),
    .i1(ds1[11]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b12  (
    .i0(1'b0),
    .i1(ds1[12]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b13  (
    .i0(1'b0),
    .i1(ds1[13]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b14  (
    .i0(1'b0),
    .i1(ds1[14]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b15  (
    .i0(1'b0),
    .i1(ds1[15]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b16  (
    .i0(1'b0),
    .i1(ds1[16]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b17  (
    .i0(1'b0),
    .i1(ds1[17]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b18  (
    .i0(1'b0),
    .i1(ds1[18]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b19  (
    .i0(1'b0),
    .i1(ds1[19]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b2  (
    .i0(1'b0),
    .i1(ds1[2]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b20  (
    .i0(1'b0),
    .i1(ds1[20]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b21  (
    .i0(1'b0),
    .i1(ds1[21]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b22  (
    .i0(1'b0),
    .i1(ds1[22]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b23  (
    .i0(1'b0),
    .i1(ds1[23]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b24  (
    .i0(1'b0),
    .i1(ds1[24]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b25  (
    .i0(1'b0),
    .i1(ds1[25]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b26  (
    .i0(1'b0),
    .i1(ds1[26]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b27  (
    .i0(1'b0),
    .i1(ds1[27]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b28  (
    .i0(1'b0),
    .i1(ds1[28]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b29  (
    .i0(1'b0),
    .i1(ds1[29]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b3  (
    .i0(1'b0),
    .i1(ds1[3]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b30  (
    .i0(1'b0),
    .i1(ds1[30]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b31  (
    .i0(1'b0),
    .i1(ds1[31]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b32  (
    .i0(1'b0),
    .i1(ds1[32]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b33  (
    .i0(1'b0),
    .i1(ds1[33]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b34  (
    .i0(1'b0),
    .i1(ds1[34]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b35  (
    .i0(1'b0),
    .i1(ds1[35]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b36  (
    .i0(1'b0),
    .i1(ds1[36]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b37  (
    .i0(1'b0),
    .i1(ds1[37]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b38  (
    .i0(1'b0),
    .i1(ds1[38]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b39  (
    .i0(1'b0),
    .i1(ds1[39]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b4  (
    .i0(1'b0),
    .i1(ds1[4]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b40  (
    .i0(1'b0),
    .i1(ds1[40]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b41  (
    .i0(1'b0),
    .i1(ds1[41]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b42  (
    .i0(1'b0),
    .i1(ds1[42]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b43  (
    .i0(1'b0),
    .i1(ds1[43]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b44  (
    .i0(1'b0),
    .i1(ds1[44]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b45  (
    .i0(1'b0),
    .i1(ds1[45]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b46  (
    .i0(1'b0),
    .i1(ds1[46]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b47  (
    .i0(1'b0),
    .i1(ds1[47]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b48  (
    .i0(1'b0),
    .i1(ds1[48]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b49  (
    .i0(1'b0),
    .i1(ds1[49]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b5  (
    .i0(1'b0),
    .i1(ds1[5]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b50  (
    .i0(1'b0),
    .i1(ds1[50]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b51  (
    .i0(1'b0),
    .i1(ds1[51]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b52  (
    .i0(1'b0),
    .i1(ds1[52]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b53  (
    .i0(1'b0),
    .i1(ds1[53]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b54  (
    .i0(1'b0),
    .i1(ds1[54]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b55  (
    .i0(1'b0),
    .i1(ds1[55]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b56  (
    .i0(1'b0),
    .i1(ds1[56]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b57  (
    .i0(1'b0),
    .i1(ds1[57]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b58  (
    .i0(1'b0),
    .i1(ds1[58]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b59  (
    .i0(1'b0),
    .i1(ds1[59]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b6  (
    .i0(1'b0),
    .i1(ds1[6]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b60  (
    .i0(1'b0),
    .i1(ds1[60]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b61  (
    .i0(1'b0),
    .i1(ds1[61]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b62  (
    .i0(1'b0),
    .i1(ds1[62]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b63  (
    .i0(1'b0),
    .i1(ds1[63]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b7  (
    .i0(1'b0),
    .i1(ds1[7]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b8  (
    .i0(1'b0),
    .i1(ds1[8]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux6_b9  (
    .i0(1'b0),
    .i1(ds1[9]),
    .sel(rd_data_ds1),
    .o(\exu/alu_au/n28 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(99)
  binary_mux_s1_w1 \exu/alu_au/mux7_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [0]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [1]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [10]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [11]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [12]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [13]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [14]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [15]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [16]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [17]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [18]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [19]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [2]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [20]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [21]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [22]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [23]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [24]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [25]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [26]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [27]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [28]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [29]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [3]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [30]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [31]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [32]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [33]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [34]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [35]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [36]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [37]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [38]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [39]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [4]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [40]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [41]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [42]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [43]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [44]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [45]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [46]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [47]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [48]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [49]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [5]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [50]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [51]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [52]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [53]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [54]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [55]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [56]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [57]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [58]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [59]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [6]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [60]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [61]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [62]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_add [63]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [7]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [8]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux7_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/add_64 [9]),
    .sel(rd_data_add),
    .o(\exu/alu_au/n29 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  binary_mux_s1_w1 \exu/alu_au/mux8_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [0]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [1]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [10]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [11]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [12]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [13]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [14]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [15]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [16]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [17]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [18]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [19]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [2]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [20]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [21]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [22]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [23]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [24]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [25]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [26]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [27]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [28]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [29]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [3]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [30]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [31]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [32]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [33]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [34]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [35]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [36]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [37]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [38]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [39]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [4]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [40]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [41]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [42]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [43]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [44]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [45]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [46]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [47]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [48]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [49]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [5]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [50]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [51]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [52]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [53]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [54]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [55]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [56]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [57]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [58]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [59]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [6]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [60]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [61]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [62]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_sub [63]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [7]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [8]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux8_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/sub_64 [9]),
    .sel(rd_data_sub),
    .o(\exu/alu_au/n31 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  binary_mux_s1_w1 \exu/alu_au/mux9_b0  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [0]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [0]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b1  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [1]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [1]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b10  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [10]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [10]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b11  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [11]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [11]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b12  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [12]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [12]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b13  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [13]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [13]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b14  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [14]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [14]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b15  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [15]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [15]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b16  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [16]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [16]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b17  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [17]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [17]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b18  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [18]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [18]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b19  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [19]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [19]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b2  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [2]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [2]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b20  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [20]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [20]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b21  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [21]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [21]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b22  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [22]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [22]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b23  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [23]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [23]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b24  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [24]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [24]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b25  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [25]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [25]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b26  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [26]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [26]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b27  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [27]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [27]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b28  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [28]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [28]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b29  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [29]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [29]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b3  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [3]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [3]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b30  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [30]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [30]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b31  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [31]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [31]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b32  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [32]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [32]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b33  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [33]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [33]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b34  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [34]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [34]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b35  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [35]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [35]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b36  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [36]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [36]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b37  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [37]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [37]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b38  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [38]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [38]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b39  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [39]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [39]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b4  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [4]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [4]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b40  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [40]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [40]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b41  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [41]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [41]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b42  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [42]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [42]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b43  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [43]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [43]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b44  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [44]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [44]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b45  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [45]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [45]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b46  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [46]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [46]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b47  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [47]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [47]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b48  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [48]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [48]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b49  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [49]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [49]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b5  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [5]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [5]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b50  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [50]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [50]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b51  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [51]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [51]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b52  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [52]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [52]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b53  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [53]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [53]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b54  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [54]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [54]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b55  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [55]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [55]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b56  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [56]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [56]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b57  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [57]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [57]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b58  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [58]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [58]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b59  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [59]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [59]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b6  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [6]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [6]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b60  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [60]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [60]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b61  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [61]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [61]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b62  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [62]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [62]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b63  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [63]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [63]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b7  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [7]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [7]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b8  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [8]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [8]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  binary_mux_s1_w1 \exu/alu_au/mux9_b9  (
    .i0(1'b0),
    .i1(\exu/alu_au/alu_and [9]),
    .sel(rd_data_and),
    .o(\exu/alu_au/n33 [9]));  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u10  (\exu/alu_au/n7 , \exu/alu_au/n2 , \exu/alu_au/n6 );  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(72)
  or \exu/alu_au/u100  (\exu/alu_data_mem_csr [51], \exu/alu_au/n54 [51], \exu/alu_au/n55 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u101  (\exu/alu_data_mem_csr [52], \exu/alu_au/n54 [52], \exu/alu_au/n55 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u102  (\exu/alu_data_mem_csr [53], \exu/alu_au/n54 [53], \exu/alu_au/n55 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u103  (\exu/alu_data_mem_csr [54], \exu/alu_au/n54 [54], \exu/alu_au/n55 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u104  (\exu/alu_data_mem_csr [55], \exu/alu_au/n54 [55], \exu/alu_au/n55 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u105  (\exu/alu_data_mem_csr [56], \exu/alu_au/n54 [56], \exu/alu_au/n55 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  xor \exu/alu_au/u1058  (\exu/alu_au/alu_xor [1], ds1[1], ds2[1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1059  (\exu/alu_au/alu_xor [2], ds1[2], ds2[2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  or \exu/alu_au/u106  (\exu/alu_data_mem_csr [57], \exu/alu_au/n54 [57], \exu/alu_au/n55 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  xor \exu/alu_au/u1060  (\exu/alu_au/alu_xor [3], ds1[3], ds2[3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1061  (\exu/alu_au/alu_xor [4], ds1[4], ds2[4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1062  (\exu/alu_au/alu_xor [5], ds1[5], ds2[5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1063  (\exu/alu_au/alu_xor [6], ds1[6], ds2[6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1064  (\exu/alu_au/alu_xor [7], ds1[7], ds2[7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1065  (\exu/alu_au/alu_xor [8], ds1[8], ds2[8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1066  (\exu/alu_au/alu_xor [9], ds1[9], ds2[9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1067  (\exu/alu_au/alu_xor [10], ds1[10], ds2[10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1068  (\exu/alu_au/alu_xor [11], ds1[11], ds2[11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1069  (\exu/alu_au/alu_xor [12], ds1[12], ds2[12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  or \exu/alu_au/u107  (\exu/alu_data_mem_csr [58], \exu/alu_au/n54 [58], \exu/alu_au/n55 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  xor \exu/alu_au/u1070  (\exu/alu_au/alu_xor [13], ds1[13], ds2[13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1071  (\exu/alu_au/alu_xor [14], ds1[14], ds2[14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1072  (\exu/alu_au/alu_xor [15], ds1[15], ds2[15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1073  (\exu/alu_au/alu_xor [16], ds1[16], ds2[16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1074  (\exu/alu_au/alu_xor [17], ds1[17], ds2[17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1075  (\exu/alu_au/alu_xor [18], ds1[18], ds2[18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1076  (\exu/alu_au/alu_xor [19], ds1[19], ds2[19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1077  (\exu/alu_au/alu_xor [20], ds1[20], ds2[20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1078  (\exu/alu_au/alu_xor [21], ds1[21], ds2[21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1079  (\exu/alu_au/alu_xor [22], ds1[22], ds2[22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  or \exu/alu_au/u108  (\exu/alu_data_mem_csr [59], \exu/alu_au/n54 [59], \exu/alu_au/n55 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  xor \exu/alu_au/u1080  (\exu/alu_au/alu_xor [23], ds1[23], ds2[23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1081  (\exu/alu_au/alu_xor [24], ds1[24], ds2[24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1082  (\exu/alu_au/alu_xor [25], ds1[25], ds2[25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1083  (\exu/alu_au/alu_xor [26], ds1[26], ds2[26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1084  (\exu/alu_au/alu_xor [27], ds1[27], ds2[27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1085  (\exu/alu_au/alu_xor [28], ds1[28], ds2[28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1086  (\exu/alu_au/alu_xor [29], ds1[29], ds2[29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1087  (\exu/alu_au/alu_xor [30], ds1[30], ds2[30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1088  (\exu/alu_au/alu_xor [31], ds1[31], ds2[31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1089  (\exu/alu_au/alu_xor [32], ds1[32], ds2[32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  or \exu/alu_au/u109  (\exu/alu_data_mem_csr [60], \exu/alu_au/n54 [60], \exu/alu_au/n55 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  xor \exu/alu_au/u1090  (\exu/alu_au/alu_xor [33], ds1[33], ds2[33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1091  (\exu/alu_au/alu_xor [34], ds1[34], ds2[34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1092  (\exu/alu_au/alu_xor [35], ds1[35], ds2[35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1093  (\exu/alu_au/alu_xor [36], ds1[36], ds2[36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1094  (\exu/alu_au/alu_xor [37], ds1[37], ds2[37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1095  (\exu/alu_au/alu_xor [38], ds1[38], ds2[38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1096  (\exu/alu_au/alu_xor [39], ds1[39], ds2[39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1097  (\exu/alu_au/alu_xor [40], ds1[40], ds2[40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1098  (\exu/alu_au/alu_xor [41], ds1[41], ds2[41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1099  (\exu/alu_au/alu_xor [42], ds1[42], ds2[42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  and \exu/alu_au/u11  (\exu/alu_au/n8 , \exu/alu_au/n0 , \exu/alu_au/n7 );  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(72)
  or \exu/alu_au/u110  (\exu/alu_data_mem_csr [61], \exu/alu_au/n54 [61], \exu/alu_au/n55 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  xor \exu/alu_au/u1100  (\exu/alu_au/alu_xor [43], ds1[43], ds2[43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1101  (\exu/alu_au/alu_xor [44], ds1[44], ds2[44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1102  (\exu/alu_au/alu_xor [45], ds1[45], ds2[45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1103  (\exu/alu_au/alu_xor [46], ds1[46], ds2[46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1104  (\exu/alu_au/alu_xor [47], ds1[47], ds2[47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1105  (\exu/alu_au/alu_xor [48], ds1[48], ds2[48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1106  (\exu/alu_au/alu_xor [49], ds1[49], ds2[49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1107  (\exu/alu_au/alu_xor [50], ds1[50], ds2[50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1108  (\exu/alu_au/alu_xor [51], ds1[51], ds2[51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1109  (\exu/alu_au/alu_xor [52], ds1[52], ds2[52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  or \exu/alu_au/u111  (\exu/alu_data_mem_csr [62], \exu/alu_au/n54 [62], \exu/alu_au/n55 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  xor \exu/alu_au/u1110  (\exu/alu_au/alu_xor [53], ds1[53], ds2[53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1111  (\exu/alu_au/alu_xor [54], ds1[54], ds2[54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1112  (\exu/alu_au/alu_xor [55], ds1[55], ds2[55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1113  (\exu/alu_au/alu_xor [56], ds1[56], ds2[56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1114  (\exu/alu_au/alu_xor [57], ds1[57], ds2[57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1115  (\exu/alu_au/alu_xor [58], ds1[58], ds2[58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1116  (\exu/alu_au/alu_xor [59], ds1[59], ds2[59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1117  (\exu/alu_au/alu_xor [60], ds1[60], ds2[60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1118  (\exu/alu_au/alu_xor [61], ds1[61], ds2[61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  xor \exu/alu_au/u1119  (\exu/alu_au/alu_xor [62], ds1[62], ds2[62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  or \exu/alu_au/u112  (\exu/alu_data_mem_csr [63], \exu/alu_au/n54 [63], \exu/alu_au/n55 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  xor \exu/alu_au/u1120  (\exu/alu_au/alu_xor [63], ds1[63], ds2[63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  or \exu/alu_au/u1121  (\exu/alu_au/alu_or [1], ds1[1], ds2[1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1122  (\exu/alu_au/alu_or [2], ds1[2], ds2[2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1123  (\exu/alu_au/alu_or [3], ds1[3], ds2[3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1124  (\exu/alu_au/alu_or [4], ds1[4], ds2[4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1125  (\exu/alu_au/alu_or [5], ds1[5], ds2[5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1126  (\exu/alu_au/alu_or [6], ds1[6], ds2[6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1127  (\exu/alu_au/alu_or [7], ds1[7], ds2[7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1128  (\exu/alu_au/alu_or [8], ds1[8], ds2[8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1129  (\exu/alu_au/alu_or [9], ds1[9], ds2[9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u113  (\exu/alu_au/n54 [1], \exu/alu_au/n52 [1], \exu/alu_au/n53 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u1130  (\exu/alu_au/alu_or [10], ds1[10], ds2[10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1131  (\exu/alu_au/alu_or [11], ds1[11], ds2[11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1132  (\exu/alu_au/alu_or [12], ds1[12], ds2[12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1133  (\exu/alu_au/alu_or [13], ds1[13], ds2[13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1134  (\exu/alu_au/alu_or [14], ds1[14], ds2[14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1135  (\exu/alu_au/alu_or [15], ds1[15], ds2[15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1136  (\exu/alu_au/alu_or [16], ds1[16], ds2[16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1137  (\exu/alu_au/alu_or [17], ds1[17], ds2[17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1138  (\exu/alu_au/alu_or [18], ds1[18], ds2[18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1139  (\exu/alu_au/alu_or [19], ds1[19], ds2[19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u114  (\exu/alu_au/n54 [2], \exu/alu_au/n52 [2], \exu/alu_au/n53 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u1140  (\exu/alu_au/alu_or [20], ds1[20], ds2[20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1141  (\exu/alu_au/alu_or [21], ds1[21], ds2[21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1142  (\exu/alu_au/alu_or [22], ds1[22], ds2[22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1143  (\exu/alu_au/alu_or [23], ds1[23], ds2[23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1144  (\exu/alu_au/alu_or [24], ds1[24], ds2[24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1145  (\exu/alu_au/alu_or [25], ds1[25], ds2[25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1146  (\exu/alu_au/alu_or [26], ds1[26], ds2[26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1147  (\exu/alu_au/alu_or [27], ds1[27], ds2[27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1148  (\exu/alu_au/alu_or [28], ds1[28], ds2[28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1149  (\exu/alu_au/alu_or [29], ds1[29], ds2[29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u115  (\exu/alu_au/n54 [3], \exu/alu_au/n52 [3], \exu/alu_au/n53 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u1150  (\exu/alu_au/alu_or [30], ds1[30], ds2[30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1151  (\exu/alu_au/alu_or [31], ds1[31], ds2[31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1152  (\exu/alu_au/alu_or [32], ds1[32], ds2[32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1153  (\exu/alu_au/alu_or [33], ds1[33], ds2[33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1154  (\exu/alu_au/alu_or [34], ds1[34], ds2[34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1155  (\exu/alu_au/alu_or [35], ds1[35], ds2[35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1156  (\exu/alu_au/alu_or [36], ds1[36], ds2[36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1157  (\exu/alu_au/alu_or [37], ds1[37], ds2[37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1158  (\exu/alu_au/alu_or [38], ds1[38], ds2[38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1159  (\exu/alu_au/alu_or [39], ds1[39], ds2[39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u116  (\exu/alu_au/n54 [4], \exu/alu_au/n52 [4], \exu/alu_au/n53 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u1160  (\exu/alu_au/alu_or [40], ds1[40], ds2[40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1161  (\exu/alu_au/alu_or [41], ds1[41], ds2[41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1162  (\exu/alu_au/alu_or [42], ds1[42], ds2[42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1163  (\exu/alu_au/alu_or [43], ds1[43], ds2[43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1164  (\exu/alu_au/alu_or [44], ds1[44], ds2[44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1165  (\exu/alu_au/alu_or [45], ds1[45], ds2[45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1166  (\exu/alu_au/alu_or [46], ds1[46], ds2[46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1167  (\exu/alu_au/alu_or [47], ds1[47], ds2[47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1168  (\exu/alu_au/alu_or [48], ds1[48], ds2[48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1169  (\exu/alu_au/alu_or [49], ds1[49], ds2[49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u117  (\exu/alu_au/n54 [5], \exu/alu_au/n52 [5], \exu/alu_au/n53 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u1170  (\exu/alu_au/alu_or [50], ds1[50], ds2[50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1171  (\exu/alu_au/alu_or [51], ds1[51], ds2[51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1172  (\exu/alu_au/alu_or [52], ds1[52], ds2[52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1173  (\exu/alu_au/alu_or [53], ds1[53], ds2[53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1174  (\exu/alu_au/alu_or [54], ds1[54], ds2[54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1175  (\exu/alu_au/alu_or [55], ds1[55], ds2[55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1176  (\exu/alu_au/alu_or [56], ds1[56], ds2[56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1177  (\exu/alu_au/alu_or [57], ds1[57], ds2[57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1178  (\exu/alu_au/alu_or [58], ds1[58], ds2[58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1179  (\exu/alu_au/alu_or [59], ds1[59], ds2[59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u118  (\exu/alu_au/n54 [6], \exu/alu_au/n52 [6], \exu/alu_au/n53 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u1180  (\exu/alu_au/alu_or [60], ds1[60], ds2[60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1181  (\exu/alu_au/alu_or [61], ds1[61], ds2[61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1182  (\exu/alu_au/alu_or [62], ds1[62], ds2[62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u1183  (\exu/alu_au/alu_or [63], ds1[63], ds2[63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  and \exu/alu_au/u1184  (\exu/alu_au/alu_and [1], ds1[1], \exu/alu_au/n18 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1185  (\exu/alu_au/alu_and [2], ds1[2], \exu/alu_au/n18 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1186  (\exu/alu_au/alu_and [3], ds1[3], \exu/alu_au/n18 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1187  (\exu/alu_au/alu_and [4], ds1[4], \exu/alu_au/n18 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1188  (\exu/alu_au/alu_and [5], ds1[5], \exu/alu_au/n18 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1189  (\exu/alu_au/alu_and [6], ds1[6], \exu/alu_au/n18 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  or \exu/alu_au/u119  (\exu/alu_au/n54 [7], \exu/alu_au/n52 [7], \exu/alu_au/n53 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  and \exu/alu_au/u1190  (\exu/alu_au/alu_and [7], ds1[7], \exu/alu_au/n18 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1191  (\exu/alu_au/alu_and [8], ds1[8], \exu/alu_au/n18 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1192  (\exu/alu_au/alu_and [9], ds1[9], \exu/alu_au/n18 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1193  (\exu/alu_au/alu_and [10], ds1[10], \exu/alu_au/n18 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1194  (\exu/alu_au/alu_and [11], ds1[11], \exu/alu_au/n18 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1195  (\exu/alu_au/alu_and [12], ds1[12], \exu/alu_au/n18 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1196  (\exu/alu_au/alu_and [13], ds1[13], \exu/alu_au/n18 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1197  (\exu/alu_au/alu_and [14], ds1[14], \exu/alu_au/n18 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1198  (\exu/alu_au/alu_and [15], ds1[15], \exu/alu_au/n18 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1199  (\exu/alu_au/alu_and [16], ds1[16], \exu/alu_au/n18 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  or \exu/alu_au/u12  (\exu/alu_data_mem_csr [6], \exu/alu_au/n54 [6], \exu/alu_au/n55 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u120  (\exu/alu_au/n54 [8], \exu/alu_au/n52 [8], \exu/alu_au/n53 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  and \exu/alu_au/u1200  (\exu/alu_au/alu_and [17], ds1[17], \exu/alu_au/n18 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1201  (\exu/alu_au/alu_and [18], ds1[18], \exu/alu_au/n18 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1202  (\exu/alu_au/alu_and [19], ds1[19], \exu/alu_au/n18 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1203  (\exu/alu_au/alu_and [20], ds1[20], \exu/alu_au/n18 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1204  (\exu/alu_au/alu_and [21], ds1[21], \exu/alu_au/n18 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1205  (\exu/alu_au/alu_and [22], ds1[22], \exu/alu_au/n18 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1206  (\exu/alu_au/alu_and [23], ds1[23], \exu/alu_au/n18 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1207  (\exu/alu_au/alu_and [24], ds1[24], \exu/alu_au/n18 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1208  (\exu/alu_au/alu_and [25], ds1[25], \exu/alu_au/n18 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1209  (\exu/alu_au/alu_and [26], ds1[26], \exu/alu_au/n18 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  or \exu/alu_au/u121  (\exu/alu_au/n54 [9], \exu/alu_au/n52 [9], \exu/alu_au/n53 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  and \exu/alu_au/u1210  (\exu/alu_au/alu_and [27], ds1[27], \exu/alu_au/n18 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1211  (\exu/alu_au/alu_and [28], ds1[28], \exu/alu_au/n18 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1212  (\exu/alu_au/alu_and [29], ds1[29], \exu/alu_au/n18 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1213  (\exu/alu_au/alu_and [30], ds1[30], \exu/alu_au/n18 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1214  (\exu/alu_au/alu_and [31], ds1[31], \exu/alu_au/n18 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1215  (\exu/alu_au/alu_and [32], ds1[32], \exu/alu_au/n18 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1216  (\exu/alu_au/alu_and [33], ds1[33], \exu/alu_au/n18 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1217  (\exu/alu_au/alu_and [34], ds1[34], \exu/alu_au/n18 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1218  (\exu/alu_au/alu_and [35], ds1[35], \exu/alu_au/n18 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1219  (\exu/alu_au/alu_and [36], ds1[36], \exu/alu_au/n18 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  or \exu/alu_au/u122  (\exu/alu_au/n54 [10], \exu/alu_au/n52 [10], \exu/alu_au/n53 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  and \exu/alu_au/u1220  (\exu/alu_au/alu_and [37], ds1[37], \exu/alu_au/n18 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1221  (\exu/alu_au/alu_and [38], ds1[38], \exu/alu_au/n18 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1222  (\exu/alu_au/alu_and [39], ds1[39], \exu/alu_au/n18 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1223  (\exu/alu_au/alu_and [40], ds1[40], \exu/alu_au/n18 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1224  (\exu/alu_au/alu_and [41], ds1[41], \exu/alu_au/n18 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1225  (\exu/alu_au/alu_and [42], ds1[42], \exu/alu_au/n18 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1226  (\exu/alu_au/alu_and [43], ds1[43], \exu/alu_au/n18 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1227  (\exu/alu_au/alu_and [44], ds1[44], \exu/alu_au/n18 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1228  (\exu/alu_au/alu_and [45], ds1[45], \exu/alu_au/n18 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1229  (\exu/alu_au/alu_and [46], ds1[46], \exu/alu_au/n18 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  or \exu/alu_au/u123  (\exu/alu_au/n54 [11], \exu/alu_au/n52 [11], \exu/alu_au/n53 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  and \exu/alu_au/u1230  (\exu/alu_au/alu_and [47], ds1[47], \exu/alu_au/n18 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1231  (\exu/alu_au/alu_and [48], ds1[48], \exu/alu_au/n18 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1232  (\exu/alu_au/alu_and [49], ds1[49], \exu/alu_au/n18 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1233  (\exu/alu_au/alu_and [50], ds1[50], \exu/alu_au/n18 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1234  (\exu/alu_au/alu_and [51], ds1[51], \exu/alu_au/n18 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1235  (\exu/alu_au/alu_and [52], ds1[52], \exu/alu_au/n18 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1236  (\exu/alu_au/alu_and [53], ds1[53], \exu/alu_au/n18 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1237  (\exu/alu_au/alu_and [54], ds1[54], \exu/alu_au/n18 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1238  (\exu/alu_au/alu_and [55], ds1[55], \exu/alu_au/n18 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1239  (\exu/alu_au/alu_and [56], ds1[56], \exu/alu_au/n18 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  or \exu/alu_au/u124  (\exu/alu_au/n54 [12], \exu/alu_au/n52 [12], \exu/alu_au/n53 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  and \exu/alu_au/u1240  (\exu/alu_au/alu_and [57], ds1[57], \exu/alu_au/n18 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1241  (\exu/alu_au/alu_and [58], ds1[58], \exu/alu_au/n18 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1242  (\exu/alu_au/alu_and [59], ds1[59], \exu/alu_au/n18 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1243  (\exu/alu_au/alu_and [60], ds1[60], \exu/alu_au/n18 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1244  (\exu/alu_au/alu_and [61], ds1[61], \exu/alu_au/n18 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1245  (\exu/alu_au/alu_and [62], ds1[62], \exu/alu_au/n18 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  and \exu/alu_au/u1246  (\exu/alu_au/alu_and [63], ds1[63], \exu/alu_au/n18 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  or \exu/alu_au/u125  (\exu/alu_au/n54 [13], \exu/alu_au/n52 [13], \exu/alu_au/n53 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u126  (\exu/alu_au/n54 [14], \exu/alu_au/n52 [14], \exu/alu_au/n53 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u127  (\exu/alu_au/n54 [15], \exu/alu_au/n52 [15], \exu/alu_au/n53 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u128  (\exu/alu_au/n54 [16], \exu/alu_au/n52 [16], \exu/alu_au/n53 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u129  (\exu/alu_au/n54 [17], \exu/alu_au/n52 [17], \exu/alu_au/n53 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  and \exu/alu_au/u13  (\exu/alu_au/n9 , unsign, \exu/alu_au/n5 );  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(73)
  or \exu/alu_au/u130  (\exu/alu_au/n54 [18], \exu/alu_au/n52 [18], \exu/alu_au/n53 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  not \exu/alu_au/u1309  (\exu/alu_au/n16 [1], ds2[1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  or \exu/alu_au/u131  (\exu/alu_au/n54 [19], \exu/alu_au/n52 [19], \exu/alu_au/n53 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  not \exu/alu_au/u1310  (\exu/alu_au/n16 [2], ds2[2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1311  (\exu/alu_au/n16 [3], ds2[3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1312  (\exu/alu_au/n16 [4], ds2[4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1313  (\exu/alu_au/n16 [5], ds2[5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1314  (\exu/alu_au/n16 [6], ds2[6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1315  (\exu/alu_au/n16 [7], ds2[7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1316  (\exu/alu_au/n16 [8], ds2[8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1317  (\exu/alu_au/n16 [9], ds2[9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1318  (\exu/alu_au/n16 [10], ds2[10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1319  (\exu/alu_au/n16 [11], ds2[11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  or \exu/alu_au/u132  (\exu/alu_au/n54 [20], \exu/alu_au/n52 [20], \exu/alu_au/n53 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  not \exu/alu_au/u1320  (\exu/alu_au/n16 [12], ds2[12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1321  (\exu/alu_au/n16 [13], ds2[13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1322  (\exu/alu_au/n16 [14], ds2[14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1323  (\exu/alu_au/n16 [15], ds2[15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1324  (\exu/alu_au/n16 [16], ds2[16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1325  (\exu/alu_au/n16 [17], ds2[17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1326  (\exu/alu_au/n16 [18], ds2[18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1327  (\exu/alu_au/n16 [19], ds2[19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1328  (\exu/alu_au/n16 [20], ds2[20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1329  (\exu/alu_au/n16 [21], ds2[21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  or \exu/alu_au/u133  (\exu/alu_au/n54 [21], \exu/alu_au/n52 [21], \exu/alu_au/n53 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  not \exu/alu_au/u1330  (\exu/alu_au/n16 [22], ds2[22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1331  (\exu/alu_au/n16 [23], ds2[23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1332  (\exu/alu_au/n16 [24], ds2[24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1333  (\exu/alu_au/n16 [25], ds2[25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1334  (\exu/alu_au/n16 [26], ds2[26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1335  (\exu/alu_au/n16 [27], ds2[27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1336  (\exu/alu_au/n16 [28], ds2[28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1337  (\exu/alu_au/n16 [29], ds2[29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1338  (\exu/alu_au/n16 [30], ds2[30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1339  (\exu/alu_au/n16 [31], ds2[31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  or \exu/alu_au/u134  (\exu/alu_au/n54 [22], \exu/alu_au/n52 [22], \exu/alu_au/n53 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  not \exu/alu_au/u1340  (\exu/alu_au/n16 [32], ds2[32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1341  (\exu/alu_au/n16 [33], ds2[33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1342  (\exu/alu_au/n16 [34], ds2[34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1343  (\exu/alu_au/n16 [35], ds2[35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1344  (\exu/alu_au/n16 [36], ds2[36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1345  (\exu/alu_au/n16 [37], ds2[37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1346  (\exu/alu_au/n16 [38], ds2[38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1347  (\exu/alu_au/n16 [39], ds2[39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1348  (\exu/alu_au/n16 [40], ds2[40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1349  (\exu/alu_au/n16 [41], ds2[41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  or \exu/alu_au/u135  (\exu/alu_au/n54 [23], \exu/alu_au/n52 [23], \exu/alu_au/n53 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  not \exu/alu_au/u1350  (\exu/alu_au/n16 [42], ds2[42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1351  (\exu/alu_au/n16 [43], ds2[43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1352  (\exu/alu_au/n16 [44], ds2[44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1353  (\exu/alu_au/n16 [45], ds2[45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1354  (\exu/alu_au/n16 [46], ds2[46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1355  (\exu/alu_au/n16 [47], ds2[47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1356  (\exu/alu_au/n16 [48], ds2[48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1357  (\exu/alu_au/n16 [49], ds2[49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1358  (\exu/alu_au/n16 [50], ds2[50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1359  (\exu/alu_au/n16 [51], ds2[51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  or \exu/alu_au/u136  (\exu/alu_au/n54 [24], \exu/alu_au/n52 [24], \exu/alu_au/n53 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  not \exu/alu_au/u1360  (\exu/alu_au/n16 [52], ds2[52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1361  (\exu/alu_au/n16 [53], ds2[53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1362  (\exu/alu_au/n16 [54], ds2[54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1363  (\exu/alu_au/n16 [55], ds2[55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1364  (\exu/alu_au/n16 [56], ds2[56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1365  (\exu/alu_au/n16 [57], ds2[57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1366  (\exu/alu_au/n16 [58], ds2[58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1367  (\exu/alu_au/n16 [59], ds2[59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1368  (\exu/alu_au/n16 [60], ds2[60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1369  (\exu/alu_au/n16 [61], ds2[61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  or \exu/alu_au/u137  (\exu/alu_au/n54 [25], \exu/alu_au/n52 [25], \exu/alu_au/n53 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  not \exu/alu_au/u1370  (\exu/alu_au/n16 [62], ds2[62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  not \exu/alu_au/u1371  (\exu/alu_au/n16 [63], ds2[63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  or \exu/alu_au/u138  (\exu/alu_au/n54 [26], \exu/alu_au/n52 [26], \exu/alu_au/n53 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u139  (\exu/alu_au/n54 [27], \exu/alu_au/n52 [27], \exu/alu_au/n53 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u14  (\exu/alu_au/ds1_light_than_ds2 , \exu/alu_au/n8 , \exu/alu_au/n9 );  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(73)
  or \exu/alu_au/u140  (\exu/alu_au/n54 [28], \exu/alu_au/n52 [28], \exu/alu_au/n53 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u141  (\exu/alu_au/n54 [29], \exu/alu_au/n52 [29], \exu/alu_au/n53 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u142  (\exu/alu_au/n54 [30], \exu/alu_au/n52 [30], \exu/alu_au/n53 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u143  (\exu/alu_au/n54 [31], \exu/alu_au/n52 [31], \exu/alu_au/n53 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u144  (\exu/alu_au/n54 [32], \exu/alu_au/n52 [32], \exu/alu_au/n53 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u145  (\exu/alu_au/n54 [33], \exu/alu_au/n52 [33], \exu/alu_au/n53 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u146  (\exu/alu_au/n54 [34], \exu/alu_au/n52 [34], \exu/alu_au/n53 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u147  (\exu/alu_au/n54 [35], \exu/alu_au/n52 [35], \exu/alu_au/n53 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u148  (\exu/alu_au/n54 [36], \exu/alu_au/n52 [36], \exu/alu_au/n53 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u149  (\exu/alu_au/n54 [37], \exu/alu_au/n52 [37], \exu/alu_au/n53 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u15  (\exu/alu_data_mem_csr [5], \exu/alu_au/n54 [5], \exu/alu_au/n55 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u150  (\exu/alu_au/n54 [38], \exu/alu_au/n52 [38], \exu/alu_au/n53 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u151  (\exu/alu_au/n54 [39], \exu/alu_au/n52 [39], \exu/alu_au/n53 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u152  (\exu/alu_au/n54 [40], \exu/alu_au/n52 [40], \exu/alu_au/n53 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u153  (\exu/alu_au/n54 [41], \exu/alu_au/n52 [41], \exu/alu_au/n53 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u154  (\exu/alu_au/n54 [42], \exu/alu_au/n52 [42], \exu/alu_au/n53 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u155  (\exu/alu_au/n54 [43], \exu/alu_au/n52 [43], \exu/alu_au/n53 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u156  (\exu/alu_au/n54 [44], \exu/alu_au/n52 [44], \exu/alu_au/n53 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u157  (\exu/alu_au/n54 [45], \exu/alu_au/n52 [45], \exu/alu_au/n53 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u158  (\exu/alu_au/n54 [46], \exu/alu_au/n52 [46], \exu/alu_au/n53 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u159  (\exu/alu_au/n54 [47], \exu/alu_au/n52 [47], \exu/alu_au/n53 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  not \exu/alu_au/u16  (\exu/alu_au/n10 , ds1[63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(74)
  or \exu/alu_au/u160  (\exu/alu_au/n54 [48], \exu/alu_au/n52 [48], \exu/alu_au/n53 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u161  (\exu/alu_au/n54 [49], \exu/alu_au/n52 [49], \exu/alu_au/n53 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u162  (\exu/alu_au/n54 [50], \exu/alu_au/n52 [50], \exu/alu_au/n53 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u163  (\exu/alu_au/n54 [51], \exu/alu_au/n52 [51], \exu/alu_au/n53 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u164  (\exu/alu_au/n54 [52], \exu/alu_au/n52 [52], \exu/alu_au/n53 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u165  (\exu/alu_au/n54 [53], \exu/alu_au/n52 [53], \exu/alu_au/n53 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u166  (\exu/alu_au/n54 [54], \exu/alu_au/n52 [54], \exu/alu_au/n53 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u167  (\exu/alu_au/n54 [55], \exu/alu_au/n52 [55], \exu/alu_au/n53 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u168  (\exu/alu_au/n54 [56], \exu/alu_au/n52 [56], \exu/alu_au/n53 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u169  (\exu/alu_au/n54 [57], \exu/alu_au/n52 [57], \exu/alu_au/n53 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  and \exu/alu_au/u17  (\exu/alu_au/n11 , \exu/alu_au/n10 , ds2[63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(74)
  or \exu/alu_au/u170  (\exu/alu_au/n54 [58], \exu/alu_au/n52 [58], \exu/alu_au/n53 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u171  (\exu/alu_au/n54 [59], \exu/alu_au/n52 [59], \exu/alu_au/n53 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u172  (\exu/alu_au/n54 [60], \exu/alu_au/n52 [60], \exu/alu_au/n53 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u173  (\exu/alu_au/n54 [61], \exu/alu_au/n52 [61], \exu/alu_au/n53 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u174  (\exu/alu_au/n54 [62], \exu/alu_au/n52 [62], \exu/alu_au/n53 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u175  (\exu/alu_au/n54 [63], \exu/alu_au/n52 [63], \exu/alu_au/n53 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u176  (\exu/alu_au/n52 [1], \exu/alu_au/n50 [1], \exu/alu_au/n51 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u177  (\exu/alu_au/n52 [2], \exu/alu_au/n50 [2], \exu/alu_au/n51 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u178  (\exu/alu_au/n52 [3], \exu/alu_au/n50 [3], \exu/alu_au/n51 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u179  (\exu/alu_au/n52 [4], \exu/alu_au/n50 [4], \exu/alu_au/n51 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u18  (\exu/alu_data_mem_csr [4], \exu/alu_au/n54 [4], \exu/alu_au/n55 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u180  (\exu/alu_au/n52 [5], \exu/alu_au/n50 [5], \exu/alu_au/n51 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u181  (\exu/alu_au/n52 [6], \exu/alu_au/n50 [6], \exu/alu_au/n51 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u182  (\exu/alu_au/n52 [7], \exu/alu_au/n50 [7], \exu/alu_au/n51 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u183  (\exu/alu_au/n52 [8], \exu/alu_au/n50 [8], \exu/alu_au/n51 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u184  (\exu/alu_au/n52 [9], \exu/alu_au/n50 [9], \exu/alu_au/n51 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u185  (\exu/alu_au/n52 [10], \exu/alu_au/n50 [10], \exu/alu_au/n51 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u186  (\exu/alu_au/n52 [11], \exu/alu_au/n50 [11], \exu/alu_au/n51 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u187  (\exu/alu_au/n52 [12], \exu/alu_au/n50 [12], \exu/alu_au/n51 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u188  (\exu/alu_au/n52 [13], \exu/alu_au/n50 [13], \exu/alu_au/n51 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u189  (\exu/alu_au/n52 [14], \exu/alu_au/n50 [14], \exu/alu_au/n51 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u19  (\exu/alu_data_mem_csr [3], \exu/alu_au/n54 [3], \exu/alu_au/n55 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u190  (\exu/alu_au/n52 [15], \exu/alu_au/n50 [15], \exu/alu_au/n51 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u191  (\exu/alu_au/n52 [16], \exu/alu_au/n50 [16], \exu/alu_au/n51 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u192  (\exu/alu_au/n52 [17], \exu/alu_au/n50 [17], \exu/alu_au/n51 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u193  (\exu/alu_au/n52 [18], \exu/alu_au/n50 [18], \exu/alu_au/n51 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u194  (\exu/alu_au/n52 [19], \exu/alu_au/n50 [19], \exu/alu_au/n51 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u195  (\exu/alu_au/n52 [20], \exu/alu_au/n50 [20], \exu/alu_au/n51 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u196  (\exu/alu_au/n52 [21], \exu/alu_au/n50 [21], \exu/alu_au/n51 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u197  (\exu/alu_au/n52 [22], \exu/alu_au/n50 [22], \exu/alu_au/n51 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u198  (\exu/alu_au/n52 [23], \exu/alu_au/n50 [23], \exu/alu_au/n51 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u199  (\exu/alu_au/n52 [24], \exu/alu_au/n50 [24], \exu/alu_au/n51 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u2  (\exu/alu_data_mem_csr [8], \exu/alu_au/n54 [8], \exu/alu_au/n55 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  and \exu/alu_au/u20  (\exu/alu_au/n13 , \exu/alu_au/n4 , \exu/alu_au/n12 );  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(75)
  or \exu/alu_au/u200  (\exu/alu_au/n52 [25], \exu/alu_au/n50 [25], \exu/alu_au/n51 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u201  (\exu/alu_au/n52 [26], \exu/alu_au/n50 [26], \exu/alu_au/n51 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u202  (\exu/alu_au/n52 [27], \exu/alu_au/n50 [27], \exu/alu_au/n51 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u203  (\exu/alu_au/n52 [28], \exu/alu_au/n50 [28], \exu/alu_au/n51 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u204  (\exu/alu_au/n52 [29], \exu/alu_au/n50 [29], \exu/alu_au/n51 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u205  (\exu/alu_au/n52 [30], \exu/alu_au/n50 [30], \exu/alu_au/n51 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u206  (\exu/alu_au/n52 [31], \exu/alu_au/n50 [31], \exu/alu_au/n51 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u207  (\exu/alu_au/n52 [32], \exu/alu_au/n50 [32], \exu/alu_au/n51 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u208  (\exu/alu_au/n52 [33], \exu/alu_au/n50 [33], \exu/alu_au/n51 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u209  (\exu/alu_au/n52 [34], \exu/alu_au/n50 [34], \exu/alu_au/n51 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u21  (\exu/alu_au/n14 , \exu/alu_au/n11 , \exu/alu_au/n13 );  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(75)
  or \exu/alu_au/u210  (\exu/alu_au/n52 [35], \exu/alu_au/n50 [35], \exu/alu_au/n51 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u211  (\exu/alu_au/n52 [36], \exu/alu_au/n50 [36], \exu/alu_au/n51 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u212  (\exu/alu_au/n52 [37], \exu/alu_au/n50 [37], \exu/alu_au/n51 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u213  (\exu/alu_au/n52 [38], \exu/alu_au/n50 [38], \exu/alu_au/n51 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u214  (\exu/alu_au/n52 [39], \exu/alu_au/n50 [39], \exu/alu_au/n51 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u215  (\exu/alu_au/n52 [40], \exu/alu_au/n50 [40], \exu/alu_au/n51 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u216  (\exu/alu_au/n52 [41], \exu/alu_au/n50 [41], \exu/alu_au/n51 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u217  (\exu/alu_au/n52 [42], \exu/alu_au/n50 [42], \exu/alu_au/n51 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u218  (\exu/alu_au/n52 [43], \exu/alu_au/n50 [43], \exu/alu_au/n51 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u219  (\exu/alu_au/n52 [44], \exu/alu_au/n50 [44], \exu/alu_au/n51 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  and \exu/alu_au/u22  (\exu/alu_au/n15 , \exu/alu_au/n0 , \exu/alu_au/n14 );  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(75)
  or \exu/alu_au/u220  (\exu/alu_au/n52 [45], \exu/alu_au/n50 [45], \exu/alu_au/n51 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u221  (\exu/alu_au/n52 [46], \exu/alu_au/n50 [46], \exu/alu_au/n51 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u222  (\exu/alu_au/n52 [47], \exu/alu_au/n50 [47], \exu/alu_au/n51 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u223  (\exu/alu_au/n52 [48], \exu/alu_au/n50 [48], \exu/alu_au/n51 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u224  (\exu/alu_au/n52 [49], \exu/alu_au/n50 [49], \exu/alu_au/n51 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u225  (\exu/alu_au/n52 [50], \exu/alu_au/n50 [50], \exu/alu_au/n51 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u226  (\exu/alu_au/n52 [51], \exu/alu_au/n50 [51], \exu/alu_au/n51 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u227  (\exu/alu_au/n52 [52], \exu/alu_au/n50 [52], \exu/alu_au/n51 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u228  (\exu/alu_au/n52 [53], \exu/alu_au/n50 [53], \exu/alu_au/n51 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u229  (\exu/alu_au/n52 [54], \exu/alu_au/n50 [54], \exu/alu_au/n51 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u23  (\exu/alu_data_mem_csr [2], \exu/alu_au/n54 [2], \exu/alu_au/n55 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u230  (\exu/alu_au/n52 [55], \exu/alu_au/n50 [55], \exu/alu_au/n51 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u231  (\exu/alu_au/n52 [56], \exu/alu_au/n50 [56], \exu/alu_au/n51 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u232  (\exu/alu_au/n52 [57], \exu/alu_au/n50 [57], \exu/alu_au/n51 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u233  (\exu/alu_au/n52 [58], \exu/alu_au/n50 [58], \exu/alu_au/n51 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u234  (\exu/alu_au/n52 [59], \exu/alu_au/n50 [59], \exu/alu_au/n51 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u235  (\exu/alu_au/n52 [60], \exu/alu_au/n50 [60], \exu/alu_au/n51 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u236  (\exu/alu_au/n52 [61], \exu/alu_au/n50 [61], \exu/alu_au/n51 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u237  (\exu/alu_au/n52 [62], \exu/alu_au/n50 [62], \exu/alu_au/n51 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u238  (\exu/alu_au/n52 [63], \exu/alu_au/n50 [63], \exu/alu_au/n51 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u239  (\exu/alu_au/n50 [1], \exu/alu_au/n48 [1], \exu/alu_au/n49 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u24  (\exu/alu_data_mem_csr [1], \exu/alu_au/n54 [1], \exu/alu_au/n55 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u240  (\exu/alu_au/n50 [2], \exu/alu_au/n48 [2], \exu/alu_au/n49 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u241  (\exu/alu_au/n50 [3], \exu/alu_au/n48 [3], \exu/alu_au/n49 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u242  (\exu/alu_au/n50 [4], \exu/alu_au/n48 [4], \exu/alu_au/n49 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u243  (\exu/alu_au/n50 [5], \exu/alu_au/n48 [5], \exu/alu_au/n49 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u244  (\exu/alu_au/n50 [6], \exu/alu_au/n48 [6], \exu/alu_au/n49 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u245  (\exu/alu_au/n50 [7], \exu/alu_au/n48 [7], \exu/alu_au/n49 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u246  (\exu/alu_au/n50 [8], \exu/alu_au/n48 [8], \exu/alu_au/n49 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u247  (\exu/alu_au/n50 [9], \exu/alu_au/n48 [9], \exu/alu_au/n49 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u248  (\exu/alu_au/n50 [10], \exu/alu_au/n48 [10], \exu/alu_au/n49 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u249  (\exu/alu_au/n50 [11], \exu/alu_au/n48 [11], \exu/alu_au/n49 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u25  (\exu/alu_au/ds1_great_than_ds2 , \exu/alu_au/n15 , \exu/alu_au/n9 );  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(76)
  or \exu/alu_au/u250  (\exu/alu_au/n50 [12], \exu/alu_au/n48 [12], \exu/alu_au/n49 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u251  (\exu/alu_au/n50 [13], \exu/alu_au/n48 [13], \exu/alu_au/n49 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u252  (\exu/alu_au/n50 [14], \exu/alu_au/n48 [14], \exu/alu_au/n49 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u253  (\exu/alu_au/n50 [15], \exu/alu_au/n48 [15], \exu/alu_au/n49 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u254  (\exu/alu_au/n50 [16], \exu/alu_au/n48 [16], \exu/alu_au/n49 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u255  (\exu/alu_au/n50 [17], \exu/alu_au/n48 [17], \exu/alu_au/n49 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u256  (\exu/alu_au/n50 [18], \exu/alu_au/n48 [18], \exu/alu_au/n49 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u257  (\exu/alu_au/n50 [19], \exu/alu_au/n48 [19], \exu/alu_au/n49 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u258  (\exu/alu_au/n50 [20], \exu/alu_au/n48 [20], \exu/alu_au/n49 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u259  (\exu/alu_au/n50 [21], \exu/alu_au/n48 [21], \exu/alu_au/n49 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  not \exu/alu_au/u26  (\exu/alu_au/n16 [0], ds2[0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(79)
  or \exu/alu_au/u260  (\exu/alu_au/n50 [22], \exu/alu_au/n48 [22], \exu/alu_au/n49 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u261  (\exu/alu_au/n50 [23], \exu/alu_au/n48 [23], \exu/alu_au/n49 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u262  (\exu/alu_au/n50 [24], \exu/alu_au/n48 [24], \exu/alu_au/n49 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u263  (\exu/alu_au/n50 [25], \exu/alu_au/n48 [25], \exu/alu_au/n49 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u264  (\exu/alu_au/n50 [26], \exu/alu_au/n48 [26], \exu/alu_au/n49 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u265  (\exu/alu_au/n50 [27], \exu/alu_au/n48 [27], \exu/alu_au/n49 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u266  (\exu/alu_au/n50 [28], \exu/alu_au/n48 [28], \exu/alu_au/n49 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u267  (\exu/alu_au/n50 [29], \exu/alu_au/n48 [29], \exu/alu_au/n49 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u268  (\exu/alu_au/n50 [30], \exu/alu_au/n48 [30], \exu/alu_au/n49 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u269  (\exu/alu_au/n50 [31], \exu/alu_au/n48 [31], \exu/alu_au/n49 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u270  (\exu/alu_au/n50 [32], \exu/alu_au/n48 [32], \exu/alu_au/n49 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u271  (\exu/alu_au/n50 [33], \exu/alu_au/n48 [33], \exu/alu_au/n49 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u272  (\exu/alu_au/n50 [34], \exu/alu_au/n48 [34], \exu/alu_au/n49 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u273  (\exu/alu_au/n50 [35], \exu/alu_au/n48 [35], \exu/alu_au/n49 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u274  (\exu/alu_au/n50 [36], \exu/alu_au/n48 [36], \exu/alu_au/n49 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u275  (\exu/alu_au/n50 [37], \exu/alu_au/n48 [37], \exu/alu_au/n49 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u276  (\exu/alu_au/n50 [38], \exu/alu_au/n48 [38], \exu/alu_au/n49 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u277  (\exu/alu_au/n50 [39], \exu/alu_au/n48 [39], \exu/alu_au/n49 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u278  (\exu/alu_au/n50 [40], \exu/alu_au/n48 [40], \exu/alu_au/n49 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u279  (\exu/alu_au/n50 [41], \exu/alu_au/n48 [41], \exu/alu_au/n49 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u28  (\exu/alu_data_mem_csr [0], \exu/alu_au/n54 [0], \exu/alu_au/n55 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u280  (\exu/alu_au/n50 [42], \exu/alu_au/n48 [42], \exu/alu_au/n49 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u281  (\exu/alu_au/n50 [43], \exu/alu_au/n48 [43], \exu/alu_au/n49 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u282  (\exu/alu_au/n50 [44], \exu/alu_au/n48 [44], \exu/alu_au/n49 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u283  (\exu/alu_au/n50 [45], \exu/alu_au/n48 [45], \exu/alu_au/n49 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u284  (\exu/alu_au/n50 [46], \exu/alu_au/n48 [46], \exu/alu_au/n49 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u285  (\exu/alu_au/n50 [47], \exu/alu_au/n48 [47], \exu/alu_au/n49 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u286  (\exu/alu_au/n50 [48], \exu/alu_au/n48 [48], \exu/alu_au/n49 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u287  (\exu/alu_au/n50 [49], \exu/alu_au/n48 [49], \exu/alu_au/n49 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u288  (\exu/alu_au/n50 [50], \exu/alu_au/n48 [50], \exu/alu_au/n49 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u289  (\exu/alu_au/n50 [51], \exu/alu_au/n48 [51], \exu/alu_au/n49 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u290  (\exu/alu_au/n50 [52], \exu/alu_au/n48 [52], \exu/alu_au/n49 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u291  (\exu/alu_au/n50 [53], \exu/alu_au/n48 [53], \exu/alu_au/n49 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u292  (\exu/alu_au/n50 [54], \exu/alu_au/n48 [54], \exu/alu_au/n49 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u293  (\exu/alu_au/n50 [55], \exu/alu_au/n48 [55], \exu/alu_au/n49 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u294  (\exu/alu_au/n50 [56], \exu/alu_au/n48 [56], \exu/alu_au/n49 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u295  (\exu/alu_au/n50 [57], \exu/alu_au/n48 [57], \exu/alu_au/n49 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u296  (\exu/alu_au/n50 [58], \exu/alu_au/n48 [58], \exu/alu_au/n49 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u297  (\exu/alu_au/n50 [59], \exu/alu_au/n48 [59], \exu/alu_au/n49 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u298  (\exu/alu_au/n50 [60], \exu/alu_au/n48 [60], \exu/alu_au/n49 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u299  (\exu/alu_au/n50 [61], \exu/alu_au/n48 [61], \exu/alu_au/n49 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u3  (\exu/alu_data_mem_csr [7], \exu/alu_au/n54 [7], \exu/alu_au/n55 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  and \exu/alu_au/u30  (\exu/alu_au/alu_and [0], ds1[0], \exu/alu_au/n18 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(87)
  or \exu/alu_au/u300  (\exu/alu_au/n50 [62], \exu/alu_au/n48 [62], \exu/alu_au/n49 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u301  (\exu/alu_au/n50 [63], \exu/alu_au/n48 [63], \exu/alu_au/n49 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u302  (\exu/alu_au/n48 [1], \exu/alu_au/n46 [1], \exu/alu_au/n47 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u303  (\exu/alu_au/n48 [2], \exu/alu_au/n46 [2], \exu/alu_au/n47 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u304  (\exu/alu_au/n48 [3], \exu/alu_au/n46 [3], \exu/alu_au/n47 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u305  (\exu/alu_au/n48 [4], \exu/alu_au/n46 [4], \exu/alu_au/n47 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u306  (\exu/alu_au/n48 [5], \exu/alu_au/n46 [5], \exu/alu_au/n47 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u307  (\exu/alu_au/n48 [6], \exu/alu_au/n46 [6], \exu/alu_au/n47 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u308  (\exu/alu_au/n48 [7], \exu/alu_au/n46 [7], \exu/alu_au/n47 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u309  (\exu/alu_au/n48 [8], \exu/alu_au/n46 [8], \exu/alu_au/n47 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u31  (\exu/alu_au/alu_or [0], ds1[0], ds2[0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(88)
  or \exu/alu_au/u310  (\exu/alu_au/n48 [9], \exu/alu_au/n46 [9], \exu/alu_au/n47 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u311  (\exu/alu_au/n48 [10], \exu/alu_au/n46 [10], \exu/alu_au/n47 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u312  (\exu/alu_au/n48 [11], \exu/alu_au/n46 [11], \exu/alu_au/n47 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u313  (\exu/alu_au/n48 [12], \exu/alu_au/n46 [12], \exu/alu_au/n47 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u314  (\exu/alu_au/n48 [13], \exu/alu_au/n46 [13], \exu/alu_au/n47 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u315  (\exu/alu_au/n48 [14], \exu/alu_au/n46 [14], \exu/alu_au/n47 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u316  (\exu/alu_au/n48 [15], \exu/alu_au/n46 [15], \exu/alu_au/n47 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u317  (\exu/alu_au/n48 [16], \exu/alu_au/n46 [16], \exu/alu_au/n47 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u318  (\exu/alu_au/n48 [17], \exu/alu_au/n46 [17], \exu/alu_au/n47 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u319  (\exu/alu_au/n48 [18], \exu/alu_au/n46 [18], \exu/alu_au/n47 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  xor \exu/alu_au/u32  (\exu/alu_au/alu_xor [0], ds1[0], ds2[0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(89)
  or \exu/alu_au/u320  (\exu/alu_au/n48 [19], \exu/alu_au/n46 [19], \exu/alu_au/n47 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u321  (\exu/alu_au/n48 [20], \exu/alu_au/n46 [20], \exu/alu_au/n47 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u322  (\exu/alu_au/n48 [21], \exu/alu_au/n46 [21], \exu/alu_au/n47 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u323  (\exu/alu_au/n48 [22], \exu/alu_au/n46 [22], \exu/alu_au/n47 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u324  (\exu/alu_au/n48 [23], \exu/alu_au/n46 [23], \exu/alu_au/n47 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u325  (\exu/alu_au/n48 [24], \exu/alu_au/n46 [24], \exu/alu_au/n47 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u326  (\exu/alu_au/n48 [25], \exu/alu_au/n46 [25], \exu/alu_au/n47 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u327  (\exu/alu_au/n48 [26], \exu/alu_au/n46 [26], \exu/alu_au/n47 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u328  (\exu/alu_au/n48 [27], \exu/alu_au/n46 [27], \exu/alu_au/n47 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u329  (\exu/alu_au/n48 [28], \exu/alu_au/n46 [28], \exu/alu_au/n47 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u330  (\exu/alu_au/n48 [29], \exu/alu_au/n46 [29], \exu/alu_au/n47 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u331  (\exu/alu_au/n48 [30], \exu/alu_au/n46 [30], \exu/alu_au/n47 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u332  (\exu/alu_au/n48 [31], \exu/alu_au/n46 [31], \exu/alu_au/n47 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u333  (\exu/alu_au/n48 [32], \exu/alu_au/n46 [32], \exu/alu_au/n47 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u334  (\exu/alu_au/n48 [33], \exu/alu_au/n46 [33], \exu/alu_au/n47 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u335  (\exu/alu_au/n48 [34], \exu/alu_au/n46 [34], \exu/alu_au/n47 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u336  (\exu/alu_au/n48 [35], \exu/alu_au/n46 [35], \exu/alu_au/n47 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u337  (\exu/alu_au/n48 [36], \exu/alu_au/n46 [36], \exu/alu_au/n47 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u338  (\exu/alu_au/n48 [37], \exu/alu_au/n46 [37], \exu/alu_au/n47 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u339  (\exu/alu_au/n48 [38], \exu/alu_au/n46 [38], \exu/alu_au/n47 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u340  (\exu/alu_au/n48 [39], \exu/alu_au/n46 [39], \exu/alu_au/n47 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u341  (\exu/alu_au/n48 [40], \exu/alu_au/n46 [40], \exu/alu_au/n47 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u342  (\exu/alu_au/n48 [41], \exu/alu_au/n46 [41], \exu/alu_au/n47 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u343  (\exu/alu_au/n48 [42], \exu/alu_au/n46 [42], \exu/alu_au/n47 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u344  (\exu/alu_au/n48 [43], \exu/alu_au/n46 [43], \exu/alu_au/n47 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u345  (\exu/alu_au/n48 [44], \exu/alu_au/n46 [44], \exu/alu_au/n47 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u346  (\exu/alu_au/n48 [45], \exu/alu_au/n46 [45], \exu/alu_au/n47 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u347  (\exu/alu_au/n48 [46], \exu/alu_au/n46 [46], \exu/alu_au/n47 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u348  (\exu/alu_au/n48 [47], \exu/alu_au/n46 [47], \exu/alu_au/n47 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u349  (\exu/alu_au/n48 [48], \exu/alu_au/n46 [48], \exu/alu_au/n47 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u350  (\exu/alu_au/n48 [49], \exu/alu_au/n46 [49], \exu/alu_au/n47 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u351  (\exu/alu_au/n48 [50], \exu/alu_au/n46 [50], \exu/alu_au/n47 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u352  (\exu/alu_au/n48 [51], \exu/alu_au/n46 [51], \exu/alu_au/n47 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u353  (\exu/alu_au/n48 [52], \exu/alu_au/n46 [52], \exu/alu_au/n47 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u354  (\exu/alu_au/n48 [53], \exu/alu_au/n46 [53], \exu/alu_au/n47 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u355  (\exu/alu_au/n48 [54], \exu/alu_au/n46 [54], \exu/alu_au/n47 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u356  (\exu/alu_au/n48 [55], \exu/alu_au/n46 [55], \exu/alu_au/n47 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u357  (\exu/alu_au/n48 [56], \exu/alu_au/n46 [56], \exu/alu_au/n47 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u358  (\exu/alu_au/n48 [57], \exu/alu_au/n46 [57], \exu/alu_au/n47 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u359  (\exu/alu_au/n48 [58], \exu/alu_au/n46 [58], \exu/alu_au/n47 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u360  (\exu/alu_au/n48 [59], \exu/alu_au/n46 [59], \exu/alu_au/n47 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u361  (\exu/alu_au/n48 [60], \exu/alu_au/n46 [60], \exu/alu_au/n47 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u362  (\exu/alu_au/n48 [61], \exu/alu_au/n46 [61], \exu/alu_au/n47 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u363  (\exu/alu_au/n48 [62], \exu/alu_au/n46 [62], \exu/alu_au/n47 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u364  (\exu/alu_au/n48 [63], \exu/alu_au/n46 [63], \exu/alu_au/n47 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u365  (\exu/alu_au/n46 [1], \exu/alu_au/n43 [1], \exu/alu_au/n45 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u366  (\exu/alu_au/n46 [2], \exu/alu_au/n43 [2], \exu/alu_au/n45 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u367  (\exu/alu_au/n46 [3], \exu/alu_au/n43 [3], \exu/alu_au/n45 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u368  (\exu/alu_au/n46 [4], \exu/alu_au/n43 [4], \exu/alu_au/n45 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u369  (\exu/alu_au/n46 [5], \exu/alu_au/n43 [5], \exu/alu_au/n45 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u370  (\exu/alu_au/n46 [6], \exu/alu_au/n43 [6], \exu/alu_au/n45 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u371  (\exu/alu_au/n46 [7], \exu/alu_au/n43 [7], \exu/alu_au/n45 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u372  (\exu/alu_au/n46 [8], \exu/alu_au/n43 [8], \exu/alu_au/n45 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u373  (\exu/alu_au/n46 [9], \exu/alu_au/n43 [9], \exu/alu_au/n45 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u374  (\exu/alu_au/n46 [10], \exu/alu_au/n43 [10], \exu/alu_au/n45 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u375  (\exu/alu_au/n46 [11], \exu/alu_au/n43 [11], \exu/alu_au/n45 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u376  (\exu/alu_au/n46 [12], \exu/alu_au/n43 [12], \exu/alu_au/n45 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u377  (\exu/alu_au/n46 [13], \exu/alu_au/n43 [13], \exu/alu_au/n45 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u378  (\exu/alu_au/n46 [14], \exu/alu_au/n43 [14], \exu/alu_au/n45 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u379  (\exu/alu_au/n46 [15], \exu/alu_au/n43 [15], \exu/alu_au/n45 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u380  (\exu/alu_au/n46 [16], \exu/alu_au/n43 [16], \exu/alu_au/n45 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u381  (\exu/alu_au/n46 [17], \exu/alu_au/n43 [17], \exu/alu_au/n45 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u382  (\exu/alu_au/n46 [18], \exu/alu_au/n43 [18], \exu/alu_au/n45 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u383  (\exu/alu_au/n46 [19], \exu/alu_au/n43 [19], \exu/alu_au/n45 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u384  (\exu/alu_au/n46 [20], \exu/alu_au/n43 [20], \exu/alu_au/n45 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u385  (\exu/alu_au/n46 [21], \exu/alu_au/n43 [21], \exu/alu_au/n45 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u386  (\exu/alu_au/n46 [22], \exu/alu_au/n43 [22], \exu/alu_au/n45 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u387  (\exu/alu_au/n46 [23], \exu/alu_au/n43 [23], \exu/alu_au/n45 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u388  (\exu/alu_au/n46 [24], \exu/alu_au/n43 [24], \exu/alu_au/n45 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u389  (\exu/alu_au/n46 [25], \exu/alu_au/n43 [25], \exu/alu_au/n45 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u390  (\exu/alu_au/n46 [26], \exu/alu_au/n43 [26], \exu/alu_au/n45 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u391  (\exu/alu_au/n46 [27], \exu/alu_au/n43 [27], \exu/alu_au/n45 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u392  (\exu/alu_au/n46 [28], \exu/alu_au/n43 [28], \exu/alu_au/n45 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u393  (\exu/alu_au/n46 [29], \exu/alu_au/n43 [29], \exu/alu_au/n45 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u394  (\exu/alu_au/n46 [30], \exu/alu_au/n43 [30], \exu/alu_au/n45 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u395  (\exu/alu_au/n46 [31], \exu/alu_au/n43 [31], \exu/alu_au/n45 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u396  (\exu/alu_au/n46 [32], \exu/alu_au/n43 [32], \exu/alu_au/n45 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u397  (\exu/alu_au/n46 [33], \exu/alu_au/n43 [33], \exu/alu_au/n45 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u398  (\exu/alu_au/n46 [34], \exu/alu_au/n43 [34], \exu/alu_au/n45 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u399  (\exu/alu_au/n46 [35], \exu/alu_au/n43 [35], \exu/alu_au/n45 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  not \exu/alu_au/u4  (\exu/alu_au/n0 , unsign);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(71)
  or \exu/alu_au/u400  (\exu/alu_au/n46 [36], \exu/alu_au/n43 [36], \exu/alu_au/n45 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u401  (\exu/alu_au/n46 [37], \exu/alu_au/n43 [37], \exu/alu_au/n45 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u402  (\exu/alu_au/n46 [38], \exu/alu_au/n43 [38], \exu/alu_au/n45 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u403  (\exu/alu_au/n46 [39], \exu/alu_au/n43 [39], \exu/alu_au/n45 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u404  (\exu/alu_au/n46 [40], \exu/alu_au/n43 [40], \exu/alu_au/n45 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u405  (\exu/alu_au/n46 [41], \exu/alu_au/n43 [41], \exu/alu_au/n45 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u406  (\exu/alu_au/n46 [42], \exu/alu_au/n43 [42], \exu/alu_au/n45 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u407  (\exu/alu_au/n46 [43], \exu/alu_au/n43 [43], \exu/alu_au/n45 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u408  (\exu/alu_au/n46 [44], \exu/alu_au/n43 [44], \exu/alu_au/n45 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u409  (\exu/alu_au/n46 [45], \exu/alu_au/n43 [45], \exu/alu_au/n45 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u410  (\exu/alu_au/n46 [46], \exu/alu_au/n43 [46], \exu/alu_au/n45 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u411  (\exu/alu_au/n46 [47], \exu/alu_au/n43 [47], \exu/alu_au/n45 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u412  (\exu/alu_au/n46 [48], \exu/alu_au/n43 [48], \exu/alu_au/n45 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u413  (\exu/alu_au/n46 [49], \exu/alu_au/n43 [49], \exu/alu_au/n45 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u414  (\exu/alu_au/n46 [50], \exu/alu_au/n43 [50], \exu/alu_au/n45 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u415  (\exu/alu_au/n46 [51], \exu/alu_au/n43 [51], \exu/alu_au/n45 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u416  (\exu/alu_au/n46 [52], \exu/alu_au/n43 [52], \exu/alu_au/n45 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u417  (\exu/alu_au/n46 [53], \exu/alu_au/n43 [53], \exu/alu_au/n45 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u418  (\exu/alu_au/n46 [54], \exu/alu_au/n43 [54], \exu/alu_au/n45 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u419  (\exu/alu_au/n46 [55], \exu/alu_au/n43 [55], \exu/alu_au/n45 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u420  (\exu/alu_au/n46 [56], \exu/alu_au/n43 [56], \exu/alu_au/n45 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u421  (\exu/alu_au/n46 [57], \exu/alu_au/n43 [57], \exu/alu_au/n45 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u422  (\exu/alu_au/n46 [58], \exu/alu_au/n43 [58], \exu/alu_au/n45 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u423  (\exu/alu_au/n46 [59], \exu/alu_au/n43 [59], \exu/alu_au/n45 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u424  (\exu/alu_au/n46 [60], \exu/alu_au/n43 [60], \exu/alu_au/n45 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u425  (\exu/alu_au/n46 [61], \exu/alu_au/n43 [61], \exu/alu_au/n45 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u426  (\exu/alu_au/n46 [62], \exu/alu_au/n43 [62], \exu/alu_au/n45 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u427  (\exu/alu_au/n46 [63], \exu/alu_au/n43 [63], \exu/alu_au/n45 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u45  (\exu/alu_au/n30 [0], \exu/alu_au/n28 [0], \exu/alu_au/n29 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u46  (\exu/alu_au/n32 [0], \exu/alu_au/n30 [0], \exu/alu_au/n31 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u47  (\exu/alu_au/n34 [0], \exu/alu_au/n32 [0], \exu/alu_au/n33 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u48  (\exu/alu_au/n36 [0], \exu/alu_au/n34 [0], \exu/alu_au/n35 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u49  (\exu/alu_au/n38 [0], \exu/alu_au/n36 [0], \exu/alu_au/n37 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u50  (\exu/alu_au/n40 [0], \exu/alu_au/n38 [0], \exu/alu_au/n39 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(105)
  or \exu/alu_au/u53  (\exu/alu_au/n46 [0], \exu/alu_au/n43 [0], \exu/alu_au/n45 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(111)
  or \exu/alu_au/u54  (\exu/alu_au/n48 [0], \exu/alu_au/n46 [0], \exu/alu_au/n47 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(112)
  or \exu/alu_au/u55  (\exu/alu_au/n50 [0], \exu/alu_au/n48 [0], \exu/alu_au/n49 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(113)
  or \exu/alu_au/u56  (\exu/alu_au/n52 [0], \exu/alu_au/n50 [0], \exu/alu_au/n51 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(114)
  or \exu/alu_au/u57  (\exu/alu_au/n54 [0], \exu/alu_au/n52 [0], \exu/alu_au/n53 [0]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(115)
  or \exu/alu_au/u58  (\exu/alu_data_mem_csr [9], \exu/alu_au/n54 [9], \exu/alu_au/n55 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u59  (\exu/alu_data_mem_csr [10], \exu/alu_au/n54 [10], \exu/alu_au/n55 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  and \exu/alu_au/u6  (\exu/alu_au/n2 , ds1[63], \exu/alu_au/n16 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(71)
  or \exu/alu_au/u60  (\exu/alu_data_mem_csr [11], \exu/alu_au/n54 [11], \exu/alu_au/n55 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u61  (\exu/alu_data_mem_csr [12], \exu/alu_au/n54 [12], \exu/alu_au/n55 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u617  (\exu/alu_au/n38 [1], \exu/alu_au/n36 [1], \exu/alu_au/n37 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u618  (\exu/alu_au/n38 [2], \exu/alu_au/n36 [2], \exu/alu_au/n37 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u619  (\exu/alu_au/n38 [3], \exu/alu_au/n36 [3], \exu/alu_au/n37 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u62  (\exu/alu_data_mem_csr [13], \exu/alu_au/n54 [13], \exu/alu_au/n55 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u620  (\exu/alu_au/n38 [4], \exu/alu_au/n36 [4], \exu/alu_au/n37 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u621  (\exu/alu_au/n38 [5], \exu/alu_au/n36 [5], \exu/alu_au/n37 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u622  (\exu/alu_au/n38 [6], \exu/alu_au/n36 [6], \exu/alu_au/n37 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u623  (\exu/alu_au/n38 [7], \exu/alu_au/n36 [7], \exu/alu_au/n37 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u624  (\exu/alu_au/n38 [8], \exu/alu_au/n36 [8], \exu/alu_au/n37 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u625  (\exu/alu_au/n38 [9], \exu/alu_au/n36 [9], \exu/alu_au/n37 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u626  (\exu/alu_au/n38 [10], \exu/alu_au/n36 [10], \exu/alu_au/n37 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u627  (\exu/alu_au/n38 [11], \exu/alu_au/n36 [11], \exu/alu_au/n37 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u628  (\exu/alu_au/n38 [12], \exu/alu_au/n36 [12], \exu/alu_au/n37 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u629  (\exu/alu_au/n38 [13], \exu/alu_au/n36 [13], \exu/alu_au/n37 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u63  (\exu/alu_data_mem_csr [14], \exu/alu_au/n54 [14], \exu/alu_au/n55 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u630  (\exu/alu_au/n38 [14], \exu/alu_au/n36 [14], \exu/alu_au/n37 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u631  (\exu/alu_au/n38 [15], \exu/alu_au/n36 [15], \exu/alu_au/n37 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u632  (\exu/alu_au/n38 [16], \exu/alu_au/n36 [16], \exu/alu_au/n37 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u633  (\exu/alu_au/n38 [17], \exu/alu_au/n36 [17], \exu/alu_au/n37 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u634  (\exu/alu_au/n38 [18], \exu/alu_au/n36 [18], \exu/alu_au/n37 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u635  (\exu/alu_au/n38 [19], \exu/alu_au/n36 [19], \exu/alu_au/n37 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u636  (\exu/alu_au/n38 [20], \exu/alu_au/n36 [20], \exu/alu_au/n37 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u637  (\exu/alu_au/n38 [21], \exu/alu_au/n36 [21], \exu/alu_au/n37 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u638  (\exu/alu_au/n38 [22], \exu/alu_au/n36 [22], \exu/alu_au/n37 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u639  (\exu/alu_au/n38 [23], \exu/alu_au/n36 [23], \exu/alu_au/n37 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u64  (\exu/alu_data_mem_csr [15], \exu/alu_au/n54 [15], \exu/alu_au/n55 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u640  (\exu/alu_au/n38 [24], \exu/alu_au/n36 [24], \exu/alu_au/n37 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u641  (\exu/alu_au/n38 [25], \exu/alu_au/n36 [25], \exu/alu_au/n37 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u642  (\exu/alu_au/n38 [26], \exu/alu_au/n36 [26], \exu/alu_au/n37 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u643  (\exu/alu_au/n38 [27], \exu/alu_au/n36 [27], \exu/alu_au/n37 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u644  (\exu/alu_au/n38 [28], \exu/alu_au/n36 [28], \exu/alu_au/n37 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u645  (\exu/alu_au/n38 [29], \exu/alu_au/n36 [29], \exu/alu_au/n37 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u646  (\exu/alu_au/n38 [30], \exu/alu_au/n36 [30], \exu/alu_au/n37 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u647  (\exu/alu_au/n38 [31], \exu/alu_au/n36 [31], \exu/alu_au/n37 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u648  (\exu/alu_au/n38 [32], \exu/alu_au/n36 [32], \exu/alu_au/n37 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u649  (\exu/alu_au/n38 [33], \exu/alu_au/n36 [33], \exu/alu_au/n37 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u65  (\exu/alu_data_mem_csr [16], \exu/alu_au/n54 [16], \exu/alu_au/n55 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u650  (\exu/alu_au/n38 [34], \exu/alu_au/n36 [34], \exu/alu_au/n37 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u651  (\exu/alu_au/n38 [35], \exu/alu_au/n36 [35], \exu/alu_au/n37 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u652  (\exu/alu_au/n38 [36], \exu/alu_au/n36 [36], \exu/alu_au/n37 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u653  (\exu/alu_au/n38 [37], \exu/alu_au/n36 [37], \exu/alu_au/n37 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u654  (\exu/alu_au/n38 [38], \exu/alu_au/n36 [38], \exu/alu_au/n37 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u655  (\exu/alu_au/n38 [39], \exu/alu_au/n36 [39], \exu/alu_au/n37 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u656  (\exu/alu_au/n38 [40], \exu/alu_au/n36 [40], \exu/alu_au/n37 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u657  (\exu/alu_au/n38 [41], \exu/alu_au/n36 [41], \exu/alu_au/n37 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u658  (\exu/alu_au/n38 [42], \exu/alu_au/n36 [42], \exu/alu_au/n37 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u659  (\exu/alu_au/n38 [43], \exu/alu_au/n36 [43], \exu/alu_au/n37 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u66  (\exu/alu_data_mem_csr [17], \exu/alu_au/n54 [17], \exu/alu_au/n55 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u660  (\exu/alu_au/n38 [44], \exu/alu_au/n36 [44], \exu/alu_au/n37 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u661  (\exu/alu_au/n38 [45], \exu/alu_au/n36 [45], \exu/alu_au/n37 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u662  (\exu/alu_au/n38 [46], \exu/alu_au/n36 [46], \exu/alu_au/n37 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u663  (\exu/alu_au/n38 [47], \exu/alu_au/n36 [47], \exu/alu_au/n37 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u664  (\exu/alu_au/n38 [48], \exu/alu_au/n36 [48], \exu/alu_au/n37 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u665  (\exu/alu_au/n38 [49], \exu/alu_au/n36 [49], \exu/alu_au/n37 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u666  (\exu/alu_au/n38 [50], \exu/alu_au/n36 [50], \exu/alu_au/n37 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u667  (\exu/alu_au/n38 [51], \exu/alu_au/n36 [51], \exu/alu_au/n37 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u668  (\exu/alu_au/n38 [52], \exu/alu_au/n36 [52], \exu/alu_au/n37 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u669  (\exu/alu_au/n38 [53], \exu/alu_au/n36 [53], \exu/alu_au/n37 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u67  (\exu/alu_data_mem_csr [18], \exu/alu_au/n54 [18], \exu/alu_au/n55 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u670  (\exu/alu_au/n38 [54], \exu/alu_au/n36 [54], \exu/alu_au/n37 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u671  (\exu/alu_au/n38 [55], \exu/alu_au/n36 [55], \exu/alu_au/n37 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u672  (\exu/alu_au/n38 [56], \exu/alu_au/n36 [56], \exu/alu_au/n37 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u673  (\exu/alu_au/n38 [57], \exu/alu_au/n36 [57], \exu/alu_au/n37 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u674  (\exu/alu_au/n38 [58], \exu/alu_au/n36 [58], \exu/alu_au/n37 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u675  (\exu/alu_au/n38 [59], \exu/alu_au/n36 [59], \exu/alu_au/n37 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u676  (\exu/alu_au/n38 [60], \exu/alu_au/n36 [60], \exu/alu_au/n37 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u677  (\exu/alu_au/n38 [61], \exu/alu_au/n36 [61], \exu/alu_au/n37 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u678  (\exu/alu_au/n38 [62], \exu/alu_au/n36 [62], \exu/alu_au/n37 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u679  (\exu/alu_au/n38 [63], \exu/alu_au/n36 [63], \exu/alu_au/n37 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(104)
  or \exu/alu_au/u68  (\exu/alu_data_mem_csr [19], \exu/alu_au/n54 [19], \exu/alu_au/n55 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u680  (\exu/alu_au/n36 [1], \exu/alu_au/n34 [1], \exu/alu_au/n35 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u681  (\exu/alu_au/n36 [2], \exu/alu_au/n34 [2], \exu/alu_au/n35 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u682  (\exu/alu_au/n36 [3], \exu/alu_au/n34 [3], \exu/alu_au/n35 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u683  (\exu/alu_au/n36 [4], \exu/alu_au/n34 [4], \exu/alu_au/n35 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u684  (\exu/alu_au/n36 [5], \exu/alu_au/n34 [5], \exu/alu_au/n35 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u685  (\exu/alu_au/n36 [6], \exu/alu_au/n34 [6], \exu/alu_au/n35 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u686  (\exu/alu_au/n36 [7], \exu/alu_au/n34 [7], \exu/alu_au/n35 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u687  (\exu/alu_au/n36 [8], \exu/alu_au/n34 [8], \exu/alu_au/n35 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u688  (\exu/alu_au/n36 [9], \exu/alu_au/n34 [9], \exu/alu_au/n35 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u689  (\exu/alu_au/n36 [10], \exu/alu_au/n34 [10], \exu/alu_au/n35 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u69  (\exu/alu_data_mem_csr [20], \exu/alu_au/n54 [20], \exu/alu_au/n55 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u690  (\exu/alu_au/n36 [11], \exu/alu_au/n34 [11], \exu/alu_au/n35 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u691  (\exu/alu_au/n36 [12], \exu/alu_au/n34 [12], \exu/alu_au/n35 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u692  (\exu/alu_au/n36 [13], \exu/alu_au/n34 [13], \exu/alu_au/n35 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u693  (\exu/alu_au/n36 [14], \exu/alu_au/n34 [14], \exu/alu_au/n35 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u694  (\exu/alu_au/n36 [15], \exu/alu_au/n34 [15], \exu/alu_au/n35 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u695  (\exu/alu_au/n36 [16], \exu/alu_au/n34 [16], \exu/alu_au/n35 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u696  (\exu/alu_au/n36 [17], \exu/alu_au/n34 [17], \exu/alu_au/n35 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u697  (\exu/alu_au/n36 [18], \exu/alu_au/n34 [18], \exu/alu_au/n35 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u698  (\exu/alu_au/n36 [19], \exu/alu_au/n34 [19], \exu/alu_au/n35 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u699  (\exu/alu_au/n36 [20], \exu/alu_au/n34 [20], \exu/alu_au/n35 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u70  (\exu/alu_data_mem_csr [21], \exu/alu_au/n54 [21], \exu/alu_au/n55 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u700  (\exu/alu_au/n36 [21], \exu/alu_au/n34 [21], \exu/alu_au/n35 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u701  (\exu/alu_au/n36 [22], \exu/alu_au/n34 [22], \exu/alu_au/n35 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u702  (\exu/alu_au/n36 [23], \exu/alu_au/n34 [23], \exu/alu_au/n35 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u703  (\exu/alu_au/n36 [24], \exu/alu_au/n34 [24], \exu/alu_au/n35 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u704  (\exu/alu_au/n36 [25], \exu/alu_au/n34 [25], \exu/alu_au/n35 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u705  (\exu/alu_au/n36 [26], \exu/alu_au/n34 [26], \exu/alu_au/n35 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u706  (\exu/alu_au/n36 [27], \exu/alu_au/n34 [27], \exu/alu_au/n35 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u707  (\exu/alu_au/n36 [28], \exu/alu_au/n34 [28], \exu/alu_au/n35 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u708  (\exu/alu_au/n36 [29], \exu/alu_au/n34 [29], \exu/alu_au/n35 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u709  (\exu/alu_au/n36 [30], \exu/alu_au/n34 [30], \exu/alu_au/n35 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u71  (\exu/alu_data_mem_csr [22], \exu/alu_au/n54 [22], \exu/alu_au/n55 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u710  (\exu/alu_au/n36 [31], \exu/alu_au/n34 [31], \exu/alu_au/n35 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u711  (\exu/alu_au/n36 [32], \exu/alu_au/n34 [32], \exu/alu_au/n35 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u712  (\exu/alu_au/n36 [33], \exu/alu_au/n34 [33], \exu/alu_au/n35 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u713  (\exu/alu_au/n36 [34], \exu/alu_au/n34 [34], \exu/alu_au/n35 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u714  (\exu/alu_au/n36 [35], \exu/alu_au/n34 [35], \exu/alu_au/n35 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u715  (\exu/alu_au/n36 [36], \exu/alu_au/n34 [36], \exu/alu_au/n35 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u716  (\exu/alu_au/n36 [37], \exu/alu_au/n34 [37], \exu/alu_au/n35 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u717  (\exu/alu_au/n36 [38], \exu/alu_au/n34 [38], \exu/alu_au/n35 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u718  (\exu/alu_au/n36 [39], \exu/alu_au/n34 [39], \exu/alu_au/n35 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u719  (\exu/alu_au/n36 [40], \exu/alu_au/n34 [40], \exu/alu_au/n35 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u72  (\exu/alu_data_mem_csr [23], \exu/alu_au/n54 [23], \exu/alu_au/n55 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u720  (\exu/alu_au/n36 [41], \exu/alu_au/n34 [41], \exu/alu_au/n35 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u721  (\exu/alu_au/n36 [42], \exu/alu_au/n34 [42], \exu/alu_au/n35 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u722  (\exu/alu_au/n36 [43], \exu/alu_au/n34 [43], \exu/alu_au/n35 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u723  (\exu/alu_au/n36 [44], \exu/alu_au/n34 [44], \exu/alu_au/n35 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u724  (\exu/alu_au/n36 [45], \exu/alu_au/n34 [45], \exu/alu_au/n35 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u725  (\exu/alu_au/n36 [46], \exu/alu_au/n34 [46], \exu/alu_au/n35 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u726  (\exu/alu_au/n36 [47], \exu/alu_au/n34 [47], \exu/alu_au/n35 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u727  (\exu/alu_au/n36 [48], \exu/alu_au/n34 [48], \exu/alu_au/n35 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u728  (\exu/alu_au/n36 [49], \exu/alu_au/n34 [49], \exu/alu_au/n35 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u729  (\exu/alu_au/n36 [50], \exu/alu_au/n34 [50], \exu/alu_au/n35 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u73  (\exu/alu_data_mem_csr [24], \exu/alu_au/n54 [24], \exu/alu_au/n55 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u730  (\exu/alu_au/n36 [51], \exu/alu_au/n34 [51], \exu/alu_au/n35 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u731  (\exu/alu_au/n36 [52], \exu/alu_au/n34 [52], \exu/alu_au/n35 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u732  (\exu/alu_au/n36 [53], \exu/alu_au/n34 [53], \exu/alu_au/n35 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u733  (\exu/alu_au/n36 [54], \exu/alu_au/n34 [54], \exu/alu_au/n35 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u734  (\exu/alu_au/n36 [55], \exu/alu_au/n34 [55], \exu/alu_au/n35 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u735  (\exu/alu_au/n36 [56], \exu/alu_au/n34 [56], \exu/alu_au/n35 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u736  (\exu/alu_au/n36 [57], \exu/alu_au/n34 [57], \exu/alu_au/n35 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u737  (\exu/alu_au/n36 [58], \exu/alu_au/n34 [58], \exu/alu_au/n35 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u738  (\exu/alu_au/n36 [59], \exu/alu_au/n34 [59], \exu/alu_au/n35 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u739  (\exu/alu_au/n36 [60], \exu/alu_au/n34 [60], \exu/alu_au/n35 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u74  (\exu/alu_data_mem_csr [25], \exu/alu_au/n54 [25], \exu/alu_au/n55 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u740  (\exu/alu_au/n36 [61], \exu/alu_au/n34 [61], \exu/alu_au/n35 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u741  (\exu/alu_au/n36 [62], \exu/alu_au/n34 [62], \exu/alu_au/n35 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u742  (\exu/alu_au/n36 [63], \exu/alu_au/n34 [63], \exu/alu_au/n35 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(103)
  or \exu/alu_au/u743  (\exu/alu_au/n34 [1], \exu/alu_au/n32 [1], \exu/alu_au/n33 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u744  (\exu/alu_au/n34 [2], \exu/alu_au/n32 [2], \exu/alu_au/n33 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u745  (\exu/alu_au/n34 [3], \exu/alu_au/n32 [3], \exu/alu_au/n33 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u746  (\exu/alu_au/n34 [4], \exu/alu_au/n32 [4], \exu/alu_au/n33 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u747  (\exu/alu_au/n34 [5], \exu/alu_au/n32 [5], \exu/alu_au/n33 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u748  (\exu/alu_au/n34 [6], \exu/alu_au/n32 [6], \exu/alu_au/n33 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u749  (\exu/alu_au/n34 [7], \exu/alu_au/n32 [7], \exu/alu_au/n33 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u75  (\exu/alu_data_mem_csr [26], \exu/alu_au/n54 [26], \exu/alu_au/n55 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u750  (\exu/alu_au/n34 [8], \exu/alu_au/n32 [8], \exu/alu_au/n33 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u751  (\exu/alu_au/n34 [9], \exu/alu_au/n32 [9], \exu/alu_au/n33 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u752  (\exu/alu_au/n34 [10], \exu/alu_au/n32 [10], \exu/alu_au/n33 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u753  (\exu/alu_au/n34 [11], \exu/alu_au/n32 [11], \exu/alu_au/n33 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u754  (\exu/alu_au/n34 [12], \exu/alu_au/n32 [12], \exu/alu_au/n33 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u755  (\exu/alu_au/n34 [13], \exu/alu_au/n32 [13], \exu/alu_au/n33 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u756  (\exu/alu_au/n34 [14], \exu/alu_au/n32 [14], \exu/alu_au/n33 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u757  (\exu/alu_au/n34 [15], \exu/alu_au/n32 [15], \exu/alu_au/n33 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u758  (\exu/alu_au/n34 [16], \exu/alu_au/n32 [16], \exu/alu_au/n33 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u759  (\exu/alu_au/n34 [17], \exu/alu_au/n32 [17], \exu/alu_au/n33 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u76  (\exu/alu_data_mem_csr [27], \exu/alu_au/n54 [27], \exu/alu_au/n55 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u760  (\exu/alu_au/n34 [18], \exu/alu_au/n32 [18], \exu/alu_au/n33 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u761  (\exu/alu_au/n34 [19], \exu/alu_au/n32 [19], \exu/alu_au/n33 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u762  (\exu/alu_au/n34 [20], \exu/alu_au/n32 [20], \exu/alu_au/n33 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u763  (\exu/alu_au/n34 [21], \exu/alu_au/n32 [21], \exu/alu_au/n33 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u764  (\exu/alu_au/n34 [22], \exu/alu_au/n32 [22], \exu/alu_au/n33 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u765  (\exu/alu_au/n34 [23], \exu/alu_au/n32 [23], \exu/alu_au/n33 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u766  (\exu/alu_au/n34 [24], \exu/alu_au/n32 [24], \exu/alu_au/n33 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u767  (\exu/alu_au/n34 [25], \exu/alu_au/n32 [25], \exu/alu_au/n33 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u768  (\exu/alu_au/n34 [26], \exu/alu_au/n32 [26], \exu/alu_au/n33 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u769  (\exu/alu_au/n34 [27], \exu/alu_au/n32 [27], \exu/alu_au/n33 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u77  (\exu/alu_data_mem_csr [28], \exu/alu_au/n54 [28], \exu/alu_au/n55 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u770  (\exu/alu_au/n34 [28], \exu/alu_au/n32 [28], \exu/alu_au/n33 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u771  (\exu/alu_au/n34 [29], \exu/alu_au/n32 [29], \exu/alu_au/n33 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u772  (\exu/alu_au/n34 [30], \exu/alu_au/n32 [30], \exu/alu_au/n33 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u773  (\exu/alu_au/n34 [31], \exu/alu_au/n32 [31], \exu/alu_au/n33 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u774  (\exu/alu_au/n34 [32], \exu/alu_au/n32 [32], \exu/alu_au/n33 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u775  (\exu/alu_au/n34 [33], \exu/alu_au/n32 [33], \exu/alu_au/n33 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u776  (\exu/alu_au/n34 [34], \exu/alu_au/n32 [34], \exu/alu_au/n33 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u777  (\exu/alu_au/n34 [35], \exu/alu_au/n32 [35], \exu/alu_au/n33 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u778  (\exu/alu_au/n34 [36], \exu/alu_au/n32 [36], \exu/alu_au/n33 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u779  (\exu/alu_au/n34 [37], \exu/alu_au/n32 [37], \exu/alu_au/n33 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u78  (\exu/alu_data_mem_csr [29], \exu/alu_au/n54 [29], \exu/alu_au/n55 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u780  (\exu/alu_au/n34 [38], \exu/alu_au/n32 [38], \exu/alu_au/n33 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u781  (\exu/alu_au/n34 [39], \exu/alu_au/n32 [39], \exu/alu_au/n33 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u782  (\exu/alu_au/n34 [40], \exu/alu_au/n32 [40], \exu/alu_au/n33 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u783  (\exu/alu_au/n34 [41], \exu/alu_au/n32 [41], \exu/alu_au/n33 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u784  (\exu/alu_au/n34 [42], \exu/alu_au/n32 [42], \exu/alu_au/n33 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u785  (\exu/alu_au/n34 [43], \exu/alu_au/n32 [43], \exu/alu_au/n33 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u786  (\exu/alu_au/n34 [44], \exu/alu_au/n32 [44], \exu/alu_au/n33 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u787  (\exu/alu_au/n34 [45], \exu/alu_au/n32 [45], \exu/alu_au/n33 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u788  (\exu/alu_au/n34 [46], \exu/alu_au/n32 [46], \exu/alu_au/n33 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u789  (\exu/alu_au/n34 [47], \exu/alu_au/n32 [47], \exu/alu_au/n33 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u79  (\exu/alu_data_mem_csr [30], \exu/alu_au/n54 [30], \exu/alu_au/n55 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u790  (\exu/alu_au/n34 [48], \exu/alu_au/n32 [48], \exu/alu_au/n33 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u791  (\exu/alu_au/n34 [49], \exu/alu_au/n32 [49], \exu/alu_au/n33 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u792  (\exu/alu_au/n34 [50], \exu/alu_au/n32 [50], \exu/alu_au/n33 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u793  (\exu/alu_au/n34 [51], \exu/alu_au/n32 [51], \exu/alu_au/n33 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u794  (\exu/alu_au/n34 [52], \exu/alu_au/n32 [52], \exu/alu_au/n33 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u795  (\exu/alu_au/n34 [53], \exu/alu_au/n32 [53], \exu/alu_au/n33 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u796  (\exu/alu_au/n34 [54], \exu/alu_au/n32 [54], \exu/alu_au/n33 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u797  (\exu/alu_au/n34 [55], \exu/alu_au/n32 [55], \exu/alu_au/n33 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u798  (\exu/alu_au/n34 [56], \exu/alu_au/n32 [56], \exu/alu_au/n33 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u799  (\exu/alu_au/n34 [57], \exu/alu_au/n32 [57], \exu/alu_au/n33 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  not \exu/alu_au/u8  (\exu/alu_au/n4 , \exu/alu_au/alu_xor [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(72)
  or \exu/alu_au/u80  (\exu/alu_data_mem_csr [31], \exu/alu_au/n54 [31], \exu/alu_au/n55 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u800  (\exu/alu_au/n34 [58], \exu/alu_au/n32 [58], \exu/alu_au/n33 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u801  (\exu/alu_au/n34 [59], \exu/alu_au/n32 [59], \exu/alu_au/n33 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u802  (\exu/alu_au/n34 [60], \exu/alu_au/n32 [60], \exu/alu_au/n33 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u803  (\exu/alu_au/n34 [61], \exu/alu_au/n32 [61], \exu/alu_au/n33 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u804  (\exu/alu_au/n34 [62], \exu/alu_au/n32 [62], \exu/alu_au/n33 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u805  (\exu/alu_au/n34 [63], \exu/alu_au/n32 [63], \exu/alu_au/n33 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(102)
  or \exu/alu_au/u806  (\exu/alu_au/n32 [1], \exu/alu_au/n30 [1], \exu/alu_au/n31 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u807  (\exu/alu_au/n32 [2], \exu/alu_au/n30 [2], \exu/alu_au/n31 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u808  (\exu/alu_au/n32 [3], \exu/alu_au/n30 [3], \exu/alu_au/n31 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u809  (\exu/alu_au/n32 [4], \exu/alu_au/n30 [4], \exu/alu_au/n31 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u81  (\exu/alu_data_mem_csr [32], \exu/alu_au/n54 [32], \exu/alu_au/n55 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u810  (\exu/alu_au/n32 [5], \exu/alu_au/n30 [5], \exu/alu_au/n31 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u811  (\exu/alu_au/n32 [6], \exu/alu_au/n30 [6], \exu/alu_au/n31 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u812  (\exu/alu_au/n32 [7], \exu/alu_au/n30 [7], \exu/alu_au/n31 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u813  (\exu/alu_au/n32 [8], \exu/alu_au/n30 [8], \exu/alu_au/n31 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u814  (\exu/alu_au/n32 [9], \exu/alu_au/n30 [9], \exu/alu_au/n31 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u815  (\exu/alu_au/n32 [10], \exu/alu_au/n30 [10], \exu/alu_au/n31 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u816  (\exu/alu_au/n32 [11], \exu/alu_au/n30 [11], \exu/alu_au/n31 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u817  (\exu/alu_au/n32 [12], \exu/alu_au/n30 [12], \exu/alu_au/n31 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u818  (\exu/alu_au/n32 [13], \exu/alu_au/n30 [13], \exu/alu_au/n31 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u819  (\exu/alu_au/n32 [14], \exu/alu_au/n30 [14], \exu/alu_au/n31 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u82  (\exu/alu_data_mem_csr [33], \exu/alu_au/n54 [33], \exu/alu_au/n55 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u820  (\exu/alu_au/n32 [15], \exu/alu_au/n30 [15], \exu/alu_au/n31 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u821  (\exu/alu_au/n32 [16], \exu/alu_au/n30 [16], \exu/alu_au/n31 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u822  (\exu/alu_au/n32 [17], \exu/alu_au/n30 [17], \exu/alu_au/n31 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u823  (\exu/alu_au/n32 [18], \exu/alu_au/n30 [18], \exu/alu_au/n31 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u824  (\exu/alu_au/n32 [19], \exu/alu_au/n30 [19], \exu/alu_au/n31 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u825  (\exu/alu_au/n32 [20], \exu/alu_au/n30 [20], \exu/alu_au/n31 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u826  (\exu/alu_au/n32 [21], \exu/alu_au/n30 [21], \exu/alu_au/n31 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u827  (\exu/alu_au/n32 [22], \exu/alu_au/n30 [22], \exu/alu_au/n31 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u828  (\exu/alu_au/n32 [23], \exu/alu_au/n30 [23], \exu/alu_au/n31 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u829  (\exu/alu_au/n32 [24], \exu/alu_au/n30 [24], \exu/alu_au/n31 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u83  (\exu/alu_data_mem_csr [34], \exu/alu_au/n54 [34], \exu/alu_au/n55 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u830  (\exu/alu_au/n32 [25], \exu/alu_au/n30 [25], \exu/alu_au/n31 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u831  (\exu/alu_au/n32 [26], \exu/alu_au/n30 [26], \exu/alu_au/n31 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u832  (\exu/alu_au/n32 [27], \exu/alu_au/n30 [27], \exu/alu_au/n31 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u833  (\exu/alu_au/n32 [28], \exu/alu_au/n30 [28], \exu/alu_au/n31 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u834  (\exu/alu_au/n32 [29], \exu/alu_au/n30 [29], \exu/alu_au/n31 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u835  (\exu/alu_au/n32 [30], \exu/alu_au/n30 [30], \exu/alu_au/n31 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u836  (\exu/alu_au/n32 [31], \exu/alu_au/n30 [31], \exu/alu_au/n31 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u837  (\exu/alu_au/n32 [32], \exu/alu_au/n30 [32], \exu/alu_au/n31 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u838  (\exu/alu_au/n32 [33], \exu/alu_au/n30 [33], \exu/alu_au/n31 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u839  (\exu/alu_au/n32 [34], \exu/alu_au/n30 [34], \exu/alu_au/n31 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u84  (\exu/alu_data_mem_csr [35], \exu/alu_au/n54 [35], \exu/alu_au/n55 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u840  (\exu/alu_au/n32 [35], \exu/alu_au/n30 [35], \exu/alu_au/n31 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u841  (\exu/alu_au/n32 [36], \exu/alu_au/n30 [36], \exu/alu_au/n31 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u842  (\exu/alu_au/n32 [37], \exu/alu_au/n30 [37], \exu/alu_au/n31 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u843  (\exu/alu_au/n32 [38], \exu/alu_au/n30 [38], \exu/alu_au/n31 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u844  (\exu/alu_au/n32 [39], \exu/alu_au/n30 [39], \exu/alu_au/n31 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u845  (\exu/alu_au/n32 [40], \exu/alu_au/n30 [40], \exu/alu_au/n31 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u846  (\exu/alu_au/n32 [41], \exu/alu_au/n30 [41], \exu/alu_au/n31 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u847  (\exu/alu_au/n32 [42], \exu/alu_au/n30 [42], \exu/alu_au/n31 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u848  (\exu/alu_au/n32 [43], \exu/alu_au/n30 [43], \exu/alu_au/n31 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u849  (\exu/alu_au/n32 [44], \exu/alu_au/n30 [44], \exu/alu_au/n31 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u85  (\exu/alu_data_mem_csr [36], \exu/alu_au/n54 [36], \exu/alu_au/n55 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u850  (\exu/alu_au/n32 [45], \exu/alu_au/n30 [45], \exu/alu_au/n31 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u851  (\exu/alu_au/n32 [46], \exu/alu_au/n30 [46], \exu/alu_au/n31 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u852  (\exu/alu_au/n32 [47], \exu/alu_au/n30 [47], \exu/alu_au/n31 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u853  (\exu/alu_au/n32 [48], \exu/alu_au/n30 [48], \exu/alu_au/n31 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u854  (\exu/alu_au/n32 [49], \exu/alu_au/n30 [49], \exu/alu_au/n31 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u855  (\exu/alu_au/n32 [50], \exu/alu_au/n30 [50], \exu/alu_au/n31 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u856  (\exu/alu_au/n32 [51], \exu/alu_au/n30 [51], \exu/alu_au/n31 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u857  (\exu/alu_au/n32 [52], \exu/alu_au/n30 [52], \exu/alu_au/n31 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u858  (\exu/alu_au/n32 [53], \exu/alu_au/n30 [53], \exu/alu_au/n31 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u859  (\exu/alu_au/n32 [54], \exu/alu_au/n30 [54], \exu/alu_au/n31 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u86  (\exu/alu_data_mem_csr [37], \exu/alu_au/n54 [37], \exu/alu_au/n55 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u860  (\exu/alu_au/n32 [55], \exu/alu_au/n30 [55], \exu/alu_au/n31 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u861  (\exu/alu_au/n32 [56], \exu/alu_au/n30 [56], \exu/alu_au/n31 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u862  (\exu/alu_au/n32 [57], \exu/alu_au/n30 [57], \exu/alu_au/n31 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u863  (\exu/alu_au/n32 [58], \exu/alu_au/n30 [58], \exu/alu_au/n31 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u864  (\exu/alu_au/n32 [59], \exu/alu_au/n30 [59], \exu/alu_au/n31 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u865  (\exu/alu_au/n32 [60], \exu/alu_au/n30 [60], \exu/alu_au/n31 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u866  (\exu/alu_au/n32 [61], \exu/alu_au/n30 [61], \exu/alu_au/n31 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u867  (\exu/alu_au/n32 [62], \exu/alu_au/n30 [62], \exu/alu_au/n31 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u868  (\exu/alu_au/n32 [63], \exu/alu_au/n30 [63], \exu/alu_au/n31 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(101)
  or \exu/alu_au/u869  (\exu/alu_au/n30 [1], \exu/alu_au/n28 [1], \exu/alu_au/n29 [1]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u87  (\exu/alu_data_mem_csr [38], \exu/alu_au/n54 [38], \exu/alu_au/n55 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u870  (\exu/alu_au/n30 [2], \exu/alu_au/n28 [2], \exu/alu_au/n29 [2]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u871  (\exu/alu_au/n30 [3], \exu/alu_au/n28 [3], \exu/alu_au/n29 [3]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u872  (\exu/alu_au/n30 [4], \exu/alu_au/n28 [4], \exu/alu_au/n29 [4]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u873  (\exu/alu_au/n30 [5], \exu/alu_au/n28 [5], \exu/alu_au/n29 [5]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u874  (\exu/alu_au/n30 [6], \exu/alu_au/n28 [6], \exu/alu_au/n29 [6]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u875  (\exu/alu_au/n30 [7], \exu/alu_au/n28 [7], \exu/alu_au/n29 [7]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u876  (\exu/alu_au/n30 [8], \exu/alu_au/n28 [8], \exu/alu_au/n29 [8]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u877  (\exu/alu_au/n30 [9], \exu/alu_au/n28 [9], \exu/alu_au/n29 [9]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u878  (\exu/alu_au/n30 [10], \exu/alu_au/n28 [10], \exu/alu_au/n29 [10]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u879  (\exu/alu_au/n30 [11], \exu/alu_au/n28 [11], \exu/alu_au/n29 [11]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u88  (\exu/alu_data_mem_csr [39], \exu/alu_au/n54 [39], \exu/alu_au/n55 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u880  (\exu/alu_au/n30 [12], \exu/alu_au/n28 [12], \exu/alu_au/n29 [12]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u881  (\exu/alu_au/n30 [13], \exu/alu_au/n28 [13], \exu/alu_au/n29 [13]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u882  (\exu/alu_au/n30 [14], \exu/alu_au/n28 [14], \exu/alu_au/n29 [14]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u883  (\exu/alu_au/n30 [15], \exu/alu_au/n28 [15], \exu/alu_au/n29 [15]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u884  (\exu/alu_au/n30 [16], \exu/alu_au/n28 [16], \exu/alu_au/n29 [16]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u885  (\exu/alu_au/n30 [17], \exu/alu_au/n28 [17], \exu/alu_au/n29 [17]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u886  (\exu/alu_au/n30 [18], \exu/alu_au/n28 [18], \exu/alu_au/n29 [18]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u887  (\exu/alu_au/n30 [19], \exu/alu_au/n28 [19], \exu/alu_au/n29 [19]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u888  (\exu/alu_au/n30 [20], \exu/alu_au/n28 [20], \exu/alu_au/n29 [20]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u889  (\exu/alu_au/n30 [21], \exu/alu_au/n28 [21], \exu/alu_au/n29 [21]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u89  (\exu/alu_data_mem_csr [40], \exu/alu_au/n54 [40], \exu/alu_au/n55 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u890  (\exu/alu_au/n30 [22], \exu/alu_au/n28 [22], \exu/alu_au/n29 [22]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u891  (\exu/alu_au/n30 [23], \exu/alu_au/n28 [23], \exu/alu_au/n29 [23]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u892  (\exu/alu_au/n30 [24], \exu/alu_au/n28 [24], \exu/alu_au/n29 [24]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u893  (\exu/alu_au/n30 [25], \exu/alu_au/n28 [25], \exu/alu_au/n29 [25]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u894  (\exu/alu_au/n30 [26], \exu/alu_au/n28 [26], \exu/alu_au/n29 [26]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u895  (\exu/alu_au/n30 [27], \exu/alu_au/n28 [27], \exu/alu_au/n29 [27]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u896  (\exu/alu_au/n30 [28], \exu/alu_au/n28 [28], \exu/alu_au/n29 [28]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u897  (\exu/alu_au/n30 [29], \exu/alu_au/n28 [29], \exu/alu_au/n29 [29]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u898  (\exu/alu_au/n30 [30], \exu/alu_au/n28 [30], \exu/alu_au/n29 [30]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u899  (\exu/alu_au/n30 [31], \exu/alu_au/n28 [31], \exu/alu_au/n29 [31]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  and \exu/alu_au/u9  (\exu/alu_au/n6 , \exu/alu_au/n4 , \exu/alu_au/n5 );  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(72)
  or \exu/alu_au/u90  (\exu/alu_data_mem_csr [41], \exu/alu_au/n54 [41], \exu/alu_au/n55 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u900  (\exu/alu_au/n30 [32], \exu/alu_au/n28 [32], \exu/alu_au/n29 [32]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u901  (\exu/alu_au/n30 [33], \exu/alu_au/n28 [33], \exu/alu_au/n29 [33]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u902  (\exu/alu_au/n30 [34], \exu/alu_au/n28 [34], \exu/alu_au/n29 [34]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u903  (\exu/alu_au/n30 [35], \exu/alu_au/n28 [35], \exu/alu_au/n29 [35]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u904  (\exu/alu_au/n30 [36], \exu/alu_au/n28 [36], \exu/alu_au/n29 [36]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u905  (\exu/alu_au/n30 [37], \exu/alu_au/n28 [37], \exu/alu_au/n29 [37]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u906  (\exu/alu_au/n30 [38], \exu/alu_au/n28 [38], \exu/alu_au/n29 [38]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u907  (\exu/alu_au/n30 [39], \exu/alu_au/n28 [39], \exu/alu_au/n29 [39]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u908  (\exu/alu_au/n30 [40], \exu/alu_au/n28 [40], \exu/alu_au/n29 [40]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u909  (\exu/alu_au/n30 [41], \exu/alu_au/n28 [41], \exu/alu_au/n29 [41]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u91  (\exu/alu_data_mem_csr [42], \exu/alu_au/n54 [42], \exu/alu_au/n55 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u910  (\exu/alu_au/n30 [42], \exu/alu_au/n28 [42], \exu/alu_au/n29 [42]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u911  (\exu/alu_au/n30 [43], \exu/alu_au/n28 [43], \exu/alu_au/n29 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u912  (\exu/alu_au/n30 [44], \exu/alu_au/n28 [44], \exu/alu_au/n29 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u913  (\exu/alu_au/n30 [45], \exu/alu_au/n28 [45], \exu/alu_au/n29 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u914  (\exu/alu_au/n30 [46], \exu/alu_au/n28 [46], \exu/alu_au/n29 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u915  (\exu/alu_au/n30 [47], \exu/alu_au/n28 [47], \exu/alu_au/n29 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u916  (\exu/alu_au/n30 [48], \exu/alu_au/n28 [48], \exu/alu_au/n29 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u917  (\exu/alu_au/n30 [49], \exu/alu_au/n28 [49], \exu/alu_au/n29 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u918  (\exu/alu_au/n30 [50], \exu/alu_au/n28 [50], \exu/alu_au/n29 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u919  (\exu/alu_au/n30 [51], \exu/alu_au/n28 [51], \exu/alu_au/n29 [51]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u92  (\exu/alu_data_mem_csr [43], \exu/alu_au/n54 [43], \exu/alu_au/n55 [43]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u920  (\exu/alu_au/n30 [52], \exu/alu_au/n28 [52], \exu/alu_au/n29 [52]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u921  (\exu/alu_au/n30 [53], \exu/alu_au/n28 [53], \exu/alu_au/n29 [53]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u922  (\exu/alu_au/n30 [54], \exu/alu_au/n28 [54], \exu/alu_au/n29 [54]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u923  (\exu/alu_au/n30 [55], \exu/alu_au/n28 [55], \exu/alu_au/n29 [55]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u924  (\exu/alu_au/n30 [56], \exu/alu_au/n28 [56], \exu/alu_au/n29 [56]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u925  (\exu/alu_au/n30 [57], \exu/alu_au/n28 [57], \exu/alu_au/n29 [57]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u926  (\exu/alu_au/n30 [58], \exu/alu_au/n28 [58], \exu/alu_au/n29 [58]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u927  (\exu/alu_au/n30 [59], \exu/alu_au/n28 [59], \exu/alu_au/n29 [59]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u928  (\exu/alu_au/n30 [60], \exu/alu_au/n28 [60], \exu/alu_au/n29 [60]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u929  (\exu/alu_au/n30 [61], \exu/alu_au/n28 [61], \exu/alu_au/n29 [61]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u93  (\exu/alu_data_mem_csr [44], \exu/alu_au/n54 [44], \exu/alu_au/n55 [44]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u930  (\exu/alu_au/n30 [62], \exu/alu_au/n28 [62], \exu/alu_au/n29 [62]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u931  (\exu/alu_au/n30 [63], \exu/alu_au/n28 [63], \exu/alu_au/n29 [63]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(100)
  or \exu/alu_au/u94  (\exu/alu_data_mem_csr [45], \exu/alu_au/n54 [45], \exu/alu_au/n55 [45]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u95  (\exu/alu_data_mem_csr [46], \exu/alu_au/n54 [46], \exu/alu_au/n55 [46]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u96  (\exu/alu_data_mem_csr [47], \exu/alu_au/n54 [47], \exu/alu_au/n55 [47]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u97  (\exu/alu_data_mem_csr [48], \exu/alu_au/n54 [48], \exu/alu_au/n55 [48]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u98  (\exu/alu_data_mem_csr [49], \exu/alu_au/n54 [49], \exu/alu_au/n55 [49]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  or \exu/alu_au/u99  (\exu/alu_data_mem_csr [50], \exu/alu_au/n54 [50], \exu/alu_au/n55 [50]);  // ../../RTL/CPU/EX/ALU&AU/alu_au.v(116)
  not \exu/c_amo_mem01_inv  (\exu/c_amo_mem01_neg , \exu/c_amo_mem01 );
  not \exu/c_amo_mem0_inv  (\exu/c_amo_mem0_neg , \exu/c_amo_mem0 );
  not \exu/c_amo_mem1_inv  (\exu/c_amo_mem1_neg , \exu/c_amo_mem1 );
  not \exu/c_load_inv  (\exu/c_load_neg , \exu/c_load );
  not \exu/c_shift_inv  (\exu/c_shift_neg , \exu/c_shift );
  not \exu/c_store_inv  (\exu/c_store_neg , \exu/c_store );
  reg_sr_as_w1 \exu/csr_write_reg  (
    .clk(clk),
    .d(ex_csr_write),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_csr_write));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/ebreak_reg  (
    .clk(clk),
    .d(ex_ebreak),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ebreak));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ecall_reg  (
    .clk(clk),
    .d(ex_ecall),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ecall));  // ../../RTL/CPU/EX/exu.v(448)
  eq_w4 \exu/eq1  (
    .i0(\exu/main_state ),
    .i1(4'b0001),
    .o(\exu/c_shift ));  // ../../RTL/CPU/EX/exu.v(215)
  eq_w4 \exu/eq10  (
    .i0(\exu/main_state ),
    .i1(4'b1011),
    .o(\exu/c_amo_mem1 ));  // ../../RTL/CPU/EX/exu.v(264)
  eq_w4 \exu/eq11  (
    .i0(\exu/main_state ),
    .i1(4'b0011),
    .o(\exu/c_load_1 ));  // ../../RTL/CPU/EX/exu.v(272)
  eq_w3 \exu/eq12  (
    .i0({mod_priv[3],mod_priv[1:0]}),
    .i1(3'b011),
    .o(\exu/n148 ));  // ../../RTL/CPU/EX/exu.v(506)
  eq_w8 \exu/eq2  (
    .i0(\exu/shift_count ),
    .i1(8'b00000001),
    .o(\exu/n9 ));  // ../../RTL/CPU/EX/exu.v(215)
  eq_w4 \exu/eq3  (
    .i0(\exu/main_state ),
    .i1(4'b0000),
    .o(\exu/c_stb ));  // ../../RTL/CPU/EX/exu.v(235)
  eq_w4 \exu/eq4  (
    .i0(\exu/main_state ),
    .i1(4'b0010),
    .o(\exu/c_load ));  // ../../RTL/CPU/EX/exu.v(243)
  eq_w4 \exu/eq5  (
    .i0(\exu/main_state ),
    .i1(4'b0100),
    .o(\exu/c_store ));  // ../../RTL/CPU/EX/exu.v(246)
  eq_w4 \exu/eq6  (
    .i0(\exu/main_state ),
    .i1(4'b1000),
    .o(\exu/c_amo_mem0 ));  // ../../RTL/CPU/EX/exu.v(252)
  eq_w4 \exu/eq7  (
    .i0(\exu/main_state ),
    .i1(4'b1100),
    .o(\exu/c_fence ));  // ../../RTL/CPU/EX/exu.v(255)
  eq_w4 \exu/eq8  (
    .i0(\exu/main_state ),
    .i1(4'b1010),
    .o(\exu/n35 ));  // ../../RTL/CPU/EX/exu.v(258)
  eq_w4 \exu/eq9  (
    .i0(\exu/main_state ),
    .i1(4'b1001),
    .o(\exu/c_amo_mem01 ));  // ../../RTL/CPU/EX/exu.v(261)
  reg_sr_as_w1 \exu/gpr_write_reg  (
    .clk(clk),
    .d(ex_gpr_write),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_gpr_write));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/id_jmp_reg  (
    .clk(clk),
    .d(ex_jmp),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_jmp));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/id_system_reg  (
    .clk(clk),
    .d(ex_system),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_system));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ill_ins_reg  (
    .clk(clk),
    .d(ex_ill_ins),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ill_ins));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ins_acc_fault_reg  (
    .clk(clk),
    .d(ex_ins_acc_fault),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ins_acc_fault));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ins_addr_mis_reg  (
    .clk(clk),
    .d(ex_ins_addr_mis),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ins_addr_mis));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ins_page_fault_reg  (
    .clk(clk),
    .d(ex_ins_page_fault),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ins_page_fault));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/int_acc_reg  (
    .clk(clk),
    .d(ex_int_acc),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_int_acc));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ld_acc_fault_reg  (
    .clk(clk),
    .d(load_acc_fault),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ld_acc_fault));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ld_addr_mis_reg  (
    .clk(clk),
    .d(\exu/load_addr_mis ),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ld_addr_mis));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/ld_page_fault_reg  (
    .clk(clk),
    .d(load_page_fault),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_ld_page_fault));  // ../../RTL/CPU/EX/exu.v(448)
  eq_w2 \exu/lsu/eq0  (
    .i0(addr_ex[1:0]),
    .i1(2'b00),
    .o(\exu/lsu/n0 ));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  eq_w2 \exu/lsu/eq1  (
    .i0(addr_ex[1:0]),
    .i1(2'b01),
    .o(\exu/lsu/n2 ));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  eq_w2 \exu/lsu/eq2  (
    .i0(addr_ex[1:0]),
    .i1(2'b10),
    .o(\exu/lsu/n5 ));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  eq_w2 \exu/lsu/eq3  (
    .i0(addr_ex[1:0]),
    .i1(2'b11),
    .o(\exu/lsu/n8 ));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux0_b0  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [0]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b1  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [1]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b10  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [10]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b11  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [11]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b12  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [12]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b13  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [13]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b14  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [14]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b15  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [15]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b16  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [16]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b17  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [17]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b18  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [18]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b19  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [19]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b2  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [2]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b20  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [20]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b21  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [21]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b22  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [22]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b23  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [23]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b24  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [24]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b25  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [25]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b26  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [26]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b27  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [27]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b28  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [28]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b29  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [29]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b3  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [3]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b30  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [30]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b31  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [31]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b32  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [32]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b33  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [33]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b34  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [34]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b35  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [35]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b36  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [36]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b37  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [37]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b38  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [38]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b39  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [39]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b4  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [4]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b40  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [40]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b41  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [41]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b42  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [42]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b43  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [43]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b44  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [44]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b45  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [45]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b46  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [46]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b47  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [47]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b48  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [48]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [48]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b49  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [49]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [49]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b5  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [5]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b50  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [50]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [50]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b51  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [51]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [51]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b52  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [52]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [52]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b53  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [53]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [53]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b54  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [54]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [54]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b55  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [55]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [55]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b56  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [56]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [56]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b57  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [57]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [57]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b58  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [58]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [58]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b59  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [59]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [59]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b6  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [6]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b60  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [60]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [60]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b61  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [61]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [61]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b62  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [62]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [62]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b63  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [63]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [63]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b7  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [7]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b8  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [8]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux0_b9  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [9]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n1 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(32)
  binary_mux_s1_w1 \exu/lsu/mux10_b0  (
    .i0(1'b0),
    .i1(uncache_data[16]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b1  (
    .i0(1'b0),
    .i1(uncache_data[17]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b10  (
    .i0(1'b0),
    .i1(uncache_data[26]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b11  (
    .i0(1'b0),
    .i1(uncache_data[27]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b12  (
    .i0(1'b0),
    .i1(uncache_data[28]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b13  (
    .i0(1'b0),
    .i1(uncache_data[29]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b14  (
    .i0(1'b0),
    .i1(uncache_data[30]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b15  (
    .i0(1'b0),
    .i1(uncache_data[31]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b16  (
    .i0(1'b0),
    .i1(uncache_data[32]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b17  (
    .i0(1'b0),
    .i1(uncache_data[33]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b18  (
    .i0(1'b0),
    .i1(uncache_data[34]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b19  (
    .i0(1'b0),
    .i1(uncache_data[35]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b2  (
    .i0(1'b0),
    .i1(uncache_data[18]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b20  (
    .i0(1'b0),
    .i1(uncache_data[36]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b21  (
    .i0(1'b0),
    .i1(uncache_data[37]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b22  (
    .i0(1'b0),
    .i1(uncache_data[38]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b23  (
    .i0(1'b0),
    .i1(uncache_data[39]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b24  (
    .i0(1'b0),
    .i1(uncache_data[40]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b25  (
    .i0(1'b0),
    .i1(uncache_data[41]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b26  (
    .i0(1'b0),
    .i1(uncache_data[42]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b27  (
    .i0(1'b0),
    .i1(uncache_data[43]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b28  (
    .i0(1'b0),
    .i1(uncache_data[44]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b29  (
    .i0(1'b0),
    .i1(uncache_data[45]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b3  (
    .i0(1'b0),
    .i1(uncache_data[19]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b30  (
    .i0(1'b0),
    .i1(uncache_data[46]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b31  (
    .i0(1'b0),
    .i1(uncache_data[47]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b32  (
    .i0(1'b0),
    .i1(uncache_data[48]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b33  (
    .i0(1'b0),
    .i1(uncache_data[49]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b34  (
    .i0(1'b0),
    .i1(uncache_data[50]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b35  (
    .i0(1'b0),
    .i1(uncache_data[51]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b36  (
    .i0(1'b0),
    .i1(uncache_data[52]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b37  (
    .i0(1'b0),
    .i1(uncache_data[53]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b38  (
    .i0(1'b0),
    .i1(uncache_data[54]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b39  (
    .i0(1'b0),
    .i1(uncache_data[55]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b4  (
    .i0(1'b0),
    .i1(uncache_data[20]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b40  (
    .i0(1'b0),
    .i1(uncache_data[56]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b41  (
    .i0(1'b0),
    .i1(uncache_data[57]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b42  (
    .i0(1'b0),
    .i1(uncache_data[58]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b43  (
    .i0(1'b0),
    .i1(uncache_data[59]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b44  (
    .i0(1'b0),
    .i1(uncache_data[60]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b45  (
    .i0(1'b0),
    .i1(uncache_data[61]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b46  (
    .i0(1'b0),
    .i1(uncache_data[62]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b47  (
    .i0(1'b0),
    .i1(uncache_data[63]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b5  (
    .i0(1'b0),
    .i1(uncache_data[21]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b6  (
    .i0(1'b0),
    .i1(uncache_data[22]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b7  (
    .i0(1'b0),
    .i1(uncache_data[23]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b8  (
    .i0(1'b0),
    .i1(uncache_data[24]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux10_b9  (
    .i0(1'b0),
    .i1(uncache_data[25]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n25 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  binary_mux_s1_w1 \exu/lsu/mux11_b0  (
    .i0(1'b0),
    .i1(uncache_data[24]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b1  (
    .i0(1'b0),
    .i1(uncache_data[25]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b10  (
    .i0(1'b0),
    .i1(uncache_data[34]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b11  (
    .i0(1'b0),
    .i1(uncache_data[35]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b12  (
    .i0(1'b0),
    .i1(uncache_data[36]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b13  (
    .i0(1'b0),
    .i1(uncache_data[37]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b14  (
    .i0(1'b0),
    .i1(uncache_data[38]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b15  (
    .i0(1'b0),
    .i1(uncache_data[39]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b16  (
    .i0(1'b0),
    .i1(uncache_data[40]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b17  (
    .i0(1'b0),
    .i1(uncache_data[41]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b18  (
    .i0(1'b0),
    .i1(uncache_data[42]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b19  (
    .i0(1'b0),
    .i1(uncache_data[43]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b2  (
    .i0(1'b0),
    .i1(uncache_data[26]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b20  (
    .i0(1'b0),
    .i1(uncache_data[44]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b21  (
    .i0(1'b0),
    .i1(uncache_data[45]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b22  (
    .i0(1'b0),
    .i1(uncache_data[46]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b23  (
    .i0(1'b0),
    .i1(uncache_data[47]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b24  (
    .i0(1'b0),
    .i1(uncache_data[48]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b25  (
    .i0(1'b0),
    .i1(uncache_data[49]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b26  (
    .i0(1'b0),
    .i1(uncache_data[50]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b27  (
    .i0(1'b0),
    .i1(uncache_data[51]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b28  (
    .i0(1'b0),
    .i1(uncache_data[52]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b29  (
    .i0(1'b0),
    .i1(uncache_data[53]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b3  (
    .i0(1'b0),
    .i1(uncache_data[27]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b30  (
    .i0(1'b0),
    .i1(uncache_data[54]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b31  (
    .i0(1'b0),
    .i1(uncache_data[55]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b32  (
    .i0(1'b0),
    .i1(uncache_data[56]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b33  (
    .i0(1'b0),
    .i1(uncache_data[57]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b34  (
    .i0(1'b0),
    .i1(uncache_data[58]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b35  (
    .i0(1'b0),
    .i1(uncache_data[59]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b36  (
    .i0(1'b0),
    .i1(uncache_data[60]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b37  (
    .i0(1'b0),
    .i1(uncache_data[61]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b38  (
    .i0(1'b0),
    .i1(uncache_data[62]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b39  (
    .i0(1'b0),
    .i1(uncache_data[63]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b4  (
    .i0(1'b0),
    .i1(uncache_data[28]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b5  (
    .i0(1'b0),
    .i1(uncache_data[29]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b6  (
    .i0(1'b0),
    .i1(uncache_data[30]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b7  (
    .i0(1'b0),
    .i1(uncache_data[31]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b8  (
    .i0(1'b0),
    .i1(uncache_data[32]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux11_b9  (
    .i0(1'b0),
    .i1(uncache_data[33]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n27 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  binary_mux_s1_w1 \exu/lsu/mux16_b0  (
    .i0(1'b0),
    .i1(data_read[0]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b1  (
    .i0(1'b0),
    .i1(data_read[1]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b10  (
    .i0(1'b0),
    .i1(data_read[10]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b11  (
    .i0(1'b0),
    .i1(data_read[11]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b12  (
    .i0(1'b0),
    .i1(data_read[12]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b13  (
    .i0(1'b0),
    .i1(data_read[13]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b14  (
    .i0(1'b0),
    .i1(data_read[14]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b15  (
    .i0(1'b0),
    .i1(data_read[15]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b16  (
    .i0(1'b0),
    .i1(data_read[16]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b17  (
    .i0(1'b0),
    .i1(data_read[17]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b18  (
    .i0(1'b0),
    .i1(data_read[18]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b19  (
    .i0(1'b0),
    .i1(data_read[19]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b2  (
    .i0(1'b0),
    .i1(data_read[2]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b20  (
    .i0(1'b0),
    .i1(data_read[20]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b21  (
    .i0(1'b0),
    .i1(data_read[21]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b22  (
    .i0(1'b0),
    .i1(data_read[22]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b23  (
    .i0(1'b0),
    .i1(data_read[23]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b24  (
    .i0(1'b0),
    .i1(data_read[24]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b25  (
    .i0(1'b0),
    .i1(data_read[25]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b26  (
    .i0(1'b0),
    .i1(data_read[26]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b27  (
    .i0(1'b0),
    .i1(data_read[27]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b28  (
    .i0(1'b0),
    .i1(data_read[28]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b29  (
    .i0(1'b0),
    .i1(data_read[29]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b3  (
    .i0(1'b0),
    .i1(data_read[3]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b30  (
    .i0(1'b0),
    .i1(data_read[30]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b31  (
    .i0(1'b0),
    .i1(data_read[31]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b32  (
    .i0(1'b0),
    .i1(data_read[32]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b33  (
    .i0(1'b0),
    .i1(data_read[33]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b34  (
    .i0(1'b0),
    .i1(data_read[34]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b35  (
    .i0(1'b0),
    .i1(data_read[35]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b36  (
    .i0(1'b0),
    .i1(data_read[36]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b37  (
    .i0(1'b0),
    .i1(data_read[37]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b38  (
    .i0(1'b0),
    .i1(data_read[38]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b39  (
    .i0(1'b0),
    .i1(data_read[39]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b4  (
    .i0(1'b0),
    .i1(data_read[4]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b40  (
    .i0(1'b0),
    .i1(data_read[40]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b41  (
    .i0(1'b0),
    .i1(data_read[41]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b42  (
    .i0(1'b0),
    .i1(data_read[42]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b43  (
    .i0(1'b0),
    .i1(data_read[43]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b44  (
    .i0(1'b0),
    .i1(data_read[44]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b45  (
    .i0(1'b0),
    .i1(data_read[45]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b46  (
    .i0(1'b0),
    .i1(data_read[46]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b47  (
    .i0(1'b0),
    .i1(data_read[47]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b48  (
    .i0(1'b0),
    .i1(data_read[48]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [48]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b49  (
    .i0(1'b0),
    .i1(data_read[49]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [49]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b5  (
    .i0(1'b0),
    .i1(data_read[5]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b50  (
    .i0(1'b0),
    .i1(data_read[50]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [50]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b51  (
    .i0(1'b0),
    .i1(data_read[51]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [51]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b52  (
    .i0(1'b0),
    .i1(data_read[52]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [52]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b53  (
    .i0(1'b0),
    .i1(data_read[53]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [53]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b54  (
    .i0(1'b0),
    .i1(data_read[54]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [54]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b55  (
    .i0(1'b0),
    .i1(data_read[55]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [55]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b6  (
    .i0(1'b0),
    .i1(data_read[6]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b7  (
    .i0(1'b0),
    .i1(data_read[7]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b8  (
    .i0(1'b0),
    .i1(data_read[8]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux16_b9  (
    .i0(1'b0),
    .i1(data_read[9]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n36 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(51)
  binary_mux_s1_w1 \exu/lsu/mux17_b0  (
    .i0(1'b0),
    .i1(data_read[8]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b1  (
    .i0(1'b0),
    .i1(data_read[9]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b10  (
    .i0(1'b0),
    .i1(data_read[18]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b11  (
    .i0(1'b0),
    .i1(data_read[19]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b12  (
    .i0(1'b0),
    .i1(data_read[20]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b13  (
    .i0(1'b0),
    .i1(data_read[21]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b14  (
    .i0(1'b0),
    .i1(data_read[22]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b15  (
    .i0(1'b0),
    .i1(data_read[23]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b16  (
    .i0(1'b0),
    .i1(data_read[24]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b17  (
    .i0(1'b0),
    .i1(data_read[25]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b18  (
    .i0(1'b0),
    .i1(data_read[26]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b19  (
    .i0(1'b0),
    .i1(data_read[27]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b2  (
    .i0(1'b0),
    .i1(data_read[10]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b20  (
    .i0(1'b0),
    .i1(data_read[28]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b21  (
    .i0(1'b0),
    .i1(data_read[29]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b22  (
    .i0(1'b0),
    .i1(data_read[30]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b23  (
    .i0(1'b0),
    .i1(data_read[31]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b24  (
    .i0(1'b0),
    .i1(data_read[32]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b25  (
    .i0(1'b0),
    .i1(data_read[33]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b26  (
    .i0(1'b0),
    .i1(data_read[34]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b27  (
    .i0(1'b0),
    .i1(data_read[35]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b28  (
    .i0(1'b0),
    .i1(data_read[36]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b29  (
    .i0(1'b0),
    .i1(data_read[37]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b3  (
    .i0(1'b0),
    .i1(data_read[11]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b30  (
    .i0(1'b0),
    .i1(data_read[38]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b31  (
    .i0(1'b0),
    .i1(data_read[39]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b32  (
    .i0(1'b0),
    .i1(data_read[40]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b33  (
    .i0(1'b0),
    .i1(data_read[41]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b34  (
    .i0(1'b0),
    .i1(data_read[42]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b35  (
    .i0(1'b0),
    .i1(data_read[43]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b36  (
    .i0(1'b0),
    .i1(data_read[44]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b37  (
    .i0(1'b0),
    .i1(data_read[45]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b38  (
    .i0(1'b0),
    .i1(data_read[46]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b39  (
    .i0(1'b0),
    .i1(data_read[47]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b4  (
    .i0(1'b0),
    .i1(data_read[12]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b40  (
    .i0(1'b0),
    .i1(data_read[48]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b41  (
    .i0(1'b0),
    .i1(data_read[49]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b42  (
    .i0(1'b0),
    .i1(data_read[50]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b43  (
    .i0(1'b0),
    .i1(data_read[51]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b44  (
    .i0(1'b0),
    .i1(data_read[52]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b45  (
    .i0(1'b0),
    .i1(data_read[53]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b46  (
    .i0(1'b0),
    .i1(data_read[54]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b47  (
    .i0(1'b0),
    .i1(data_read[55]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b48  (
    .i0(1'b0),
    .i1(data_read[56]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [48]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b49  (
    .i0(1'b0),
    .i1(data_read[57]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [49]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b5  (
    .i0(1'b0),
    .i1(data_read[13]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b50  (
    .i0(1'b0),
    .i1(data_read[58]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [50]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b51  (
    .i0(1'b0),
    .i1(data_read[59]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [51]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b52  (
    .i0(1'b0),
    .i1(data_read[60]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [52]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b53  (
    .i0(1'b0),
    .i1(data_read[61]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [53]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b54  (
    .i0(1'b0),
    .i1(data_read[62]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [54]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b55  (
    .i0(1'b0),
    .i1(data_read[63]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [55]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b6  (
    .i0(1'b0),
    .i1(data_read[14]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b7  (
    .i0(1'b0),
    .i1(data_read[15]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b8  (
    .i0(1'b0),
    .i1(data_read[16]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux17_b9  (
    .i0(1'b0),
    .i1(data_read[17]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n37 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  binary_mux_s1_w1 \exu/lsu/mux18_b0  (
    .i0(1'b0),
    .i1(data_read[16]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b1  (
    .i0(1'b0),
    .i1(data_read[17]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b10  (
    .i0(1'b0),
    .i1(data_read[26]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b11  (
    .i0(1'b0),
    .i1(data_read[27]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b12  (
    .i0(1'b0),
    .i1(data_read[28]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b13  (
    .i0(1'b0),
    .i1(data_read[29]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b14  (
    .i0(1'b0),
    .i1(data_read[30]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b15  (
    .i0(1'b0),
    .i1(data_read[31]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b16  (
    .i0(1'b0),
    .i1(data_read[32]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b17  (
    .i0(1'b0),
    .i1(data_read[33]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b18  (
    .i0(1'b0),
    .i1(data_read[34]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b19  (
    .i0(1'b0),
    .i1(data_read[35]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b2  (
    .i0(1'b0),
    .i1(data_read[18]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b20  (
    .i0(1'b0),
    .i1(data_read[36]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b21  (
    .i0(1'b0),
    .i1(data_read[37]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b22  (
    .i0(1'b0),
    .i1(data_read[38]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b23  (
    .i0(1'b0),
    .i1(data_read[39]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b24  (
    .i0(1'b0),
    .i1(data_read[40]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b25  (
    .i0(1'b0),
    .i1(data_read[41]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b26  (
    .i0(1'b0),
    .i1(data_read[42]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b27  (
    .i0(1'b0),
    .i1(data_read[43]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b28  (
    .i0(1'b0),
    .i1(data_read[44]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b29  (
    .i0(1'b0),
    .i1(data_read[45]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b3  (
    .i0(1'b0),
    .i1(data_read[19]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b30  (
    .i0(1'b0),
    .i1(data_read[46]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b31  (
    .i0(1'b0),
    .i1(data_read[47]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b32  (
    .i0(1'b0),
    .i1(data_read[48]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b33  (
    .i0(1'b0),
    .i1(data_read[49]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b34  (
    .i0(1'b0),
    .i1(data_read[50]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b35  (
    .i0(1'b0),
    .i1(data_read[51]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b36  (
    .i0(1'b0),
    .i1(data_read[52]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b37  (
    .i0(1'b0),
    .i1(data_read[53]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b38  (
    .i0(1'b0),
    .i1(data_read[54]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b39  (
    .i0(1'b0),
    .i1(data_read[55]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b4  (
    .i0(1'b0),
    .i1(data_read[20]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b40  (
    .i0(1'b0),
    .i1(data_read[56]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b41  (
    .i0(1'b0),
    .i1(data_read[57]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b42  (
    .i0(1'b0),
    .i1(data_read[58]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b43  (
    .i0(1'b0),
    .i1(data_read[59]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b44  (
    .i0(1'b0),
    .i1(data_read[60]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b45  (
    .i0(1'b0),
    .i1(data_read[61]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b46  (
    .i0(1'b0),
    .i1(data_read[62]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b47  (
    .i0(1'b0),
    .i1(data_read[63]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b5  (
    .i0(1'b0),
    .i1(data_read[21]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b6  (
    .i0(1'b0),
    .i1(data_read[22]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b7  (
    .i0(1'b0),
    .i1(data_read[23]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b8  (
    .i0(1'b0),
    .i1(data_read[24]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux18_b9  (
    .i0(1'b0),
    .i1(data_read[25]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n39 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  binary_mux_s1_w1 \exu/lsu/mux19_b0  (
    .i0(1'b0),
    .i1(data_read[24]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b1  (
    .i0(1'b0),
    .i1(data_read[25]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b10  (
    .i0(1'b0),
    .i1(data_read[34]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b11  (
    .i0(1'b0),
    .i1(data_read[35]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b12  (
    .i0(1'b0),
    .i1(data_read[36]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b13  (
    .i0(1'b0),
    .i1(data_read[37]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b14  (
    .i0(1'b0),
    .i1(data_read[38]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b15  (
    .i0(1'b0),
    .i1(data_read[39]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b16  (
    .i0(1'b0),
    .i1(data_read[40]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b17  (
    .i0(1'b0),
    .i1(data_read[41]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b18  (
    .i0(1'b0),
    .i1(data_read[42]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b19  (
    .i0(1'b0),
    .i1(data_read[43]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b2  (
    .i0(1'b0),
    .i1(data_read[26]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b20  (
    .i0(1'b0),
    .i1(data_read[44]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b21  (
    .i0(1'b0),
    .i1(data_read[45]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b22  (
    .i0(1'b0),
    .i1(data_read[46]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b23  (
    .i0(1'b0),
    .i1(data_read[47]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b24  (
    .i0(1'b0),
    .i1(data_read[48]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b25  (
    .i0(1'b0),
    .i1(data_read[49]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b26  (
    .i0(1'b0),
    .i1(data_read[50]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b27  (
    .i0(1'b0),
    .i1(data_read[51]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b28  (
    .i0(1'b0),
    .i1(data_read[52]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b29  (
    .i0(1'b0),
    .i1(data_read[53]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b3  (
    .i0(1'b0),
    .i1(data_read[27]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b30  (
    .i0(1'b0),
    .i1(data_read[54]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b31  (
    .i0(1'b0),
    .i1(data_read[55]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b32  (
    .i0(1'b0),
    .i1(data_read[56]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b33  (
    .i0(1'b0),
    .i1(data_read[57]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b34  (
    .i0(1'b0),
    .i1(data_read[58]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b35  (
    .i0(1'b0),
    .i1(data_read[59]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b36  (
    .i0(1'b0),
    .i1(data_read[60]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b37  (
    .i0(1'b0),
    .i1(data_read[61]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b38  (
    .i0(1'b0),
    .i1(data_read[62]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b39  (
    .i0(1'b0),
    .i1(data_read[63]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b4  (
    .i0(1'b0),
    .i1(data_read[28]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b5  (
    .i0(1'b0),
    .i1(data_read[29]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b6  (
    .i0(1'b0),
    .i1(data_read[30]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b7  (
    .i0(1'b0),
    .i1(data_read[31]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b8  (
    .i0(1'b0),
    .i1(data_read[32]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux19_b9  (
    .i0(1'b0),
    .i1(data_read[33]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n41 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  binary_mux_s1_w1 \exu/lsu/mux1_b10  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [2]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b11  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [3]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b12  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [4]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b13  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [5]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b14  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [6]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b15  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [7]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b16  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [8]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b17  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [9]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b18  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [10]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b19  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [11]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b20  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [12]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b21  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [13]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b22  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [14]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b23  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [15]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b24  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [16]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b25  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [17]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b26  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [18]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b27  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [19]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b28  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [20]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b29  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [21]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b30  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [22]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b31  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [23]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b32  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [24]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b33  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [25]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b34  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [26]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b35  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [27]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b36  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [28]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b37  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [29]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b38  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [30]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b39  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [31]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b40  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [32]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b41  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [33]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b42  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [34]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b43  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [35]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b44  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [36]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b45  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [37]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b46  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [38]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b47  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [39]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b48  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [40]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [48]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b49  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [41]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [49]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b50  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [42]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [50]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b51  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [43]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [51]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b52  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [44]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [52]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b53  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [45]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [53]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b54  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [46]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [54]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b55  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [47]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [55]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b56  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [48]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [56]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b57  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [49]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [57]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b58  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [50]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [58]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b59  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [51]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [59]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b60  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [52]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [60]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b61  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [53]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [61]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b62  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [54]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [62]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b63  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [55]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [63]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b8  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [0]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux1_b9  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [1]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n3 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  binary_mux_s1_w1 \exu/lsu/mux24_b0  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [0]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n52 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(61)
  binary_mux_s1_w1 \exu/lsu/mux24_b1  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [1]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n52 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(61)
  binary_mux_s1_w1 \exu/lsu/mux24_b10  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [7]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n52 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(61)
  binary_mux_s1_w1 \exu/lsu/mux24_b2  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [2]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n52 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(61)
  binary_mux_s1_w1 \exu/lsu/mux24_b3  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [3]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n52 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(61)
  binary_mux_s1_w1 \exu/lsu/mux24_b4  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [4]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n52 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(61)
  binary_mux_s1_w1 \exu/lsu/mux24_b5  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [5]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n52 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(61)
  binary_mux_s1_w1 \exu/lsu/mux24_b6  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [6]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n52 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(61)
  binary_mux_s1_w1 \exu/lsu/mux25_b0  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [0]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b1  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [1]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b10  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [10]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b11  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [11]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b12  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [12]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b13  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [13]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b14  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [14]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b15  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [15]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b2  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [2]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b3  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [3]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b4  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [4]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b5  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [5]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b6  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [6]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b7  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [7]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b8  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [8]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux25_b9  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [9]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n54 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  binary_mux_s1_w1 \exu/lsu/mux26_b0  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [0]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b1  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [1]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b10  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [10]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b11  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [11]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b12  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [12]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b13  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [13]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b14  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [14]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b15  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [15]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b16  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [16]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b17  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [17]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b18  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [18]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b19  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [19]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b2  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [2]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b20  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [20]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b21  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [21]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b22  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [22]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b23  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [23]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b24  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [24]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b25  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [25]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b26  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [26]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b27  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [27]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b28  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [28]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b29  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [29]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b3  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [3]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b30  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [30]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b31  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [31]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b4  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [4]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b5  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [5]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b6  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [6]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b7  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [7]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b8  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [8]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux26_b9  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [9]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n57 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  binary_mux_s1_w1 \exu/lsu/mux27_b0  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [0]),
    .sel(unsign),
    .o(\exu/lsu/n59 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b1  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [1]),
    .sel(unsign),
    .o(\exu/lsu/n59 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b10  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [10]),
    .sel(unsign),
    .o(\exu/lsu/n59 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b11  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [11]),
    .sel(unsign),
    .o(\exu/lsu/n59 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b12  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [12]),
    .sel(unsign),
    .o(\exu/lsu/n59 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b13  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [13]),
    .sel(unsign),
    .o(\exu/lsu/n59 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b14  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [14]),
    .sel(unsign),
    .o(\exu/lsu/n59 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b15  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [15]),
    .sel(unsign),
    .o(\exu/lsu/n59 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b16  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [16]),
    .sel(unsign),
    .o(\exu/lsu/n59 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b17  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [17]),
    .sel(unsign),
    .o(\exu/lsu/n59 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b18  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [18]),
    .sel(unsign),
    .o(\exu/lsu/n59 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b19  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [19]),
    .sel(unsign),
    .o(\exu/lsu/n59 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b2  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [2]),
    .sel(unsign),
    .o(\exu/lsu/n59 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b20  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [20]),
    .sel(unsign),
    .o(\exu/lsu/n59 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b21  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [21]),
    .sel(unsign),
    .o(\exu/lsu/n59 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b22  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [22]),
    .sel(unsign),
    .o(\exu/lsu/n59 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b23  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [23]),
    .sel(unsign),
    .o(\exu/lsu/n59 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b24  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [24]),
    .sel(unsign),
    .o(\exu/lsu/n59 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b25  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [25]),
    .sel(unsign),
    .o(\exu/lsu/n59 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b26  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [26]),
    .sel(unsign),
    .o(\exu/lsu/n59 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b27  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [27]),
    .sel(unsign),
    .o(\exu/lsu/n59 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b28  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [28]),
    .sel(unsign),
    .o(\exu/lsu/n59 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b29  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [29]),
    .sel(unsign),
    .o(\exu/lsu/n59 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b3  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [3]),
    .sel(unsign),
    .o(\exu/lsu/n59 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b30  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [30]),
    .sel(unsign),
    .o(\exu/lsu/n59 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b31  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [31]),
    .sel(unsign),
    .o(\exu/lsu/n59 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b32  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [32]),
    .sel(unsign),
    .o(\exu/lsu/n59 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b33  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [33]),
    .sel(unsign),
    .o(\exu/lsu/n59 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b34  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [34]),
    .sel(unsign),
    .o(\exu/lsu/n59 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b35  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [35]),
    .sel(unsign),
    .o(\exu/lsu/n59 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b36  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [36]),
    .sel(unsign),
    .o(\exu/lsu/n59 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b37  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [37]),
    .sel(unsign),
    .o(\exu/lsu/n59 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b38  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [38]),
    .sel(unsign),
    .o(\exu/lsu/n59 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b39  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [39]),
    .sel(unsign),
    .o(\exu/lsu/n59 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b4  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [4]),
    .sel(unsign),
    .o(\exu/lsu/n59 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b40  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [40]),
    .sel(unsign),
    .o(\exu/lsu/n59 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b41  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [41]),
    .sel(unsign),
    .o(\exu/lsu/n59 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b42  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [42]),
    .sel(unsign),
    .o(\exu/lsu/n59 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b43  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [43]),
    .sel(unsign),
    .o(\exu/lsu/n59 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b44  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [44]),
    .sel(unsign),
    .o(\exu/lsu/n59 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b45  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [45]),
    .sel(unsign),
    .o(\exu/lsu/n59 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b46  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [46]),
    .sel(unsign),
    .o(\exu/lsu/n59 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b47  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [47]),
    .sel(unsign),
    .o(\exu/lsu/n59 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b48  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [48]),
    .sel(unsign),
    .o(\exu/lsu/n59 [48]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b49  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [49]),
    .sel(unsign),
    .o(\exu/lsu/n59 [49]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b5  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [5]),
    .sel(unsign),
    .o(\exu/lsu/n59 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b50  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [50]),
    .sel(unsign),
    .o(\exu/lsu/n59 [50]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b51  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [51]),
    .sel(unsign),
    .o(\exu/lsu/n59 [51]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b52  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [52]),
    .sel(unsign),
    .o(\exu/lsu/n59 [52]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b53  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [53]),
    .sel(unsign),
    .o(\exu/lsu/n59 [53]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b54  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [54]),
    .sel(unsign),
    .o(\exu/lsu/n59 [54]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b55  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_uncache_shift [55]),
    .sel(unsign),
    .o(\exu/lsu/n59 [55]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  AL_MUX \exu/lsu/mux27_b56  (
    .i0(1'b0),
    .i1(uncache_data[56]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [56]));
  and \exu/lsu/mux27_b56_sel_is_3  (\exu/lsu/mux27_b56_sel_is_3_o , unsign, \exu/lsu/n0 );
  AL_MUX \exu/lsu/mux27_b57  (
    .i0(1'b0),
    .i1(uncache_data[57]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [57]));
  AL_MUX \exu/lsu/mux27_b58  (
    .i0(1'b0),
    .i1(uncache_data[58]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [58]));
  AL_MUX \exu/lsu/mux27_b59  (
    .i0(1'b0),
    .i1(uncache_data[59]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [59]));
  binary_mux_s1_w1 \exu/lsu/mux27_b6  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [6]),
    .sel(unsign),
    .o(\exu/lsu/n59 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  AL_MUX \exu/lsu/mux27_b60  (
    .i0(1'b0),
    .i1(uncache_data[60]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [60]));
  AL_MUX \exu/lsu/mux27_b61  (
    .i0(1'b0),
    .i1(uncache_data[61]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [61]));
  AL_MUX \exu/lsu/mux27_b62  (
    .i0(1'b0),
    .i1(uncache_data[62]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [62]));
  AL_MUX \exu/lsu/mux27_b63  (
    .i0(1'b0),
    .i1(uncache_data[63]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n59 [63]));
  binary_mux_s1_w1 \exu/lsu/mux27_b7  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [7]),
    .sel(unsign),
    .o(\exu/lsu/n59 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b8  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [8]),
    .sel(unsign),
    .o(\exu/lsu/n59 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux27_b9  (
    .i0(1'b0),
    .i1(\exu/lsu/n28 [9]),
    .sel(unsign),
    .o(\exu/lsu/n59 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  binary_mux_s1_w1 \exu/lsu/mux28_b0  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [0]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n60 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(67)
  binary_mux_s1_w1 \exu/lsu/mux28_b1  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [1]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n60 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(67)
  binary_mux_s1_w1 \exu/lsu/mux28_b10  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [7]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n60 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(67)
  binary_mux_s1_w1 \exu/lsu/mux28_b2  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [2]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n60 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(67)
  binary_mux_s1_w1 \exu/lsu/mux28_b3  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [3]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n60 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(67)
  binary_mux_s1_w1 \exu/lsu/mux28_b4  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [4]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n60 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(67)
  binary_mux_s1_w1 \exu/lsu/mux28_b5  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [5]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n60 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(67)
  binary_mux_s1_w1 \exu/lsu/mux28_b6  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [6]),
    .sel(\exu/lsu/n51 ),
    .o(\exu/lsu/n60 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(67)
  binary_mux_s1_w1 \exu/lsu/mux29_b0  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [0]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b1  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [1]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b10  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [10]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b11  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [11]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b12  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [12]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b13  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [13]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b14  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [14]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b15  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [15]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b2  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [2]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b3  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [3]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b4  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [4]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b5  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [5]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b6  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [6]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b7  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [7]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b8  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [8]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux29_b9  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [9]),
    .sel(\exu/lsu/n53 ),
    .o(\exu/lsu/n61 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  binary_mux_s1_w1 \exu/lsu/mux2_b16  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [0]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b17  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [1]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b18  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [2]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b19  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [3]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b20  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [4]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b21  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [5]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b22  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [6]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b23  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [7]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b24  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [8]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b25  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [9]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b26  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [10]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b27  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [11]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b28  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [12]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b29  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [13]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b30  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [14]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b31  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [15]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b32  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [16]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b33  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [17]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b34  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [18]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b35  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [19]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b36  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [20]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b37  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [21]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b38  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [22]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b39  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [23]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b40  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [24]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b41  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [25]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b42  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [26]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b43  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [27]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b44  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [28]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b45  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [29]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b46  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [30]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b47  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [31]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b48  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [32]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [48]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b49  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [33]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [49]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b50  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [34]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [50]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b51  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [35]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [51]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b52  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [36]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [52]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b53  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [37]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [53]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b54  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [38]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [54]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b55  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [39]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [55]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b56  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [40]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [56]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b57  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [41]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [57]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b58  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [42]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [58]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b59  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [43]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [59]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b60  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [44]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [60]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b61  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [45]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [61]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b62  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [46]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [62]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux2_b63  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [47]),
    .sel(\exu/lsu/n5 ),
    .o(\exu/lsu/n6 [63]));  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  binary_mux_s1_w1 \exu/lsu/mux30_b0  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [0]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b1  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [1]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b10  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [10]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b11  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [11]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b12  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [12]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b13  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [13]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b14  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [14]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b15  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [15]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b16  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [16]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b17  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [17]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b18  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [18]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b19  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [19]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b2  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [2]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b20  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [20]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b21  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [21]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b22  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [22]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b23  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [23]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b24  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [24]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b25  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [25]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b26  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [26]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b27  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [27]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b28  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [28]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b29  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [29]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b3  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [3]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b30  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [30]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b31  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [31]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b4  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [4]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b5  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [5]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b6  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [6]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b7  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [7]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b8  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [8]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux30_b9  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [9]),
    .sel(\exu/lsu/n56 ),
    .o(\exu/lsu/n63 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  binary_mux_s1_w1 \exu/lsu/mux31_b0  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [0]),
    .sel(unsign),
    .o(\exu/lsu/n65 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b1  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [1]),
    .sel(unsign),
    .o(\exu/lsu/n65 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b10  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [10]),
    .sel(unsign),
    .o(\exu/lsu/n65 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b11  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [11]),
    .sel(unsign),
    .o(\exu/lsu/n65 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b12  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [12]),
    .sel(unsign),
    .o(\exu/lsu/n65 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b13  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [13]),
    .sel(unsign),
    .o(\exu/lsu/n65 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b14  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [14]),
    .sel(unsign),
    .o(\exu/lsu/n65 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b15  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [15]),
    .sel(unsign),
    .o(\exu/lsu/n65 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b16  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [16]),
    .sel(unsign),
    .o(\exu/lsu/n65 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b17  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [17]),
    .sel(unsign),
    .o(\exu/lsu/n65 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b18  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [18]),
    .sel(unsign),
    .o(\exu/lsu/n65 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b19  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [19]),
    .sel(unsign),
    .o(\exu/lsu/n65 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b2  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [2]),
    .sel(unsign),
    .o(\exu/lsu/n65 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b20  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [20]),
    .sel(unsign),
    .o(\exu/lsu/n65 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b21  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [21]),
    .sel(unsign),
    .o(\exu/lsu/n65 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b22  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [22]),
    .sel(unsign),
    .o(\exu/lsu/n65 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b23  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [23]),
    .sel(unsign),
    .o(\exu/lsu/n65 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b24  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [24]),
    .sel(unsign),
    .o(\exu/lsu/n65 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b25  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [25]),
    .sel(unsign),
    .o(\exu/lsu/n65 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b26  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [26]),
    .sel(unsign),
    .o(\exu/lsu/n65 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b27  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [27]),
    .sel(unsign),
    .o(\exu/lsu/n65 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b28  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [28]),
    .sel(unsign),
    .o(\exu/lsu/n65 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b29  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [29]),
    .sel(unsign),
    .o(\exu/lsu/n65 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b3  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [3]),
    .sel(unsign),
    .o(\exu/lsu/n65 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b30  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [30]),
    .sel(unsign),
    .o(\exu/lsu/n65 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b31  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [31]),
    .sel(unsign),
    .o(\exu/lsu/n65 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b32  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [32]),
    .sel(unsign),
    .o(\exu/lsu/n65 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b33  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [33]),
    .sel(unsign),
    .o(\exu/lsu/n65 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b34  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [34]),
    .sel(unsign),
    .o(\exu/lsu/n65 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b35  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [35]),
    .sel(unsign),
    .o(\exu/lsu/n65 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b36  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [36]),
    .sel(unsign),
    .o(\exu/lsu/n65 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b37  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [37]),
    .sel(unsign),
    .o(\exu/lsu/n65 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b38  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [38]),
    .sel(unsign),
    .o(\exu/lsu/n65 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b39  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [39]),
    .sel(unsign),
    .o(\exu/lsu/n65 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b4  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [4]),
    .sel(unsign),
    .o(\exu/lsu/n65 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b40  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [40]),
    .sel(unsign),
    .o(\exu/lsu/n65 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b41  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [41]),
    .sel(unsign),
    .o(\exu/lsu/n65 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b42  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [42]),
    .sel(unsign),
    .o(\exu/lsu/n65 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b43  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [43]),
    .sel(unsign),
    .o(\exu/lsu/n65 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b44  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [44]),
    .sel(unsign),
    .o(\exu/lsu/n65 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b45  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [45]),
    .sel(unsign),
    .o(\exu/lsu/n65 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b46  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [46]),
    .sel(unsign),
    .o(\exu/lsu/n65 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b47  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [47]),
    .sel(unsign),
    .o(\exu/lsu/n65 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b48  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [48]),
    .sel(unsign),
    .o(\exu/lsu/n65 [48]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b49  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [49]),
    .sel(unsign),
    .o(\exu/lsu/n65 [49]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b5  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [5]),
    .sel(unsign),
    .o(\exu/lsu/n65 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b50  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [50]),
    .sel(unsign),
    .o(\exu/lsu/n65 [50]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b51  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [51]),
    .sel(unsign),
    .o(\exu/lsu/n65 [51]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b52  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [52]),
    .sel(unsign),
    .o(\exu/lsu/n65 [52]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b53  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [53]),
    .sel(unsign),
    .o(\exu/lsu/n65 [53]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b54  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [54]),
    .sel(unsign),
    .o(\exu/lsu/n65 [54]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b55  (
    .i0(1'b0),
    .i1(\exu/lsu/data_lsu_cache_shift [55]),
    .sel(unsign),
    .o(\exu/lsu/n65 [55]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  AL_MUX \exu/lsu/mux31_b56  (
    .i0(1'b0),
    .i1(data_read[56]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n65 [56]));
  AL_MUX \exu/lsu/mux31_b57  (
    .i0(1'b0),
    .i1(data_read[57]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n65 [57]));
  AL_MUX \exu/lsu/mux31_b58  (
    .i0(1'b0),
    .i1(data_read[58]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n65 [58]));
  AL_MUX \exu/lsu/mux31_b59  (
    .i0(1'b0),
    .i1(data_read[59]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n65 [59]));
  binary_mux_s1_w1 \exu/lsu/mux31_b6  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [6]),
    .sel(unsign),
    .o(\exu/lsu/n65 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  AL_MUX \exu/lsu/mux31_b60  (
    .i0(1'b0),
    .i1(data_read[60]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n65 [60]));
  AL_MUX \exu/lsu/mux31_b61  (
    .i0(1'b0),
    .i1(data_read[61]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n65 [61]));
  AL_MUX \exu/lsu/mux31_b62  (
    .i0(1'b0),
    .i1(data_read[62]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n65 [62]));
  AL_MUX \exu/lsu/mux31_b63  (
    .i0(1'b0),
    .i1(data_read[63]),
    .sel(\exu/lsu/mux27_b56_sel_is_3_o ),
    .o(\exu/lsu/n65 [63]));
  binary_mux_s1_w1 \exu/lsu/mux31_b7  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [7]),
    .sel(unsign),
    .o(\exu/lsu/n65 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b8  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [8]),
    .sel(unsign),
    .o(\exu/lsu/n65 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux31_b9  (
    .i0(1'b0),
    .i1(\exu/lsu/n42 [9]),
    .sel(unsign),
    .o(\exu/lsu/n65 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  binary_mux_s1_w1 \exu/lsu/mux3_b24  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [0]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b25  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [1]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b26  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [2]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b27  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [3]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b28  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [4]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b29  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [5]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b30  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [6]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b31  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [7]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b32  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [8]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b33  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [9]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b34  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [10]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b35  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [11]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b36  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [12]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b37  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [13]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b38  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [14]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b39  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [15]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b40  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [16]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b41  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [17]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b42  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [18]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b43  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [19]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b44  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [20]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b45  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [21]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b46  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [22]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b47  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [23]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b48  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [24]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [48]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b49  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [25]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [49]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b50  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [26]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [50]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b51  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [27]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [51]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b52  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [28]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [52]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b53  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [29]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [53]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b54  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [30]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [54]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b55  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [31]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [55]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b56  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [32]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [56]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b57  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [33]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [57]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b58  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [34]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [58]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b59  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [35]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [59]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b60  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [36]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [60]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b61  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [37]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [61]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b62  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [38]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [62]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux3_b63  (
    .i0(1'b0),
    .i1(\exu/alu_data_mem_csr [39]),
    .sel(\exu/lsu/n8 ),
    .o(\exu/lsu/n9 [63]));  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  binary_mux_s1_w1 \exu/lsu/mux8_b0  (
    .i0(1'b0),
    .i1(uncache_data[0]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b1  (
    .i0(1'b0),
    .i1(uncache_data[1]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b10  (
    .i0(1'b0),
    .i1(uncache_data[10]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b11  (
    .i0(1'b0),
    .i1(uncache_data[11]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b12  (
    .i0(1'b0),
    .i1(uncache_data[12]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b13  (
    .i0(1'b0),
    .i1(uncache_data[13]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b14  (
    .i0(1'b0),
    .i1(uncache_data[14]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b15  (
    .i0(1'b0),
    .i1(uncache_data[15]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b16  (
    .i0(1'b0),
    .i1(uncache_data[16]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b17  (
    .i0(1'b0),
    .i1(uncache_data[17]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b18  (
    .i0(1'b0),
    .i1(uncache_data[18]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b19  (
    .i0(1'b0),
    .i1(uncache_data[19]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b2  (
    .i0(1'b0),
    .i1(uncache_data[2]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b20  (
    .i0(1'b0),
    .i1(uncache_data[20]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b21  (
    .i0(1'b0),
    .i1(uncache_data[21]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b22  (
    .i0(1'b0),
    .i1(uncache_data[22]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b23  (
    .i0(1'b0),
    .i1(uncache_data[23]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b24  (
    .i0(1'b0),
    .i1(uncache_data[24]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b25  (
    .i0(1'b0),
    .i1(uncache_data[25]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b26  (
    .i0(1'b0),
    .i1(uncache_data[26]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b27  (
    .i0(1'b0),
    .i1(uncache_data[27]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b28  (
    .i0(1'b0),
    .i1(uncache_data[28]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b29  (
    .i0(1'b0),
    .i1(uncache_data[29]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b3  (
    .i0(1'b0),
    .i1(uncache_data[3]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b30  (
    .i0(1'b0),
    .i1(uncache_data[30]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b31  (
    .i0(1'b0),
    .i1(uncache_data[31]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b32  (
    .i0(1'b0),
    .i1(uncache_data[32]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b33  (
    .i0(1'b0),
    .i1(uncache_data[33]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b34  (
    .i0(1'b0),
    .i1(uncache_data[34]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b35  (
    .i0(1'b0),
    .i1(uncache_data[35]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b36  (
    .i0(1'b0),
    .i1(uncache_data[36]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b37  (
    .i0(1'b0),
    .i1(uncache_data[37]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b38  (
    .i0(1'b0),
    .i1(uncache_data[38]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b39  (
    .i0(1'b0),
    .i1(uncache_data[39]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b4  (
    .i0(1'b0),
    .i1(uncache_data[4]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b40  (
    .i0(1'b0),
    .i1(uncache_data[40]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b41  (
    .i0(1'b0),
    .i1(uncache_data[41]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b42  (
    .i0(1'b0),
    .i1(uncache_data[42]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b43  (
    .i0(1'b0),
    .i1(uncache_data[43]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b44  (
    .i0(1'b0),
    .i1(uncache_data[44]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b45  (
    .i0(1'b0),
    .i1(uncache_data[45]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b46  (
    .i0(1'b0),
    .i1(uncache_data[46]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b47  (
    .i0(1'b0),
    .i1(uncache_data[47]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b48  (
    .i0(1'b0),
    .i1(uncache_data[48]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [48]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b49  (
    .i0(1'b0),
    .i1(uncache_data[49]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [49]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b5  (
    .i0(1'b0),
    .i1(uncache_data[5]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b50  (
    .i0(1'b0),
    .i1(uncache_data[50]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [50]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b51  (
    .i0(1'b0),
    .i1(uncache_data[51]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [51]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b52  (
    .i0(1'b0),
    .i1(uncache_data[52]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [52]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b53  (
    .i0(1'b0),
    .i1(uncache_data[53]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [53]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b54  (
    .i0(1'b0),
    .i1(uncache_data[54]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [54]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b55  (
    .i0(1'b0),
    .i1(uncache_data[55]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [55]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b6  (
    .i0(1'b0),
    .i1(uncache_data[6]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b7  (
    .i0(1'b0),
    .i1(uncache_data[7]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b8  (
    .i0(1'b0),
    .i1(uncache_data[8]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux8_b9  (
    .i0(1'b0),
    .i1(uncache_data[9]),
    .sel(\exu/lsu/n0 ),
    .o(\exu/lsu/n22 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(42)
  binary_mux_s1_w1 \exu/lsu/mux9_b0  (
    .i0(1'b0),
    .i1(uncache_data[8]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [0]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b1  (
    .i0(1'b0),
    .i1(uncache_data[9]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [1]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b10  (
    .i0(1'b0),
    .i1(uncache_data[18]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [10]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b11  (
    .i0(1'b0),
    .i1(uncache_data[19]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [11]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b12  (
    .i0(1'b0),
    .i1(uncache_data[20]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [12]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b13  (
    .i0(1'b0),
    .i1(uncache_data[21]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [13]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b14  (
    .i0(1'b0),
    .i1(uncache_data[22]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [14]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b15  (
    .i0(1'b0),
    .i1(uncache_data[23]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [15]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b16  (
    .i0(1'b0),
    .i1(uncache_data[24]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [16]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b17  (
    .i0(1'b0),
    .i1(uncache_data[25]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [17]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b18  (
    .i0(1'b0),
    .i1(uncache_data[26]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [18]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b19  (
    .i0(1'b0),
    .i1(uncache_data[27]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [19]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b2  (
    .i0(1'b0),
    .i1(uncache_data[10]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [2]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b20  (
    .i0(1'b0),
    .i1(uncache_data[28]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [20]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b21  (
    .i0(1'b0),
    .i1(uncache_data[29]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [21]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b22  (
    .i0(1'b0),
    .i1(uncache_data[30]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [22]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b23  (
    .i0(1'b0),
    .i1(uncache_data[31]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [23]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b24  (
    .i0(1'b0),
    .i1(uncache_data[32]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [24]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b25  (
    .i0(1'b0),
    .i1(uncache_data[33]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [25]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b26  (
    .i0(1'b0),
    .i1(uncache_data[34]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [26]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b27  (
    .i0(1'b0),
    .i1(uncache_data[35]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [27]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b28  (
    .i0(1'b0),
    .i1(uncache_data[36]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [28]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b29  (
    .i0(1'b0),
    .i1(uncache_data[37]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [29]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b3  (
    .i0(1'b0),
    .i1(uncache_data[11]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [3]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b30  (
    .i0(1'b0),
    .i1(uncache_data[38]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [30]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b31  (
    .i0(1'b0),
    .i1(uncache_data[39]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [31]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b32  (
    .i0(1'b0),
    .i1(uncache_data[40]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [32]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b33  (
    .i0(1'b0),
    .i1(uncache_data[41]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [33]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b34  (
    .i0(1'b0),
    .i1(uncache_data[42]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [34]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b35  (
    .i0(1'b0),
    .i1(uncache_data[43]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [35]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b36  (
    .i0(1'b0),
    .i1(uncache_data[44]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [36]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b37  (
    .i0(1'b0),
    .i1(uncache_data[45]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [37]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b38  (
    .i0(1'b0),
    .i1(uncache_data[46]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [38]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b39  (
    .i0(1'b0),
    .i1(uncache_data[47]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [39]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b4  (
    .i0(1'b0),
    .i1(uncache_data[12]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [4]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b40  (
    .i0(1'b0),
    .i1(uncache_data[48]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [40]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b41  (
    .i0(1'b0),
    .i1(uncache_data[49]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [41]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b42  (
    .i0(1'b0),
    .i1(uncache_data[50]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [42]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b43  (
    .i0(1'b0),
    .i1(uncache_data[51]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [43]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b44  (
    .i0(1'b0),
    .i1(uncache_data[52]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [44]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b45  (
    .i0(1'b0),
    .i1(uncache_data[53]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [45]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b46  (
    .i0(1'b0),
    .i1(uncache_data[54]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [46]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b47  (
    .i0(1'b0),
    .i1(uncache_data[55]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [47]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b48  (
    .i0(1'b0),
    .i1(uncache_data[56]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [48]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b49  (
    .i0(1'b0),
    .i1(uncache_data[57]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [49]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b5  (
    .i0(1'b0),
    .i1(uncache_data[13]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [5]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b50  (
    .i0(1'b0),
    .i1(uncache_data[58]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [50]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b51  (
    .i0(1'b0),
    .i1(uncache_data[59]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [51]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b52  (
    .i0(1'b0),
    .i1(uncache_data[60]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [52]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b53  (
    .i0(1'b0),
    .i1(uncache_data[61]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [53]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b54  (
    .i0(1'b0),
    .i1(uncache_data[62]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [54]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b55  (
    .i0(1'b0),
    .i1(uncache_data[63]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [55]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b6  (
    .i0(1'b0),
    .i1(uncache_data[14]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [6]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b7  (
    .i0(1'b0),
    .i1(uncache_data[15]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [7]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b8  (
    .i0(1'b0),
    .i1(uncache_data[16]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [8]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  binary_mux_s1_w1 \exu/lsu/mux9_b9  (
    .i0(1'b0),
    .i1(uncache_data[17]),
    .sel(\exu/lsu/n2 ),
    .o(\exu/lsu/n23 [9]));  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u10  (\exu/data_lsu_cache [23], \exu/lsu/n64 [23], \exu/lsu/n65 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u100  (\exu/lsu/n64 [5], \exu/lsu/n62 [5], \exu/lsu/n63 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u101  (\exu/lsu/n64 [6], \exu/lsu/n62 [6], \exu/lsu/n63 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u102  (\exu/lsu/n64 [7], \exu/lsu/n62 [7], \exu/lsu/n63 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u103  (\exu/lsu/n64 [8], \exu/lsu/n62 [8], \exu/lsu/n63 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u104  (\exu/lsu/n64 [9], \exu/lsu/n62 [9], \exu/lsu/n63 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u105  (\exu/lsu/n64 [10], \exu/lsu/n62 [10], \exu/lsu/n63 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u106  (\exu/lsu/n64 [11], \exu/lsu/n62 [11], \exu/lsu/n63 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u107  (\exu/lsu/n64 [12], \exu/lsu/n62 [12], \exu/lsu/n63 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u108  (\exu/lsu/n64 [13], \exu/lsu/n62 [13], \exu/lsu/n63 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u109  (\exu/lsu/n64 [14], \exu/lsu/n62 [14], \exu/lsu/n63 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u11  (\exu/data_lsu_cache [22], \exu/lsu/n64 [22], \exu/lsu/n65 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u110  (\exu/lsu/n64 [15], \exu/lsu/n62 [15], \exu/lsu/n63 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u111  (\exu/lsu/n64 [16], \exu/lsu/n62 [15], \exu/lsu/n63 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u112  (\exu/lsu/n64 [17], \exu/lsu/n62 [15], \exu/lsu/n63 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1120  (\exu/lsu/n10 [24], \exu/lsu/n7 [24], \exu/lsu/n9 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1121  (\exu/lsu/n10 [25], \exu/lsu/n7 [25], \exu/lsu/n9 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1122  (\exu/lsu/n10 [26], \exu/lsu/n7 [26], \exu/lsu/n9 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1123  (\exu/lsu/n10 [27], \exu/lsu/n7 [27], \exu/lsu/n9 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1124  (\exu/lsu/n10 [28], \exu/lsu/n7 [28], \exu/lsu/n9 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1125  (\exu/lsu/n10 [29], \exu/lsu/n7 [29], \exu/lsu/n9 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1126  (\exu/lsu/n10 [30], \exu/lsu/n7 [30], \exu/lsu/n9 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1127  (\exu/lsu/n10 [31], \exu/lsu/n7 [31], \exu/lsu/n9 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1128  (\exu/lsu/n10 [32], \exu/lsu/n7 [32], \exu/lsu/n9 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1129  (\exu/lsu/n10 [33], \exu/lsu/n7 [33], \exu/lsu/n9 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u113  (\exu/lsu/n64 [18], \exu/lsu/n62 [15], \exu/lsu/n63 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1130  (\exu/lsu/n10 [34], \exu/lsu/n7 [34], \exu/lsu/n9 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1131  (\exu/lsu/n10 [35], \exu/lsu/n7 [35], \exu/lsu/n9 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1132  (\exu/lsu/n10 [36], \exu/lsu/n7 [36], \exu/lsu/n9 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1133  (\exu/lsu/n10 [37], \exu/lsu/n7 [37], \exu/lsu/n9 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1134  (\exu/lsu/n10 [38], \exu/lsu/n7 [38], \exu/lsu/n9 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1135  (\exu/lsu/n10 [39], \exu/lsu/n7 [39], \exu/lsu/n9 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1136  (\exu/lsu/n10 [40], \exu/lsu/n7 [40], \exu/lsu/n9 [40]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1137  (\exu/lsu/n10 [41], \exu/lsu/n7 [41], \exu/lsu/n9 [41]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1138  (\exu/lsu/n10 [42], \exu/lsu/n7 [42], \exu/lsu/n9 [42]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1139  (\exu/lsu/n10 [43], \exu/lsu/n7 [43], \exu/lsu/n9 [43]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u114  (\exu/lsu/n64 [19], \exu/lsu/n62 [15], \exu/lsu/n63 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1140  (\exu/lsu/n10 [44], \exu/lsu/n7 [44], \exu/lsu/n9 [44]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1141  (\exu/lsu/n10 [45], \exu/lsu/n7 [45], \exu/lsu/n9 [45]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1142  (\exu/lsu/n10 [46], \exu/lsu/n7 [46], \exu/lsu/n9 [46]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1143  (\exu/lsu/n10 [47], \exu/lsu/n7 [47], \exu/lsu/n9 [47]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1144  (\exu/lsu/n10 [48], \exu/lsu/n7 [48], \exu/lsu/n9 [48]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1145  (\exu/lsu/n10 [49], \exu/lsu/n7 [49], \exu/lsu/n9 [49]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1146  (\exu/lsu/n10 [50], \exu/lsu/n7 [50], \exu/lsu/n9 [50]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1147  (\exu/lsu/n10 [51], \exu/lsu/n7 [51], \exu/lsu/n9 [51]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1148  (\exu/lsu/n10 [52], \exu/lsu/n7 [52], \exu/lsu/n9 [52]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1149  (\exu/lsu/n10 [53], \exu/lsu/n7 [53], \exu/lsu/n9 [53]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u115  (\exu/lsu/n64 [20], \exu/lsu/n62 [15], \exu/lsu/n63 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1150  (\exu/lsu/n10 [54], \exu/lsu/n7 [54], \exu/lsu/n9 [54]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1151  (\exu/lsu/n10 [55], \exu/lsu/n7 [55], \exu/lsu/n9 [55]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1152  (\exu/lsu/n10 [56], \exu/lsu/n7 [56], \exu/lsu/n9 [56]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1153  (\exu/lsu/n10 [57], \exu/lsu/n7 [57], \exu/lsu/n9 [57]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1154  (\exu/lsu/n10 [58], \exu/lsu/n7 [58], \exu/lsu/n9 [58]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1155  (\exu/lsu/n10 [59], \exu/lsu/n7 [59], \exu/lsu/n9 [59]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1156  (\exu/lsu/n10 [60], \exu/lsu/n7 [60], \exu/lsu/n9 [60]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1157  (\exu/lsu/n10 [61], \exu/lsu/n7 [61], \exu/lsu/n9 [61]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1158  (\exu/lsu/n10 [62], \exu/lsu/n7 [62], \exu/lsu/n9 [62]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u1159  (\exu/lsu/n10 [63], \exu/lsu/n7 [63], \exu/lsu/n9 [63]);  // ../../RTL/CPU/EX/LSU/lsu.v(35)
  or \exu/lsu/u116  (\exu/lsu/n64 [21], \exu/lsu/n62 [15], \exu/lsu/n63 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u117  (\exu/lsu/n64 [22], \exu/lsu/n62 [15], \exu/lsu/n63 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1175  (\exu/lsu/n7 [16], \exu/lsu/n4 [16], \exu/lsu/n6 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1176  (\exu/lsu/n7 [17], \exu/lsu/n4 [17], \exu/lsu/n6 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1177  (\exu/lsu/n7 [18], \exu/lsu/n4 [18], \exu/lsu/n6 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1178  (\exu/lsu/n7 [19], \exu/lsu/n4 [19], \exu/lsu/n6 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1179  (\exu/lsu/n7 [20], \exu/lsu/n4 [20], \exu/lsu/n6 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u118  (\exu/lsu/n64 [23], \exu/lsu/n62 [15], \exu/lsu/n63 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1180  (\exu/lsu/n7 [21], \exu/lsu/n4 [21], \exu/lsu/n6 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1181  (\exu/lsu/n7 [22], \exu/lsu/n4 [22], \exu/lsu/n6 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1182  (\exu/lsu/n7 [23], \exu/lsu/n4 [23], \exu/lsu/n6 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1183  (\exu/lsu/n7 [24], \exu/lsu/n4 [24], \exu/lsu/n6 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1184  (\exu/lsu/n7 [25], \exu/lsu/n4 [25], \exu/lsu/n6 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1185  (\exu/lsu/n7 [26], \exu/lsu/n4 [26], \exu/lsu/n6 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1186  (\exu/lsu/n7 [27], \exu/lsu/n4 [27], \exu/lsu/n6 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1187  (\exu/lsu/n7 [28], \exu/lsu/n4 [28], \exu/lsu/n6 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1188  (\exu/lsu/n7 [29], \exu/lsu/n4 [29], \exu/lsu/n6 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1189  (\exu/lsu/n7 [30], \exu/lsu/n4 [30], \exu/lsu/n6 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u119  (\exu/lsu/n64 [24], \exu/lsu/n62 [15], \exu/lsu/n63 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1190  (\exu/lsu/n7 [31], \exu/lsu/n4 [31], \exu/lsu/n6 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1191  (\exu/lsu/n7 [32], \exu/lsu/n4 [32], \exu/lsu/n6 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1192  (\exu/lsu/n7 [33], \exu/lsu/n4 [33], \exu/lsu/n6 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1193  (\exu/lsu/n7 [34], \exu/lsu/n4 [34], \exu/lsu/n6 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1194  (\exu/lsu/n7 [35], \exu/lsu/n4 [35], \exu/lsu/n6 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1195  (\exu/lsu/n7 [36], \exu/lsu/n4 [36], \exu/lsu/n6 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1196  (\exu/lsu/n7 [37], \exu/lsu/n4 [37], \exu/lsu/n6 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1197  (\exu/lsu/n7 [38], \exu/lsu/n4 [38], \exu/lsu/n6 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1198  (\exu/lsu/n7 [39], \exu/lsu/n4 [39], \exu/lsu/n6 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1199  (\exu/lsu/n7 [40], \exu/lsu/n4 [40], \exu/lsu/n6 [40]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u120  (\exu/lsu/n64 [25], \exu/lsu/n62 [15], \exu/lsu/n63 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1200  (\exu/lsu/n7 [41], \exu/lsu/n4 [41], \exu/lsu/n6 [41]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1201  (\exu/lsu/n7 [42], \exu/lsu/n4 [42], \exu/lsu/n6 [42]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1202  (\exu/lsu/n7 [43], \exu/lsu/n4 [43], \exu/lsu/n6 [43]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1203  (\exu/lsu/n7 [44], \exu/lsu/n4 [44], \exu/lsu/n6 [44]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1204  (\exu/lsu/n7 [45], \exu/lsu/n4 [45], \exu/lsu/n6 [45]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1205  (\exu/lsu/n7 [46], \exu/lsu/n4 [46], \exu/lsu/n6 [46]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1206  (\exu/lsu/n7 [47], \exu/lsu/n4 [47], \exu/lsu/n6 [47]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1207  (\exu/lsu/n7 [48], \exu/lsu/n4 [48], \exu/lsu/n6 [48]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1208  (\exu/lsu/n7 [49], \exu/lsu/n4 [49], \exu/lsu/n6 [49]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1209  (\exu/lsu/n7 [50], \exu/lsu/n4 [50], \exu/lsu/n6 [50]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u121  (\exu/lsu/n64 [26], \exu/lsu/n62 [15], \exu/lsu/n63 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1210  (\exu/lsu/n7 [51], \exu/lsu/n4 [51], \exu/lsu/n6 [51]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1211  (\exu/lsu/n7 [52], \exu/lsu/n4 [52], \exu/lsu/n6 [52]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1212  (\exu/lsu/n7 [53], \exu/lsu/n4 [53], \exu/lsu/n6 [53]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1213  (\exu/lsu/n7 [54], \exu/lsu/n4 [54], \exu/lsu/n6 [54]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1214  (\exu/lsu/n7 [55], \exu/lsu/n4 [55], \exu/lsu/n6 [55]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1215  (\exu/lsu/n7 [56], \exu/lsu/n4 [56], \exu/lsu/n6 [56]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1216  (\exu/lsu/n7 [57], \exu/lsu/n4 [57], \exu/lsu/n6 [57]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1217  (\exu/lsu/n7 [58], \exu/lsu/n4 [58], \exu/lsu/n6 [58]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1218  (\exu/lsu/n7 [59], \exu/lsu/n4 [59], \exu/lsu/n6 [59]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1219  (\exu/lsu/n7 [60], \exu/lsu/n4 [60], \exu/lsu/n6 [60]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u122  (\exu/lsu/n64 [27], \exu/lsu/n62 [15], \exu/lsu/n63 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1220  (\exu/lsu/n7 [61], \exu/lsu/n4 [61], \exu/lsu/n6 [61]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1221  (\exu/lsu/n7 [62], \exu/lsu/n4 [62], \exu/lsu/n6 [62]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u1222  (\exu/lsu/n7 [63], \exu/lsu/n4 [63], \exu/lsu/n6 [63]);  // ../../RTL/CPU/EX/LSU/lsu.v(34)
  or \exu/lsu/u123  (\exu/lsu/n64 [28], \exu/lsu/n62 [15], \exu/lsu/n63 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1230  (\exu/lsu/n4 [8], \exu/lsu/n1 [8], \exu/lsu/n3 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1231  (\exu/lsu/n4 [9], \exu/lsu/n1 [9], \exu/lsu/n3 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1232  (\exu/lsu/n4 [10], \exu/lsu/n1 [10], \exu/lsu/n3 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1233  (\exu/lsu/n4 [11], \exu/lsu/n1 [11], \exu/lsu/n3 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1234  (\exu/lsu/n4 [12], \exu/lsu/n1 [12], \exu/lsu/n3 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1235  (\exu/lsu/n4 [13], \exu/lsu/n1 [13], \exu/lsu/n3 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1236  (\exu/lsu/n4 [14], \exu/lsu/n1 [14], \exu/lsu/n3 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1237  (\exu/lsu/n4 [15], \exu/lsu/n1 [15], \exu/lsu/n3 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1238  (\exu/lsu/n4 [16], \exu/lsu/n1 [16], \exu/lsu/n3 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1239  (\exu/lsu/n4 [17], \exu/lsu/n1 [17], \exu/lsu/n3 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u124  (\exu/lsu/n64 [29], \exu/lsu/n62 [15], \exu/lsu/n63 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1240  (\exu/lsu/n4 [18], \exu/lsu/n1 [18], \exu/lsu/n3 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1241  (\exu/lsu/n4 [19], \exu/lsu/n1 [19], \exu/lsu/n3 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1242  (\exu/lsu/n4 [20], \exu/lsu/n1 [20], \exu/lsu/n3 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1243  (\exu/lsu/n4 [21], \exu/lsu/n1 [21], \exu/lsu/n3 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1244  (\exu/lsu/n4 [22], \exu/lsu/n1 [22], \exu/lsu/n3 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1245  (\exu/lsu/n4 [23], \exu/lsu/n1 [23], \exu/lsu/n3 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1246  (\exu/lsu/n4 [24], \exu/lsu/n1 [24], \exu/lsu/n3 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1247  (\exu/lsu/n4 [25], \exu/lsu/n1 [25], \exu/lsu/n3 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1248  (\exu/lsu/n4 [26], \exu/lsu/n1 [26], \exu/lsu/n3 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1249  (\exu/lsu/n4 [27], \exu/lsu/n1 [27], \exu/lsu/n3 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u125  (\exu/lsu/n64 [30], \exu/lsu/n62 [15], \exu/lsu/n63 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1250  (\exu/lsu/n4 [28], \exu/lsu/n1 [28], \exu/lsu/n3 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1251  (\exu/lsu/n4 [29], \exu/lsu/n1 [29], \exu/lsu/n3 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1252  (\exu/lsu/n4 [30], \exu/lsu/n1 [30], \exu/lsu/n3 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1253  (\exu/lsu/n4 [31], \exu/lsu/n1 [31], \exu/lsu/n3 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1254  (\exu/lsu/n4 [32], \exu/lsu/n1 [32], \exu/lsu/n3 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1255  (\exu/lsu/n4 [33], \exu/lsu/n1 [33], \exu/lsu/n3 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1256  (\exu/lsu/n4 [34], \exu/lsu/n1 [34], \exu/lsu/n3 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1257  (\exu/lsu/n4 [35], \exu/lsu/n1 [35], \exu/lsu/n3 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1258  (\exu/lsu/n4 [36], \exu/lsu/n1 [36], \exu/lsu/n3 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1259  (\exu/lsu/n4 [37], \exu/lsu/n1 [37], \exu/lsu/n3 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u126  (\exu/lsu/n64 [31], \exu/lsu/n62 [15], \exu/lsu/n63 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u1260  (\exu/lsu/n4 [38], \exu/lsu/n1 [38], \exu/lsu/n3 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1261  (\exu/lsu/n4 [39], \exu/lsu/n1 [39], \exu/lsu/n3 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1262  (\exu/lsu/n4 [40], \exu/lsu/n1 [40], \exu/lsu/n3 [40]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1263  (\exu/lsu/n4 [41], \exu/lsu/n1 [41], \exu/lsu/n3 [41]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1264  (\exu/lsu/n4 [42], \exu/lsu/n1 [42], \exu/lsu/n3 [42]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1265  (\exu/lsu/n4 [43], \exu/lsu/n1 [43], \exu/lsu/n3 [43]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1266  (\exu/lsu/n4 [44], \exu/lsu/n1 [44], \exu/lsu/n3 [44]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1267  (\exu/lsu/n4 [45], \exu/lsu/n1 [45], \exu/lsu/n3 [45]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1268  (\exu/lsu/n4 [46], \exu/lsu/n1 [46], \exu/lsu/n3 [46]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1269  (\exu/lsu/n4 [47], \exu/lsu/n1 [47], \exu/lsu/n3 [47]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1270  (\exu/lsu/n4 [48], \exu/lsu/n1 [48], \exu/lsu/n3 [48]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1271  (\exu/lsu/n4 [49], \exu/lsu/n1 [49], \exu/lsu/n3 [49]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1272  (\exu/lsu/n4 [50], \exu/lsu/n1 [50], \exu/lsu/n3 [50]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1273  (\exu/lsu/n4 [51], \exu/lsu/n1 [51], \exu/lsu/n3 [51]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1274  (\exu/lsu/n4 [52], \exu/lsu/n1 [52], \exu/lsu/n3 [52]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1275  (\exu/lsu/n4 [53], \exu/lsu/n1 [53], \exu/lsu/n3 [53]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1276  (\exu/lsu/n4 [54], \exu/lsu/n1 [54], \exu/lsu/n3 [54]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1277  (\exu/lsu/n4 [55], \exu/lsu/n1 [55], \exu/lsu/n3 [55]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1278  (\exu/lsu/n4 [56], \exu/lsu/n1 [56], \exu/lsu/n3 [56]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1279  (\exu/lsu/n4 [57], \exu/lsu/n1 [57], \exu/lsu/n3 [57]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1280  (\exu/lsu/n4 [58], \exu/lsu/n1 [58], \exu/lsu/n3 [58]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1281  (\exu/lsu/n4 [59], \exu/lsu/n1 [59], \exu/lsu/n3 [59]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1282  (\exu/lsu/n4 [60], \exu/lsu/n1 [60], \exu/lsu/n3 [60]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1283  (\exu/lsu/n4 [61], \exu/lsu/n1 [61], \exu/lsu/n3 [61]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1284  (\exu/lsu/n4 [62], \exu/lsu/n1 [62], \exu/lsu/n3 [62]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u1285  (\exu/lsu/n4 [63], \exu/lsu/n1 [63], \exu/lsu/n3 [63]);  // ../../RTL/CPU/EX/LSU/lsu.v(33)
  or \exu/lsu/u13  (\exu/data_lsu_cache [21], \exu/lsu/n64 [21], \exu/lsu/n65 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u14  (\exu/lsu/n24 [0], \exu/lsu/n22 [0], \exu/lsu/n23 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u15  (\exu/data_lsu_cache [20], \exu/lsu/n64 [20], \exu/lsu/n65 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u159  (\exu/lsu/n62 [1], \exu/lsu/n60 [1], \exu/lsu/n61 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u16  (\exu/lsu/n26 [0], \exu/lsu/n24 [0], \exu/lsu/n25 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u160  (\exu/lsu/n62 [2], \exu/lsu/n60 [2], \exu/lsu/n61 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u161  (\exu/lsu/n62 [3], \exu/lsu/n60 [3], \exu/lsu/n61 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u162  (\exu/lsu/n62 [4], \exu/lsu/n60 [4], \exu/lsu/n61 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u163  (\exu/lsu/n62 [5], \exu/lsu/n60 [5], \exu/lsu/n61 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u164  (\exu/lsu/n62 [6], \exu/lsu/n60 [6], \exu/lsu/n61 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u165  (\exu/lsu/n62 [7], \exu/lsu/n60 [10], \exu/lsu/n61 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u166  (\exu/lsu/n62 [8], \exu/lsu/n60 [10], \exu/lsu/n61 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u167  (\exu/lsu/n62 [9], \exu/lsu/n60 [10], \exu/lsu/n61 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u168  (\exu/lsu/n62 [10], \exu/lsu/n60 [10], \exu/lsu/n61 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u169  (\exu/lsu/n62 [11], \exu/lsu/n60 [10], \exu/lsu/n61 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u17  (\exu/data_lsu_cache [19], \exu/lsu/n64 [19], \exu/lsu/n65 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u170  (\exu/lsu/n62 [12], \exu/lsu/n60 [10], \exu/lsu/n61 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u171  (\exu/lsu/n62 [13], \exu/lsu/n60 [10], \exu/lsu/n61 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u172  (\exu/lsu/n62 [14], \exu/lsu/n60 [10], \exu/lsu/n61 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u173  (\exu/lsu/n62 [15], \exu/lsu/n60 [10], \exu/lsu/n61 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u18  (\exu/lsu/n28 [0], \exu/lsu/n26 [0], \exu/lsu/n27 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u19  (\exu/data_lsu_cache [18], \exu/lsu/n64 [18], \exu/lsu/n65 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u2  (\exu/data_lsu_cache [25], \exu/lsu/n64 [25], \exu/lsu/n65 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u21  (\exu/data_lsu_cache [17], \exu/lsu/n64 [17], \exu/lsu/n65 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u222  (\exu/data_lsu_uncache [1], \exu/lsu/n58 [1], \exu/lsu/n59 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u223  (\exu/data_lsu_uncache [2], \exu/lsu/n58 [2], \exu/lsu/n59 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u224  (\exu/data_lsu_uncache [3], \exu/lsu/n58 [3], \exu/lsu/n59 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u225  (\exu/data_lsu_uncache [4], \exu/lsu/n58 [4], \exu/lsu/n59 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u226  (\exu/data_lsu_uncache [5], \exu/lsu/n58 [5], \exu/lsu/n59 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u227  (\exu/data_lsu_uncache [6], \exu/lsu/n58 [6], \exu/lsu/n59 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u228  (\exu/data_lsu_uncache [7], \exu/lsu/n58 [7], \exu/lsu/n59 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u229  (\exu/data_lsu_uncache [8], \exu/lsu/n58 [8], \exu/lsu/n59 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u23  (\exu/data_lsu_cache [16], \exu/lsu/n64 [16], \exu/lsu/n65 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u230  (\exu/data_lsu_uncache [9], \exu/lsu/n58 [9], \exu/lsu/n59 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u231  (\exu/data_lsu_uncache [10], \exu/lsu/n58 [10], \exu/lsu/n59 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u232  (\exu/data_lsu_uncache [11], \exu/lsu/n58 [11], \exu/lsu/n59 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u233  (\exu/data_lsu_uncache [12], \exu/lsu/n58 [12], \exu/lsu/n59 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u234  (\exu/data_lsu_uncache [13], \exu/lsu/n58 [13], \exu/lsu/n59 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u235  (\exu/data_lsu_uncache [14], \exu/lsu/n58 [14], \exu/lsu/n59 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u236  (\exu/data_lsu_uncache [15], \exu/lsu/n58 [15], \exu/lsu/n59 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u237  (\exu/data_lsu_uncache [16], \exu/lsu/n58 [16], \exu/lsu/n59 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u238  (\exu/data_lsu_uncache [17], \exu/lsu/n58 [17], \exu/lsu/n59 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u239  (\exu/data_lsu_uncache [18], \exu/lsu/n58 [18], \exu/lsu/n59 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u240  (\exu/data_lsu_uncache [19], \exu/lsu/n58 [19], \exu/lsu/n59 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u241  (\exu/data_lsu_uncache [20], \exu/lsu/n58 [20], \exu/lsu/n59 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u242  (\exu/data_lsu_uncache [21], \exu/lsu/n58 [21], \exu/lsu/n59 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u243  (\exu/data_lsu_uncache [22], \exu/lsu/n58 [22], \exu/lsu/n59 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u244  (\exu/data_lsu_uncache [23], \exu/lsu/n58 [23], \exu/lsu/n59 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u245  (\exu/data_lsu_uncache [24], \exu/lsu/n58 [24], \exu/lsu/n59 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u246  (\exu/data_lsu_uncache [25], \exu/lsu/n58 [25], \exu/lsu/n59 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u247  (\exu/data_lsu_uncache [26], \exu/lsu/n58 [26], \exu/lsu/n59 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u248  (\exu/data_lsu_uncache [27], \exu/lsu/n58 [27], \exu/lsu/n59 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u249  (\exu/data_lsu_uncache [28], \exu/lsu/n58 [28], \exu/lsu/n59 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u25  (\exu/data_lsu_cache [15], \exu/lsu/n64 [15], \exu/lsu/n65 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u250  (\exu/data_lsu_uncache [29], \exu/lsu/n58 [29], \exu/lsu/n59 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u251  (\exu/data_lsu_uncache [30], \exu/lsu/n58 [30], \exu/lsu/n59 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u252  (\exu/data_lsu_uncache [31], \exu/lsu/n58 [31], \exu/lsu/n59 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u253  (\exu/data_lsu_uncache [32], \exu/lsu/n58 [31], \exu/lsu/n59 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u254  (\exu/data_lsu_uncache [33], \exu/lsu/n58 [31], \exu/lsu/n59 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u255  (\exu/data_lsu_uncache [34], \exu/lsu/n58 [31], \exu/lsu/n59 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u256  (\exu/data_lsu_uncache [35], \exu/lsu/n58 [31], \exu/lsu/n59 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u257  (\exu/data_lsu_uncache [36], \exu/lsu/n58 [31], \exu/lsu/n59 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u258  (\exu/data_lsu_uncache [37], \exu/lsu/n58 [31], \exu/lsu/n59 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u259  (\exu/data_lsu_uncache [38], \exu/lsu/n58 [31], \exu/lsu/n59 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u26  (\exu/data_lsu_cache [14], \exu/lsu/n64 [14], \exu/lsu/n65 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u260  (\exu/data_lsu_uncache [39], \exu/lsu/n58 [31], \exu/lsu/n59 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u261  (\exu/data_lsu_uncache [40], \exu/lsu/n58 [31], \exu/lsu/n59 [40]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u262  (\exu/data_lsu_uncache [41], \exu/lsu/n58 [31], \exu/lsu/n59 [41]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u263  (\exu/data_lsu_uncache [42], \exu/lsu/n58 [31], \exu/lsu/n59 [42]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u264  (\exu/data_lsu_uncache [43], \exu/lsu/n58 [31], \exu/lsu/n59 [43]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u265  (\exu/data_lsu_uncache [44], \exu/lsu/n58 [31], \exu/lsu/n59 [44]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u266  (\exu/data_lsu_uncache [45], \exu/lsu/n58 [31], \exu/lsu/n59 [45]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u267  (\exu/data_lsu_uncache [46], \exu/lsu/n58 [31], \exu/lsu/n59 [46]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u268  (\exu/data_lsu_uncache [47], \exu/lsu/n58 [31], \exu/lsu/n59 [47]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u269  (\exu/data_lsu_uncache [48], \exu/lsu/n58 [31], \exu/lsu/n59 [48]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u270  (\exu/data_lsu_uncache [49], \exu/lsu/n58 [31], \exu/lsu/n59 [49]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u271  (\exu/data_lsu_uncache [50], \exu/lsu/n58 [31], \exu/lsu/n59 [50]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u272  (\exu/data_lsu_uncache [51], \exu/lsu/n58 [31], \exu/lsu/n59 [51]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u273  (\exu/data_lsu_uncache [52], \exu/lsu/n58 [31], \exu/lsu/n59 [52]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u274  (\exu/data_lsu_uncache [53], \exu/lsu/n58 [31], \exu/lsu/n59 [53]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u275  (\exu/data_lsu_uncache [54], \exu/lsu/n58 [31], \exu/lsu/n59 [54]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u276  (\exu/data_lsu_uncache [55], \exu/lsu/n58 [31], \exu/lsu/n59 [55]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u277  (\exu/data_lsu_uncache [56], \exu/lsu/n58 [31], \exu/lsu/n59 [56]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u278  (\exu/data_lsu_uncache [57], \exu/lsu/n58 [31], \exu/lsu/n59 [57]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u279  (\exu/data_lsu_uncache [58], \exu/lsu/n58 [31], \exu/lsu/n59 [58]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u28  (\exu/data_lsu_cache [13], \exu/lsu/n64 [13], \exu/lsu/n65 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u280  (\exu/data_lsu_uncache [59], \exu/lsu/n58 [31], \exu/lsu/n59 [59]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u281  (\exu/data_lsu_uncache [60], \exu/lsu/n58 [31], \exu/lsu/n59 [60]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u282  (\exu/data_lsu_uncache [61], \exu/lsu/n58 [31], \exu/lsu/n59 [61]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u283  (\exu/data_lsu_uncache [62], \exu/lsu/n58 [31], \exu/lsu/n59 [62]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u284  (\exu/data_lsu_uncache [63], \exu/lsu/n58 [31], \exu/lsu/n59 [63]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u285  (\exu/lsu/n58 [1], \exu/lsu/n55 [1], \exu/lsu/n57 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u286  (\exu/lsu/n58 [2], \exu/lsu/n55 [2], \exu/lsu/n57 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u287  (\exu/lsu/n58 [3], \exu/lsu/n55 [3], \exu/lsu/n57 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u288  (\exu/lsu/n58 [4], \exu/lsu/n55 [4], \exu/lsu/n57 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u289  (\exu/lsu/n58 [5], \exu/lsu/n55 [5], \exu/lsu/n57 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u29  (\exu/lsu/n38 [0], \exu/lsu/n36 [0], \exu/lsu/n37 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u290  (\exu/lsu/n58 [6], \exu/lsu/n55 [6], \exu/lsu/n57 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u291  (\exu/lsu/n58 [7], \exu/lsu/n55 [7], \exu/lsu/n57 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u292  (\exu/lsu/n58 [8], \exu/lsu/n55 [8], \exu/lsu/n57 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u293  (\exu/lsu/n58 [9], \exu/lsu/n55 [9], \exu/lsu/n57 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u294  (\exu/lsu/n58 [10], \exu/lsu/n55 [10], \exu/lsu/n57 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u295  (\exu/lsu/n58 [11], \exu/lsu/n55 [11], \exu/lsu/n57 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u296  (\exu/lsu/n58 [12], \exu/lsu/n55 [12], \exu/lsu/n57 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u297  (\exu/lsu/n58 [13], \exu/lsu/n55 [13], \exu/lsu/n57 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u298  (\exu/lsu/n58 [14], \exu/lsu/n55 [14], \exu/lsu/n57 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u299  (\exu/lsu/n58 [15], \exu/lsu/n55 [15], \exu/lsu/n57 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u3  (\exu/data_lsu_cache [24], \exu/lsu/n64 [24], \exu/lsu/n65 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u30  (\exu/data_lsu_cache [12], \exu/lsu/n64 [12], \exu/lsu/n65 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u300  (\exu/lsu/n58 [16], \exu/lsu/n55 [15], \exu/lsu/n57 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u301  (\exu/lsu/n58 [17], \exu/lsu/n55 [15], \exu/lsu/n57 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u302  (\exu/lsu/n58 [18], \exu/lsu/n55 [15], \exu/lsu/n57 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u303  (\exu/lsu/n58 [19], \exu/lsu/n55 [15], \exu/lsu/n57 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u304  (\exu/lsu/n58 [20], \exu/lsu/n55 [15], \exu/lsu/n57 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u305  (\exu/lsu/n58 [21], \exu/lsu/n55 [15], \exu/lsu/n57 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u306  (\exu/lsu/n58 [22], \exu/lsu/n55 [15], \exu/lsu/n57 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u307  (\exu/lsu/n58 [23], \exu/lsu/n55 [15], \exu/lsu/n57 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u308  (\exu/lsu/n58 [24], \exu/lsu/n55 [15], \exu/lsu/n57 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u309  (\exu/lsu/n58 [25], \exu/lsu/n55 [15], \exu/lsu/n57 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u31  (\exu/lsu/n40 [0], \exu/lsu/n38 [0], \exu/lsu/n39 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u310  (\exu/lsu/n58 [26], \exu/lsu/n55 [15], \exu/lsu/n57 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u311  (\exu/lsu/n58 [27], \exu/lsu/n55 [15], \exu/lsu/n57 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u312  (\exu/lsu/n58 [28], \exu/lsu/n55 [15], \exu/lsu/n57 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u313  (\exu/lsu/n58 [29], \exu/lsu/n55 [15], \exu/lsu/n57 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u314  (\exu/lsu/n58 [30], \exu/lsu/n55 [15], \exu/lsu/n57 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u315  (\exu/lsu/n58 [31], \exu/lsu/n55 [15], \exu/lsu/n57 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u32  (\exu/data_lsu_cache [11], \exu/lsu/n64 [11], \exu/lsu/n65 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u33  (\exu/lsu/n42 [0], \exu/lsu/n40 [0], \exu/lsu/n41 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u34  (\exu/data_lsu_cache [10], \exu/lsu/n64 [10], \exu/lsu/n65 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u348  (\exu/lsu/n55 [1], \exu/lsu/n52 [1], \exu/lsu/n54 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u349  (\exu/lsu/n55 [2], \exu/lsu/n52 [2], \exu/lsu/n54 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u350  (\exu/lsu/n55 [3], \exu/lsu/n52 [3], \exu/lsu/n54 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u351  (\exu/lsu/n55 [4], \exu/lsu/n52 [4], \exu/lsu/n54 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u352  (\exu/lsu/n55 [5], \exu/lsu/n52 [5], \exu/lsu/n54 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u353  (\exu/lsu/n55 [6], \exu/lsu/n52 [6], \exu/lsu/n54 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u354  (\exu/lsu/n55 [7], \exu/lsu/n52 [10], \exu/lsu/n54 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u355  (\exu/lsu/n55 [8], \exu/lsu/n52 [10], \exu/lsu/n54 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u356  (\exu/lsu/n55 [9], \exu/lsu/n52 [10], \exu/lsu/n54 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u357  (\exu/lsu/n55 [10], \exu/lsu/n52 [10], \exu/lsu/n54 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u358  (\exu/lsu/n55 [11], \exu/lsu/n52 [10], \exu/lsu/n54 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u359  (\exu/lsu/n55 [12], \exu/lsu/n52 [10], \exu/lsu/n54 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u36  (\exu/data_lsu_cache [9], \exu/lsu/n64 [9], \exu/lsu/n65 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u360  (\exu/lsu/n55 [13], \exu/lsu/n52 [10], \exu/lsu/n54 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u361  (\exu/lsu/n55 [14], \exu/lsu/n52 [10], \exu/lsu/n54 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u362  (\exu/lsu/n55 [15], \exu/lsu/n52 [10], \exu/lsu/n54 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u38  (\exu/data_lsu_cache [8], \exu/lsu/n64 [8], \exu/lsu/n65 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  and \exu/lsu/u41  (\exu/lsu/n51 , ex_size[0], \exu/alu_au/n0 );  // ../../RTL/CPU/EX/LSU/lsu.v(61)
  or \exu/lsu/u42  (\exu/data_lsu_cache [7], \exu/lsu/n64 [7], \exu/lsu/n65 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  and \exu/lsu/u43  (\exu/lsu/n53 , ex_size[1], \exu/alu_au/n0 );  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u45  (\exu/data_lsu_cache [6], \exu/lsu/n64 [6], \exu/lsu/n65 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  and \exu/lsu/u46  (\exu/lsu/n56 , ex_size[2], \exu/alu_au/n0 );  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u47  (\exu/lsu/n55 [0], \exu/lsu/n52 [0], \exu/lsu/n54 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(62)
  or \exu/lsu/u48  (\exu/lsu/n58 [0], \exu/lsu/n55 [0], \exu/lsu/n57 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(63)
  or \exu/lsu/u487  (\exu/lsu/n42 [1], \exu/lsu/n40 [1], \exu/lsu/n41 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u488  (\exu/lsu/n42 [2], \exu/lsu/n40 [2], \exu/lsu/n41 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u489  (\exu/lsu/n42 [3], \exu/lsu/n40 [3], \exu/lsu/n41 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u49  (\exu/data_lsu_cache [5], \exu/lsu/n64 [5], \exu/lsu/n65 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u490  (\exu/lsu/n42 [4], \exu/lsu/n40 [4], \exu/lsu/n41 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u491  (\exu/lsu/n42 [5], \exu/lsu/n40 [5], \exu/lsu/n41 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u492  (\exu/lsu/n42 [6], \exu/lsu/n40 [6], \exu/lsu/n41 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u493  (\exu/lsu/n42 [7], \exu/lsu/n40 [7], \exu/lsu/n41 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u494  (\exu/lsu/n42 [8], \exu/lsu/n40 [8], \exu/lsu/n41 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u495  (\exu/lsu/n42 [9], \exu/lsu/n40 [9], \exu/lsu/n41 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u496  (\exu/lsu/n42 [10], \exu/lsu/n40 [10], \exu/lsu/n41 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u497  (\exu/lsu/n42 [11], \exu/lsu/n40 [11], \exu/lsu/n41 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u498  (\exu/lsu/n42 [12], \exu/lsu/n40 [12], \exu/lsu/n41 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u499  (\exu/lsu/n42 [13], \exu/lsu/n40 [13], \exu/lsu/n41 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u50  (\exu/data_lsu_cache [4], \exu/lsu/n64 [4], \exu/lsu/n65 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u500  (\exu/lsu/n42 [14], \exu/lsu/n40 [14], \exu/lsu/n41 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u501  (\exu/lsu/n42 [15], \exu/lsu/n40 [15], \exu/lsu/n41 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u502  (\exu/lsu/n42 [16], \exu/lsu/n40 [16], \exu/lsu/n41 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u503  (\exu/lsu/n42 [17], \exu/lsu/n40 [17], \exu/lsu/n41 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u504  (\exu/lsu/n42 [18], \exu/lsu/n40 [18], \exu/lsu/n41 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u505  (\exu/lsu/n42 [19], \exu/lsu/n40 [19], \exu/lsu/n41 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u506  (\exu/lsu/n42 [20], \exu/lsu/n40 [20], \exu/lsu/n41 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u507  (\exu/lsu/n42 [21], \exu/lsu/n40 [21], \exu/lsu/n41 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u508  (\exu/lsu/n42 [22], \exu/lsu/n40 [22], \exu/lsu/n41 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u509  (\exu/lsu/n42 [23], \exu/lsu/n40 [23], \exu/lsu/n41 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u51  (\exu/data_lsu_cache [3], \exu/lsu/n64 [3], \exu/lsu/n65 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u510  (\exu/lsu/n42 [24], \exu/lsu/n40 [24], \exu/lsu/n41 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u511  (\exu/lsu/n42 [25], \exu/lsu/n40 [25], \exu/lsu/n41 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u512  (\exu/lsu/n42 [26], \exu/lsu/n40 [26], \exu/lsu/n41 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u513  (\exu/lsu/n42 [27], \exu/lsu/n40 [27], \exu/lsu/n41 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u514  (\exu/lsu/n42 [28], \exu/lsu/n40 [28], \exu/lsu/n41 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u515  (\exu/lsu/n42 [29], \exu/lsu/n40 [29], \exu/lsu/n41 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u516  (\exu/lsu/n42 [30], \exu/lsu/n40 [30], \exu/lsu/n41 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u517  (\exu/lsu/n42 [31], \exu/lsu/n40 [31], \exu/lsu/n41 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u518  (\exu/lsu/data_lsu_cache_shift [32], \exu/lsu/n40 [32], \exu/lsu/n41 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u519  (\exu/lsu/data_lsu_cache_shift [33], \exu/lsu/n40 [33], \exu/lsu/n41 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u52  (\exu/data_lsu_cache [2], \exu/lsu/n64 [2], \exu/lsu/n65 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u520  (\exu/lsu/data_lsu_cache_shift [34], \exu/lsu/n40 [34], \exu/lsu/n41 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u521  (\exu/lsu/data_lsu_cache_shift [35], \exu/lsu/n40 [35], \exu/lsu/n41 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u522  (\exu/lsu/data_lsu_cache_shift [36], \exu/lsu/n40 [36], \exu/lsu/n41 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u523  (\exu/lsu/data_lsu_cache_shift [37], \exu/lsu/n40 [37], \exu/lsu/n41 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u524  (\exu/lsu/data_lsu_cache_shift [38], \exu/lsu/n40 [38], \exu/lsu/n41 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u525  (\exu/lsu/data_lsu_cache_shift [39], \exu/lsu/n40 [39], \exu/lsu/n41 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(54)
  or \exu/lsu/u526  (\exu/lsu/n40 [1], \exu/lsu/n38 [1], \exu/lsu/n39 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u527  (\exu/lsu/n40 [2], \exu/lsu/n38 [2], \exu/lsu/n39 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u528  (\exu/lsu/n40 [3], \exu/lsu/n38 [3], \exu/lsu/n39 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u529  (\exu/lsu/n40 [4], \exu/lsu/n38 [4], \exu/lsu/n39 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u53  (\exu/data_lsu_uncache [0], \exu/lsu/n58 [0], \exu/lsu/n59 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(64)
  or \exu/lsu/u530  (\exu/lsu/n40 [5], \exu/lsu/n38 [5], \exu/lsu/n39 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u531  (\exu/lsu/n40 [6], \exu/lsu/n38 [6], \exu/lsu/n39 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u532  (\exu/lsu/n40 [7], \exu/lsu/n38 [7], \exu/lsu/n39 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u533  (\exu/lsu/n40 [8], \exu/lsu/n38 [8], \exu/lsu/n39 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u534  (\exu/lsu/n40 [9], \exu/lsu/n38 [9], \exu/lsu/n39 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u535  (\exu/lsu/n40 [10], \exu/lsu/n38 [10], \exu/lsu/n39 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u536  (\exu/lsu/n40 [11], \exu/lsu/n38 [11], \exu/lsu/n39 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u537  (\exu/lsu/n40 [12], \exu/lsu/n38 [12], \exu/lsu/n39 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u538  (\exu/lsu/n40 [13], \exu/lsu/n38 [13], \exu/lsu/n39 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u539  (\exu/lsu/n40 [14], \exu/lsu/n38 [14], \exu/lsu/n39 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u54  (\exu/data_lsu_cache [1], \exu/lsu/n64 [1], \exu/lsu/n65 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u540  (\exu/lsu/n40 [15], \exu/lsu/n38 [15], \exu/lsu/n39 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u541  (\exu/lsu/n40 [16], \exu/lsu/n38 [16], \exu/lsu/n39 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u542  (\exu/lsu/n40 [17], \exu/lsu/n38 [17], \exu/lsu/n39 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u543  (\exu/lsu/n40 [18], \exu/lsu/n38 [18], \exu/lsu/n39 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u544  (\exu/lsu/n40 [19], \exu/lsu/n38 [19], \exu/lsu/n39 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u545  (\exu/lsu/n40 [20], \exu/lsu/n38 [20], \exu/lsu/n39 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u546  (\exu/lsu/n40 [21], \exu/lsu/n38 [21], \exu/lsu/n39 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u547  (\exu/lsu/n40 [22], \exu/lsu/n38 [22], \exu/lsu/n39 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u548  (\exu/lsu/n40 [23], \exu/lsu/n38 [23], \exu/lsu/n39 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u549  (\exu/lsu/n40 [24], \exu/lsu/n38 [24], \exu/lsu/n39 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u55  (\exu/data_lsu_cache [0], \exu/lsu/n64 [0], \exu/lsu/n65 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u550  (\exu/lsu/n40 [25], \exu/lsu/n38 [25], \exu/lsu/n39 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u551  (\exu/lsu/n40 [26], \exu/lsu/n38 [26], \exu/lsu/n39 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u552  (\exu/lsu/n40 [27], \exu/lsu/n38 [27], \exu/lsu/n39 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u553  (\exu/lsu/n40 [28], \exu/lsu/n38 [28], \exu/lsu/n39 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u554  (\exu/lsu/n40 [29], \exu/lsu/n38 [29], \exu/lsu/n39 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u555  (\exu/lsu/n40 [30], \exu/lsu/n38 [30], \exu/lsu/n39 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u556  (\exu/lsu/n40 [31], \exu/lsu/n38 [31], \exu/lsu/n39 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u557  (\exu/lsu/n40 [32], \exu/lsu/n38 [32], \exu/lsu/n39 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u558  (\exu/lsu/n40 [33], \exu/lsu/n38 [33], \exu/lsu/n39 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u559  (\exu/lsu/n40 [34], \exu/lsu/n38 [34], \exu/lsu/n39 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u56  (\exu/lsu/n62 [0], \exu/lsu/n60 [0], \exu/lsu/n61 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(68)
  or \exu/lsu/u560  (\exu/lsu/n40 [35], \exu/lsu/n38 [35], \exu/lsu/n39 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u561  (\exu/lsu/n40 [36], \exu/lsu/n38 [36], \exu/lsu/n39 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u562  (\exu/lsu/n40 [37], \exu/lsu/n38 [37], \exu/lsu/n39 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u563  (\exu/lsu/n40 [38], \exu/lsu/n38 [38], \exu/lsu/n39 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u564  (\exu/lsu/n40 [39], \exu/lsu/n38 [39], \exu/lsu/n39 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u565  (\exu/lsu/data_lsu_cache_shift [40], \exu/lsu/n38 [40], \exu/lsu/n39 [40]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u566  (\exu/lsu/data_lsu_cache_shift [41], \exu/lsu/n38 [41], \exu/lsu/n39 [41]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u567  (\exu/lsu/data_lsu_cache_shift [42], \exu/lsu/n38 [42], \exu/lsu/n39 [42]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u568  (\exu/lsu/data_lsu_cache_shift [43], \exu/lsu/n38 [43], \exu/lsu/n39 [43]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u569  (\exu/lsu/data_lsu_cache_shift [44], \exu/lsu/n38 [44], \exu/lsu/n39 [44]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u57  (\exu/lsu/n64 [0], \exu/lsu/n62 [0], \exu/lsu/n63 [0]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u570  (\exu/lsu/data_lsu_cache_shift [45], \exu/lsu/n38 [45], \exu/lsu/n39 [45]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u571  (\exu/lsu/data_lsu_cache_shift [46], \exu/lsu/n38 [46], \exu/lsu/n39 [46]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u572  (\exu/lsu/data_lsu_cache_shift [47], \exu/lsu/n38 [47], \exu/lsu/n39 [47]);  // ../../RTL/CPU/EX/LSU/lsu.v(53)
  or \exu/lsu/u573  (\exu/lsu/n38 [1], \exu/lsu/n36 [1], \exu/lsu/n37 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u574  (\exu/lsu/n38 [2], \exu/lsu/n36 [2], \exu/lsu/n37 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u575  (\exu/lsu/n38 [3], \exu/lsu/n36 [3], \exu/lsu/n37 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u576  (\exu/lsu/n38 [4], \exu/lsu/n36 [4], \exu/lsu/n37 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u577  (\exu/lsu/n38 [5], \exu/lsu/n36 [5], \exu/lsu/n37 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u578  (\exu/lsu/n38 [6], \exu/lsu/n36 [6], \exu/lsu/n37 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u579  (\exu/lsu/n38 [7], \exu/lsu/n36 [7], \exu/lsu/n37 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u58  (\exu/data_lsu_cache [26], \exu/lsu/n64 [26], \exu/lsu/n65 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u580  (\exu/lsu/n38 [8], \exu/lsu/n36 [8], \exu/lsu/n37 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u581  (\exu/lsu/n38 [9], \exu/lsu/n36 [9], \exu/lsu/n37 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u582  (\exu/lsu/n38 [10], \exu/lsu/n36 [10], \exu/lsu/n37 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u583  (\exu/lsu/n38 [11], \exu/lsu/n36 [11], \exu/lsu/n37 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u584  (\exu/lsu/n38 [12], \exu/lsu/n36 [12], \exu/lsu/n37 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u585  (\exu/lsu/n38 [13], \exu/lsu/n36 [13], \exu/lsu/n37 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u586  (\exu/lsu/n38 [14], \exu/lsu/n36 [14], \exu/lsu/n37 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u587  (\exu/lsu/n38 [15], \exu/lsu/n36 [15], \exu/lsu/n37 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u588  (\exu/lsu/n38 [16], \exu/lsu/n36 [16], \exu/lsu/n37 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u589  (\exu/lsu/n38 [17], \exu/lsu/n36 [17], \exu/lsu/n37 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u59  (\exu/data_lsu_cache [27], \exu/lsu/n64 [27], \exu/lsu/n65 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u590  (\exu/lsu/n38 [18], \exu/lsu/n36 [18], \exu/lsu/n37 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u591  (\exu/lsu/n38 [19], \exu/lsu/n36 [19], \exu/lsu/n37 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u592  (\exu/lsu/n38 [20], \exu/lsu/n36 [20], \exu/lsu/n37 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u593  (\exu/lsu/n38 [21], \exu/lsu/n36 [21], \exu/lsu/n37 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u594  (\exu/lsu/n38 [22], \exu/lsu/n36 [22], \exu/lsu/n37 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u595  (\exu/lsu/n38 [23], \exu/lsu/n36 [23], \exu/lsu/n37 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u596  (\exu/lsu/n38 [24], \exu/lsu/n36 [24], \exu/lsu/n37 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u597  (\exu/lsu/n38 [25], \exu/lsu/n36 [25], \exu/lsu/n37 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u598  (\exu/lsu/n38 [26], \exu/lsu/n36 [26], \exu/lsu/n37 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u599  (\exu/lsu/n38 [27], \exu/lsu/n36 [27], \exu/lsu/n37 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u60  (\exu/data_lsu_cache [28], \exu/lsu/n64 [28], \exu/lsu/n65 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u600  (\exu/lsu/n38 [28], \exu/lsu/n36 [28], \exu/lsu/n37 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u601  (\exu/lsu/n38 [29], \exu/lsu/n36 [29], \exu/lsu/n37 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u602  (\exu/lsu/n38 [30], \exu/lsu/n36 [30], \exu/lsu/n37 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u603  (\exu/lsu/n38 [31], \exu/lsu/n36 [31], \exu/lsu/n37 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u604  (\exu/lsu/n38 [32], \exu/lsu/n36 [32], \exu/lsu/n37 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u605  (\exu/lsu/n38 [33], \exu/lsu/n36 [33], \exu/lsu/n37 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u606  (\exu/lsu/n38 [34], \exu/lsu/n36 [34], \exu/lsu/n37 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u607  (\exu/lsu/n38 [35], \exu/lsu/n36 [35], \exu/lsu/n37 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u608  (\exu/lsu/n38 [36], \exu/lsu/n36 [36], \exu/lsu/n37 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u609  (\exu/lsu/n38 [37], \exu/lsu/n36 [37], \exu/lsu/n37 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u61  (\exu/data_lsu_cache [29], \exu/lsu/n64 [29], \exu/lsu/n65 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u610  (\exu/lsu/n38 [38], \exu/lsu/n36 [38], \exu/lsu/n37 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u611  (\exu/lsu/n38 [39], \exu/lsu/n36 [39], \exu/lsu/n37 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u612  (\exu/lsu/n38 [40], \exu/lsu/n36 [40], \exu/lsu/n37 [40]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u613  (\exu/lsu/n38 [41], \exu/lsu/n36 [41], \exu/lsu/n37 [41]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u614  (\exu/lsu/n38 [42], \exu/lsu/n36 [42], \exu/lsu/n37 [42]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u615  (\exu/lsu/n38 [43], \exu/lsu/n36 [43], \exu/lsu/n37 [43]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u616  (\exu/lsu/n38 [44], \exu/lsu/n36 [44], \exu/lsu/n37 [44]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u617  (\exu/lsu/n38 [45], \exu/lsu/n36 [45], \exu/lsu/n37 [45]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u618  (\exu/lsu/n38 [46], \exu/lsu/n36 [46], \exu/lsu/n37 [46]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u619  (\exu/lsu/n38 [47], \exu/lsu/n36 [47], \exu/lsu/n37 [47]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u62  (\exu/data_lsu_cache [30], \exu/lsu/n64 [30], \exu/lsu/n65 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u620  (\exu/lsu/data_lsu_cache_shift [48], \exu/lsu/n36 [48], \exu/lsu/n37 [48]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u621  (\exu/lsu/data_lsu_cache_shift [49], \exu/lsu/n36 [49], \exu/lsu/n37 [49]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u622  (\exu/lsu/data_lsu_cache_shift [50], \exu/lsu/n36 [50], \exu/lsu/n37 [50]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u623  (\exu/lsu/data_lsu_cache_shift [51], \exu/lsu/n36 [51], \exu/lsu/n37 [51]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u624  (\exu/lsu/data_lsu_cache_shift [52], \exu/lsu/n36 [52], \exu/lsu/n37 [52]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u625  (\exu/lsu/data_lsu_cache_shift [53], \exu/lsu/n36 [53], \exu/lsu/n37 [53]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u626  (\exu/lsu/data_lsu_cache_shift [54], \exu/lsu/n36 [54], \exu/lsu/n37 [54]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u627  (\exu/lsu/data_lsu_cache_shift [55], \exu/lsu/n36 [55], \exu/lsu/n37 [55]);  // ../../RTL/CPU/EX/LSU/lsu.v(52)
  or \exu/lsu/u63  (\exu/data_lsu_cache [31], \exu/lsu/n64 [31], \exu/lsu/n65 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u64  (\exu/data_lsu_cache [32], \exu/lsu/n64 [31], \exu/lsu/n65 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u65  (\exu/data_lsu_cache [33], \exu/lsu/n64 [31], \exu/lsu/n65 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u66  (\exu/data_lsu_cache [34], \exu/lsu/n64 [31], \exu/lsu/n65 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u67  (\exu/data_lsu_cache [35], \exu/lsu/n64 [31], \exu/lsu/n65 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u68  (\exu/data_lsu_cache [36], \exu/lsu/n64 [31], \exu/lsu/n65 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u69  (\exu/data_lsu_cache [37], \exu/lsu/n64 [31], \exu/lsu/n65 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u70  (\exu/data_lsu_cache [38], \exu/lsu/n64 [31], \exu/lsu/n65 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u704  (\exu/lsu/n28 [1], \exu/lsu/n26 [1], \exu/lsu/n27 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u705  (\exu/lsu/n28 [2], \exu/lsu/n26 [2], \exu/lsu/n27 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u706  (\exu/lsu/n28 [3], \exu/lsu/n26 [3], \exu/lsu/n27 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u707  (\exu/lsu/n28 [4], \exu/lsu/n26 [4], \exu/lsu/n27 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u708  (\exu/lsu/n28 [5], \exu/lsu/n26 [5], \exu/lsu/n27 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u709  (\exu/lsu/n28 [6], \exu/lsu/n26 [6], \exu/lsu/n27 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u71  (\exu/data_lsu_cache [39], \exu/lsu/n64 [31], \exu/lsu/n65 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u710  (\exu/lsu/n28 [7], \exu/lsu/n26 [7], \exu/lsu/n27 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u711  (\exu/lsu/n28 [8], \exu/lsu/n26 [8], \exu/lsu/n27 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u712  (\exu/lsu/n28 [9], \exu/lsu/n26 [9], \exu/lsu/n27 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u713  (\exu/lsu/n28 [10], \exu/lsu/n26 [10], \exu/lsu/n27 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u714  (\exu/lsu/n28 [11], \exu/lsu/n26 [11], \exu/lsu/n27 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u715  (\exu/lsu/n28 [12], \exu/lsu/n26 [12], \exu/lsu/n27 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u716  (\exu/lsu/n28 [13], \exu/lsu/n26 [13], \exu/lsu/n27 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u717  (\exu/lsu/n28 [14], \exu/lsu/n26 [14], \exu/lsu/n27 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u718  (\exu/lsu/n28 [15], \exu/lsu/n26 [15], \exu/lsu/n27 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u719  (\exu/lsu/n28 [16], \exu/lsu/n26 [16], \exu/lsu/n27 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u72  (\exu/data_lsu_cache [40], \exu/lsu/n64 [31], \exu/lsu/n65 [40]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u720  (\exu/lsu/n28 [17], \exu/lsu/n26 [17], \exu/lsu/n27 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u721  (\exu/lsu/n28 [18], \exu/lsu/n26 [18], \exu/lsu/n27 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u722  (\exu/lsu/n28 [19], \exu/lsu/n26 [19], \exu/lsu/n27 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u723  (\exu/lsu/n28 [20], \exu/lsu/n26 [20], \exu/lsu/n27 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u724  (\exu/lsu/n28 [21], \exu/lsu/n26 [21], \exu/lsu/n27 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u725  (\exu/lsu/n28 [22], \exu/lsu/n26 [22], \exu/lsu/n27 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u726  (\exu/lsu/n28 [23], \exu/lsu/n26 [23], \exu/lsu/n27 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u727  (\exu/lsu/n28 [24], \exu/lsu/n26 [24], \exu/lsu/n27 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u728  (\exu/lsu/n28 [25], \exu/lsu/n26 [25], \exu/lsu/n27 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u729  (\exu/lsu/n28 [26], \exu/lsu/n26 [26], \exu/lsu/n27 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u73  (\exu/data_lsu_cache [41], \exu/lsu/n64 [31], \exu/lsu/n65 [41]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u730  (\exu/lsu/n28 [27], \exu/lsu/n26 [27], \exu/lsu/n27 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u731  (\exu/lsu/n28 [28], \exu/lsu/n26 [28], \exu/lsu/n27 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u732  (\exu/lsu/n28 [29], \exu/lsu/n26 [29], \exu/lsu/n27 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u733  (\exu/lsu/n28 [30], \exu/lsu/n26 [30], \exu/lsu/n27 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u734  (\exu/lsu/n28 [31], \exu/lsu/n26 [31], \exu/lsu/n27 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u735  (\exu/lsu/data_lsu_uncache_shift [32], \exu/lsu/n26 [32], \exu/lsu/n27 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u736  (\exu/lsu/data_lsu_uncache_shift [33], \exu/lsu/n26 [33], \exu/lsu/n27 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u737  (\exu/lsu/data_lsu_uncache_shift [34], \exu/lsu/n26 [34], \exu/lsu/n27 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u738  (\exu/lsu/data_lsu_uncache_shift [35], \exu/lsu/n26 [35], \exu/lsu/n27 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u739  (\exu/lsu/data_lsu_uncache_shift [36], \exu/lsu/n26 [36], \exu/lsu/n27 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u74  (\exu/data_lsu_cache [42], \exu/lsu/n64 [31], \exu/lsu/n65 [42]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u740  (\exu/lsu/data_lsu_uncache_shift [37], \exu/lsu/n26 [37], \exu/lsu/n27 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u741  (\exu/lsu/data_lsu_uncache_shift [38], \exu/lsu/n26 [38], \exu/lsu/n27 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u742  (\exu/lsu/data_lsu_uncache_shift [39], \exu/lsu/n26 [39], \exu/lsu/n27 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(45)
  or \exu/lsu/u743  (\exu/lsu/n26 [1], \exu/lsu/n24 [1], \exu/lsu/n25 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u744  (\exu/lsu/n26 [2], \exu/lsu/n24 [2], \exu/lsu/n25 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u745  (\exu/lsu/n26 [3], \exu/lsu/n24 [3], \exu/lsu/n25 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u746  (\exu/lsu/n26 [4], \exu/lsu/n24 [4], \exu/lsu/n25 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u747  (\exu/lsu/n26 [5], \exu/lsu/n24 [5], \exu/lsu/n25 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u748  (\exu/lsu/n26 [6], \exu/lsu/n24 [6], \exu/lsu/n25 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u749  (\exu/lsu/n26 [7], \exu/lsu/n24 [7], \exu/lsu/n25 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u75  (\exu/data_lsu_cache [43], \exu/lsu/n64 [31], \exu/lsu/n65 [43]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u750  (\exu/lsu/n26 [8], \exu/lsu/n24 [8], \exu/lsu/n25 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u751  (\exu/lsu/n26 [9], \exu/lsu/n24 [9], \exu/lsu/n25 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u752  (\exu/lsu/n26 [10], \exu/lsu/n24 [10], \exu/lsu/n25 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u753  (\exu/lsu/n26 [11], \exu/lsu/n24 [11], \exu/lsu/n25 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u754  (\exu/lsu/n26 [12], \exu/lsu/n24 [12], \exu/lsu/n25 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u755  (\exu/lsu/n26 [13], \exu/lsu/n24 [13], \exu/lsu/n25 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u756  (\exu/lsu/n26 [14], \exu/lsu/n24 [14], \exu/lsu/n25 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u757  (\exu/lsu/n26 [15], \exu/lsu/n24 [15], \exu/lsu/n25 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u758  (\exu/lsu/n26 [16], \exu/lsu/n24 [16], \exu/lsu/n25 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u759  (\exu/lsu/n26 [17], \exu/lsu/n24 [17], \exu/lsu/n25 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u76  (\exu/data_lsu_cache [44], \exu/lsu/n64 [31], \exu/lsu/n65 [44]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u760  (\exu/lsu/n26 [18], \exu/lsu/n24 [18], \exu/lsu/n25 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u761  (\exu/lsu/n26 [19], \exu/lsu/n24 [19], \exu/lsu/n25 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u762  (\exu/lsu/n26 [20], \exu/lsu/n24 [20], \exu/lsu/n25 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u763  (\exu/lsu/n26 [21], \exu/lsu/n24 [21], \exu/lsu/n25 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u764  (\exu/lsu/n26 [22], \exu/lsu/n24 [22], \exu/lsu/n25 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u765  (\exu/lsu/n26 [23], \exu/lsu/n24 [23], \exu/lsu/n25 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u766  (\exu/lsu/n26 [24], \exu/lsu/n24 [24], \exu/lsu/n25 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u767  (\exu/lsu/n26 [25], \exu/lsu/n24 [25], \exu/lsu/n25 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u768  (\exu/lsu/n26 [26], \exu/lsu/n24 [26], \exu/lsu/n25 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u769  (\exu/lsu/n26 [27], \exu/lsu/n24 [27], \exu/lsu/n25 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u77  (\exu/data_lsu_cache [45], \exu/lsu/n64 [31], \exu/lsu/n65 [45]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u770  (\exu/lsu/n26 [28], \exu/lsu/n24 [28], \exu/lsu/n25 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u771  (\exu/lsu/n26 [29], \exu/lsu/n24 [29], \exu/lsu/n25 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u772  (\exu/lsu/n26 [30], \exu/lsu/n24 [30], \exu/lsu/n25 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u773  (\exu/lsu/n26 [31], \exu/lsu/n24 [31], \exu/lsu/n25 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u774  (\exu/lsu/n26 [32], \exu/lsu/n24 [32], \exu/lsu/n25 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u775  (\exu/lsu/n26 [33], \exu/lsu/n24 [33], \exu/lsu/n25 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u776  (\exu/lsu/n26 [34], \exu/lsu/n24 [34], \exu/lsu/n25 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u777  (\exu/lsu/n26 [35], \exu/lsu/n24 [35], \exu/lsu/n25 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u778  (\exu/lsu/n26 [36], \exu/lsu/n24 [36], \exu/lsu/n25 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u779  (\exu/lsu/n26 [37], \exu/lsu/n24 [37], \exu/lsu/n25 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u78  (\exu/data_lsu_cache [46], \exu/lsu/n64 [31], \exu/lsu/n65 [46]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u780  (\exu/lsu/n26 [38], \exu/lsu/n24 [38], \exu/lsu/n25 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u781  (\exu/lsu/n26 [39], \exu/lsu/n24 [39], \exu/lsu/n25 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u782  (\exu/lsu/data_lsu_uncache_shift [40], \exu/lsu/n24 [40], \exu/lsu/n25 [40]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u783  (\exu/lsu/data_lsu_uncache_shift [41], \exu/lsu/n24 [41], \exu/lsu/n25 [41]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u784  (\exu/lsu/data_lsu_uncache_shift [42], \exu/lsu/n24 [42], \exu/lsu/n25 [42]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u785  (\exu/lsu/data_lsu_uncache_shift [43], \exu/lsu/n24 [43], \exu/lsu/n25 [43]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u786  (\exu/lsu/data_lsu_uncache_shift [44], \exu/lsu/n24 [44], \exu/lsu/n25 [44]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u787  (\exu/lsu/data_lsu_uncache_shift [45], \exu/lsu/n24 [45], \exu/lsu/n25 [45]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u788  (\exu/lsu/data_lsu_uncache_shift [46], \exu/lsu/n24 [46], \exu/lsu/n25 [46]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u789  (\exu/lsu/data_lsu_uncache_shift [47], \exu/lsu/n24 [47], \exu/lsu/n25 [47]);  // ../../RTL/CPU/EX/LSU/lsu.v(44)
  or \exu/lsu/u79  (\exu/data_lsu_cache [47], \exu/lsu/n64 [31], \exu/lsu/n65 [47]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u790  (\exu/lsu/n24 [1], \exu/lsu/n22 [1], \exu/lsu/n23 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u791  (\exu/lsu/n24 [2], \exu/lsu/n22 [2], \exu/lsu/n23 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u792  (\exu/lsu/n24 [3], \exu/lsu/n22 [3], \exu/lsu/n23 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u793  (\exu/lsu/n24 [4], \exu/lsu/n22 [4], \exu/lsu/n23 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u794  (\exu/lsu/n24 [5], \exu/lsu/n22 [5], \exu/lsu/n23 [5]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u795  (\exu/lsu/n24 [6], \exu/lsu/n22 [6], \exu/lsu/n23 [6]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u796  (\exu/lsu/n24 [7], \exu/lsu/n22 [7], \exu/lsu/n23 [7]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u797  (\exu/lsu/n24 [8], \exu/lsu/n22 [8], \exu/lsu/n23 [8]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u798  (\exu/lsu/n24 [9], \exu/lsu/n22 [9], \exu/lsu/n23 [9]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u799  (\exu/lsu/n24 [10], \exu/lsu/n22 [10], \exu/lsu/n23 [10]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u80  (\exu/data_lsu_cache [48], \exu/lsu/n64 [31], \exu/lsu/n65 [48]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u800  (\exu/lsu/n24 [11], \exu/lsu/n22 [11], \exu/lsu/n23 [11]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u801  (\exu/lsu/n24 [12], \exu/lsu/n22 [12], \exu/lsu/n23 [12]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u802  (\exu/lsu/n24 [13], \exu/lsu/n22 [13], \exu/lsu/n23 [13]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u803  (\exu/lsu/n24 [14], \exu/lsu/n22 [14], \exu/lsu/n23 [14]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u804  (\exu/lsu/n24 [15], \exu/lsu/n22 [15], \exu/lsu/n23 [15]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u805  (\exu/lsu/n24 [16], \exu/lsu/n22 [16], \exu/lsu/n23 [16]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u806  (\exu/lsu/n24 [17], \exu/lsu/n22 [17], \exu/lsu/n23 [17]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u807  (\exu/lsu/n24 [18], \exu/lsu/n22 [18], \exu/lsu/n23 [18]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u808  (\exu/lsu/n24 [19], \exu/lsu/n22 [19], \exu/lsu/n23 [19]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u809  (\exu/lsu/n24 [20], \exu/lsu/n22 [20], \exu/lsu/n23 [20]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u81  (\exu/data_lsu_cache [49], \exu/lsu/n64 [31], \exu/lsu/n65 [49]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u810  (\exu/lsu/n24 [21], \exu/lsu/n22 [21], \exu/lsu/n23 [21]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u811  (\exu/lsu/n24 [22], \exu/lsu/n22 [22], \exu/lsu/n23 [22]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u812  (\exu/lsu/n24 [23], \exu/lsu/n22 [23], \exu/lsu/n23 [23]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u813  (\exu/lsu/n24 [24], \exu/lsu/n22 [24], \exu/lsu/n23 [24]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u814  (\exu/lsu/n24 [25], \exu/lsu/n22 [25], \exu/lsu/n23 [25]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u815  (\exu/lsu/n24 [26], \exu/lsu/n22 [26], \exu/lsu/n23 [26]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u816  (\exu/lsu/n24 [27], \exu/lsu/n22 [27], \exu/lsu/n23 [27]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u817  (\exu/lsu/n24 [28], \exu/lsu/n22 [28], \exu/lsu/n23 [28]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u818  (\exu/lsu/n24 [29], \exu/lsu/n22 [29], \exu/lsu/n23 [29]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u819  (\exu/lsu/n24 [30], \exu/lsu/n22 [30], \exu/lsu/n23 [30]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u82  (\exu/data_lsu_cache [50], \exu/lsu/n64 [31], \exu/lsu/n65 [50]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u820  (\exu/lsu/n24 [31], \exu/lsu/n22 [31], \exu/lsu/n23 [31]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u821  (\exu/lsu/n24 [32], \exu/lsu/n22 [32], \exu/lsu/n23 [32]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u822  (\exu/lsu/n24 [33], \exu/lsu/n22 [33], \exu/lsu/n23 [33]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u823  (\exu/lsu/n24 [34], \exu/lsu/n22 [34], \exu/lsu/n23 [34]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u824  (\exu/lsu/n24 [35], \exu/lsu/n22 [35], \exu/lsu/n23 [35]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u825  (\exu/lsu/n24 [36], \exu/lsu/n22 [36], \exu/lsu/n23 [36]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u826  (\exu/lsu/n24 [37], \exu/lsu/n22 [37], \exu/lsu/n23 [37]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u827  (\exu/lsu/n24 [38], \exu/lsu/n22 [38], \exu/lsu/n23 [38]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u828  (\exu/lsu/n24 [39], \exu/lsu/n22 [39], \exu/lsu/n23 [39]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u829  (\exu/lsu/n24 [40], \exu/lsu/n22 [40], \exu/lsu/n23 [40]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u83  (\exu/data_lsu_cache [51], \exu/lsu/n64 [31], \exu/lsu/n65 [51]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u830  (\exu/lsu/n24 [41], \exu/lsu/n22 [41], \exu/lsu/n23 [41]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u831  (\exu/lsu/n24 [42], \exu/lsu/n22 [42], \exu/lsu/n23 [42]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u832  (\exu/lsu/n24 [43], \exu/lsu/n22 [43], \exu/lsu/n23 [43]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u833  (\exu/lsu/n24 [44], \exu/lsu/n22 [44], \exu/lsu/n23 [44]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u834  (\exu/lsu/n24 [45], \exu/lsu/n22 [45], \exu/lsu/n23 [45]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u835  (\exu/lsu/n24 [46], \exu/lsu/n22 [46], \exu/lsu/n23 [46]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u836  (\exu/lsu/n24 [47], \exu/lsu/n22 [47], \exu/lsu/n23 [47]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u837  (\exu/lsu/data_lsu_uncache_shift [48], \exu/lsu/n22 [48], \exu/lsu/n23 [48]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u838  (\exu/lsu/data_lsu_uncache_shift [49], \exu/lsu/n22 [49], \exu/lsu/n23 [49]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u839  (\exu/lsu/data_lsu_uncache_shift [50], \exu/lsu/n22 [50], \exu/lsu/n23 [50]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u84  (\exu/data_lsu_cache [52], \exu/lsu/n64 [31], \exu/lsu/n65 [52]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u840  (\exu/lsu/data_lsu_uncache_shift [51], \exu/lsu/n22 [51], \exu/lsu/n23 [51]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u841  (\exu/lsu/data_lsu_uncache_shift [52], \exu/lsu/n22 [52], \exu/lsu/n23 [52]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u842  (\exu/lsu/data_lsu_uncache_shift [53], \exu/lsu/n22 [53], \exu/lsu/n23 [53]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u843  (\exu/lsu/data_lsu_uncache_shift [54], \exu/lsu/n22 [54], \exu/lsu/n23 [54]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u844  (\exu/lsu/data_lsu_uncache_shift [55], \exu/lsu/n22 [55], \exu/lsu/n23 [55]);  // ../../RTL/CPU/EX/LSU/lsu.v(43)
  or \exu/lsu/u85  (\exu/data_lsu_cache [53], \exu/lsu/n64 [31], \exu/lsu/n65 [53]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u86  (\exu/data_lsu_cache [54], \exu/lsu/n64 [31], \exu/lsu/n65 [54]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u87  (\exu/data_lsu_cache [55], \exu/lsu/n64 [31], \exu/lsu/n65 [55]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u88  (\exu/data_lsu_cache [56], \exu/lsu/n64 [31], \exu/lsu/n65 [56]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u89  (\exu/data_lsu_cache [57], \exu/lsu/n64 [31], \exu/lsu/n65 [57]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u90  (\exu/data_lsu_cache [58], \exu/lsu/n64 [31], \exu/lsu/n65 [58]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u91  (\exu/data_lsu_cache [59], \exu/lsu/n64 [31], \exu/lsu/n65 [59]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u92  (\exu/data_lsu_cache [60], \exu/lsu/n64 [31], \exu/lsu/n65 [60]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u93  (\exu/data_lsu_cache [61], \exu/lsu/n64 [31], \exu/lsu/n65 [61]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u94  (\exu/data_lsu_cache [62], \exu/lsu/n64 [31], \exu/lsu/n65 [62]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u95  (\exu/data_lsu_cache [63], \exu/lsu/n64 [31], \exu/lsu/n65 [63]);  // ../../RTL/CPU/EX/LSU/lsu.v(70)
  or \exu/lsu/u96  (\exu/lsu/n64 [1], \exu/lsu/n62 [1], \exu/lsu/n63 [1]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u97  (\exu/lsu/n64 [2], \exu/lsu/n62 [2], \exu/lsu/n63 [2]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u98  (\exu/lsu/n64 [3], \exu/lsu/n62 [3], \exu/lsu/n63 [3]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  or \exu/lsu/u99  (\exu/lsu/n64 [4], \exu/lsu/n62 [4], \exu/lsu/n63 [4]);  // ../../RTL/CPU/EX/LSU/lsu.v(69)
  reg_sr_as_w1 \exu/m_ret_reg  (
    .clk(clk),
    .d(ex_m_ret),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_m_ret));  // ../../RTL/CPU/EX/exu.v(448)
  binary_mux_s1_w1 \exu/mux0_b2  (
    .i0(\exu/main_state [2]),
    .i1(1'b1),
    .sel(\exu/n21 ),
    .o(\exu/n22 [2]));  // ../../RTL/CPU/EX/exu.v(240)
  binary_mux_s1_w1 \exu/mux10_b0  (
    .i0(\exu/n29 [2]),
    .i1(1'b0),
    .sel(ex_more_exception),
    .o(\exu/n36 [0]));  // ../../RTL/CPU/EX/exu.v(265)
  binary_mux_s1_w1 \exu/mux11_b0  (
    .i0(\exu/main_state [0]),
    .i1(\exu/n36 [0]),
    .sel(\exu/c_amo_mem1 ),
    .o(\exu/n37 [0]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux11_b1  (
    .i0(\exu/main_state [1]),
    .i1(\exu/n36 [0]),
    .sel(\exu/c_amo_mem1 ),
    .o(\exu/n37 [1]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux11_b3  (
    .i0(\exu/main_state [3]),
    .i1(\exu/n36 [0]),
    .sel(\exu/c_amo_mem1 ),
    .o(\exu/n37 [3]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux12_b0  (
    .i0(\exu/n37 [0]),
    .i1(1'b0),
    .sel(\exu/c_amo_mem01 ),
    .o(\exu/n38 [0]));  // ../../RTL/CPU/EX/exu.v(266)
  and \exu/mux12_b2_sel_is_0  (\exu/mux12_b2_sel_is_0_o , \exu/c_amo_mem01_neg , \exu/c_amo_mem1_neg );
  binary_mux_s1_w1 \exu/mux13_b0  (
    .i0(\exu/n38 [0]),
    .i1(1'b1),
    .sel(\exu/n35 ),
    .o(\exu/n39 [0]));  // ../../RTL/CPU/EX/exu.v(266)
  AL_MUX \exu/mux13_b1  (
    .i0(1'b1),
    .i1(\exu/n37 [1]),
    .sel(\exu/mux13_b1_sel_is_0_o ),
    .o(\exu/n39 [1]));
  and \exu/mux13_b1_sel_is_0  (\exu/mux13_b1_sel_is_0_o , \exu/n35_neg , \exu/c_amo_mem01_neg );
  AL_MUX \exu/mux13_b2  (
    .i0(1'b0),
    .i1(\exu/main_state [2]),
    .sel(\exu/mux13_b2_sel_is_2_o ),
    .o(\exu/n39 [2]));
  and \exu/mux13_b2_sel_is_2  (\exu/mux13_b2_sel_is_2_o , \exu/n35_neg , \exu/mux12_b2_sel_is_0_o );
  AL_MUX \exu/mux13_b3  (
    .i0(1'b1),
    .i1(\exu/n37 [3]),
    .sel(\exu/mux13_b1_sel_is_0_o ),
    .o(\exu/n39 [3]));
  binary_mux_s1_w1 \exu/mux14_b0  (
    .i0(\exu/n39 [0]),
    .i1(1'b0),
    .sel(\exu/c_fence ),
    .o(\exu/n40 [0]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux14_b1  (
    .i0(\exu/n39 [1]),
    .i1(1'b0),
    .sel(\exu/c_fence ),
    .o(\exu/n40 [1]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux14_b2  (
    .i0(\exu/n39 [2]),
    .i1(\exu/n36 [0]),
    .sel(\exu/c_fence ),
    .o(\exu/n40 [2]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux14_b3  (
    .i0(\exu/n39 [3]),
    .i1(\exu/n36 [0]),
    .sel(\exu/c_fence ),
    .o(\exu/n40 [3]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux15_b0  (
    .i0(\exu/n40 [0]),
    .i1(\exu/n33 [0]),
    .sel(\exu/c_amo_mem0 ),
    .o(\exu/n41 [0]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux15_b1  (
    .i0(\exu/n40 [1]),
    .i1(\exu/n33 [1]),
    .sel(\exu/c_amo_mem0 ),
    .o(\exu/n41 [1]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux15_b3  (
    .i0(\exu/n40 [3]),
    .i1(\exu/n33 [3]),
    .sel(\exu/c_amo_mem0 ),
    .o(\exu/n41 [3]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux16_b0  (
    .i0(\exu/n41 [0]),
    .i1(\exu/n31 ),
    .sel(\exu/c_shift ),
    .o(\exu/n42 [0]));  // ../../RTL/CPU/EX/exu.v(266)
  AL_MUX \exu/mux16_b2  (
    .i0(1'b0),
    .i1(\exu/n40 [2]),
    .sel(\exu/mux16_b2_sel_is_0_o ),
    .o(\exu/n42 [2]));
  and \exu/mux16_b2_sel_is_0  (\exu/mux16_b2_sel_is_0_o , \exu/c_shift_neg , \exu/c_amo_mem0_neg );
  binary_mux_s1_w1 \exu/mux17_b0  (
    .i0(\exu/n42 [0]),
    .i1(1'b0),
    .sel(\exu/c_store ),
    .o(\exu/n43 [0]));  // ../../RTL/CPU/EX/exu.v(266)
  AL_MUX \exu/mux17_b1  (
    .i0(1'b0),
    .i1(\exu/n41 [1]),
    .sel(\exu/mux17_b1_sel_is_0_o ),
    .o(\exu/n43 [1]));
  and \exu/mux17_b1_sel_is_0  (\exu/mux17_b1_sel_is_0_o , \exu/c_store_neg , \exu/c_shift_neg );
  binary_mux_s1_w1 \exu/mux17_b2  (
    .i0(\exu/n42 [2]),
    .i1(\exu/n36 [0]),
    .sel(\exu/c_store ),
    .o(\exu/n43 [2]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux18_b0  (
    .i0(\exu/n43 [0]),
    .i1(\exu/n27 [0]),
    .sel(\exu/c_load ),
    .o(\exu/n44 [0]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux18_b1  (
    .i0(\exu/n43 [1]),
    .i1(\exu/n27 [1]),
    .sel(\exu/c_load ),
    .o(\exu/n44 [1]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux18_b2  (
    .i0(\exu/n43 [2]),
    .i1(1'b0),
    .sel(\exu/c_load ),
    .o(\exu/n44 [2]));  // ../../RTL/CPU/EX/exu.v(266)
  AL_MUX \exu/mux18_b3  (
    .i0(1'b0),
    .i1(\exu/n41 [3]),
    .sel(\exu/mux18_b3_sel_is_2_o ),
    .o(\exu/n44 [3]));
  and \exu/mux18_b3_sel_is_2  (\exu/mux18_b3_sel_is_2_o , \exu/c_load_neg , \exu/mux17_b1_sel_is_0_o );
  binary_mux_s1_w1 \exu/mux19_b0  (
    .i0(\exu/n44 [0]),
    .i1(\exu/n26 [0]),
    .sel(\exu/n19 ),
    .o(\exu/n45 [0]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux19_b1  (
    .i0(\exu/n44 [1]),
    .i1(\exu/n26 [1]),
    .sel(\exu/n19 ),
    .o(\exu/n45 [1]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux19_b2  (
    .i0(\exu/n44 [2]),
    .i1(\exu/n26 [2]),
    .sel(\exu/n19 ),
    .o(\exu/n45 [2]));  // ../../RTL/CPU/EX/exu.v(266)
  binary_mux_s1_w1 \exu/mux19_b3  (
    .i0(\exu/n44 [3]),
    .i1(\exu/n26 [3]),
    .sel(\exu/n19 ),
    .o(\exu/n45 [3]));  // ../../RTL/CPU/EX/exu.v(266)
  AL_MUX \exu/mux1_b0  (
    .i0(1'b0),
    .i1(\exu/main_state [0]),
    .sel(\exu/mux1_b0_sel_is_0_o ),
    .o(\exu/n23 [0]));
  and \exu/mux1_b0_sel_is_0  (\exu/mux1_b0_sel_is_0_o , amo_neg, \exu/n21_neg );
  AL_MUX \exu/mux1_b3  (
    .i0(1'b1),
    .i1(\exu/main_state [3]),
    .sel(\exu/mux1_b0_sel_is_0_o ),
    .o(\exu/n23 [3]));
  binary_mux_s1_w1 \exu/mux22_b0  (
    .i0(\exu/shift_count [0]),
    .i1(\exu/n50 [0]),
    .sel(\exu/c_shift ),
    .o(\exu/n51 [0]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux22_b1  (
    .i0(\exu/shift_count [1]),
    .i1(\exu/n50 [1]),
    .sel(\exu/c_shift ),
    .o(\exu/n51 [1]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux22_b2  (
    .i0(\exu/shift_count [2]),
    .i1(\exu/n50 [2]),
    .sel(\exu/c_shift ),
    .o(\exu/n51 [2]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux22_b3  (
    .i0(\exu/shift_count [3]),
    .i1(\exu/n50 [3]),
    .sel(\exu/c_shift ),
    .o(\exu/n51 [3]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux22_b4  (
    .i0(\exu/shift_count [4]),
    .i1(\exu/n50 [4]),
    .sel(\exu/c_shift ),
    .o(\exu/n51 [4]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux22_b5  (
    .i0(\exu/shift_count [5]),
    .i1(\exu/n50 [5]),
    .sel(\exu/c_shift ),
    .o(\exu/n51 [5]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux22_b6  (
    .i0(\exu/shift_count [6]),
    .i1(\exu/n50 [6]),
    .sel(\exu/c_shift ),
    .o(\exu/n51 [6]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux22_b7  (
    .i0(\exu/shift_count [7]),
    .i1(\exu/n50 [7]),
    .sel(\exu/c_shift ),
    .o(\exu/n51 [7]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux23_b0  (
    .i0(\exu/n51 [0]),
    .i1(op_count[0]),
    .sel(\exu/n49 ),
    .o(\exu/n52 [0]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux23_b1  (
    .i0(\exu/n51 [1]),
    .i1(op_count[1]),
    .sel(\exu/n49 ),
    .o(\exu/n52 [1]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux23_b2  (
    .i0(\exu/n51 [2]),
    .i1(op_count[2]),
    .sel(\exu/n49 ),
    .o(\exu/n52 [2]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux23_b3  (
    .i0(\exu/n51 [3]),
    .i1(op_count[3]),
    .sel(\exu/n49 ),
    .o(\exu/n52 [3]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux23_b4  (
    .i0(\exu/n51 [4]),
    .i1(op_count[4]),
    .sel(\exu/n49 ),
    .o(\exu/n52 [4]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux23_b5  (
    .i0(\exu/n51 [5]),
    .i1(op_count[5]),
    .sel(\exu/n49 ),
    .o(\exu/n52 [5]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux23_b6  (
    .i0(\exu/n51 [6]),
    .i1(op_count[6]),
    .sel(\exu/n49 ),
    .o(\exu/n52 [6]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux23_b7  (
    .i0(\exu/n51 [7]),
    .i1(op_count[7]),
    .sel(\exu/n49 ),
    .o(\exu/n52 [7]));  // ../../RTL/CPU/EX/exu.v(289)
  binary_mux_s1_w1 \exu/mux25_b0  (
    .i0(data_rd[31]),
    .i1(data_rd[32]),
    .sel(ex_size[2]),
    .o(\exu/n54 [0]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b1  (
    .i0(data_rd[32]),
    .i1(data_rd[33]),
    .sel(ex_size[2]),
    .o(\exu/n54 [1]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b10  (
    .i0(data_rd[41]),
    .i1(data_rd[42]),
    .sel(ex_size[2]),
    .o(\exu/n54 [10]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b11  (
    .i0(data_rd[42]),
    .i1(data_rd[43]),
    .sel(ex_size[2]),
    .o(\exu/n54 [11]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b12  (
    .i0(data_rd[43]),
    .i1(data_rd[44]),
    .sel(ex_size[2]),
    .o(\exu/n54 [12]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b13  (
    .i0(data_rd[44]),
    .i1(data_rd[45]),
    .sel(ex_size[2]),
    .o(\exu/n54 [13]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b14  (
    .i0(data_rd[45]),
    .i1(data_rd[46]),
    .sel(ex_size[2]),
    .o(\exu/n54 [14]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b15  (
    .i0(data_rd[46]),
    .i1(data_rd[47]),
    .sel(ex_size[2]),
    .o(\exu/n54 [15]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b16  (
    .i0(data_rd[47]),
    .i1(data_rd[48]),
    .sel(ex_size[2]),
    .o(\exu/n54 [16]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b17  (
    .i0(data_rd[48]),
    .i1(data_rd[49]),
    .sel(ex_size[2]),
    .o(\exu/n54 [17]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b18  (
    .i0(data_rd[49]),
    .i1(data_rd[50]),
    .sel(ex_size[2]),
    .o(\exu/n54 [18]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b19  (
    .i0(data_rd[50]),
    .i1(data_rd[51]),
    .sel(ex_size[2]),
    .o(\exu/n54 [19]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b2  (
    .i0(data_rd[33]),
    .i1(data_rd[34]),
    .sel(ex_size[2]),
    .o(\exu/n54 [2]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b20  (
    .i0(data_rd[51]),
    .i1(data_rd[52]),
    .sel(ex_size[2]),
    .o(\exu/n54 [20]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b21  (
    .i0(data_rd[52]),
    .i1(data_rd[53]),
    .sel(ex_size[2]),
    .o(\exu/n54 [21]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b22  (
    .i0(data_rd[53]),
    .i1(data_rd[54]),
    .sel(ex_size[2]),
    .o(\exu/n54 [22]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b23  (
    .i0(data_rd[54]),
    .i1(data_rd[55]),
    .sel(ex_size[2]),
    .o(\exu/n54 [23]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b24  (
    .i0(data_rd[55]),
    .i1(data_rd[56]),
    .sel(ex_size[2]),
    .o(\exu/n54 [24]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b25  (
    .i0(data_rd[56]),
    .i1(data_rd[57]),
    .sel(ex_size[2]),
    .o(\exu/n54 [25]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b26  (
    .i0(data_rd[57]),
    .i1(data_rd[58]),
    .sel(ex_size[2]),
    .o(\exu/n54 [26]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b27  (
    .i0(data_rd[58]),
    .i1(data_rd[59]),
    .sel(ex_size[2]),
    .o(\exu/n54 [27]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b28  (
    .i0(data_rd[59]),
    .i1(data_rd[60]),
    .sel(ex_size[2]),
    .o(\exu/n54 [28]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b29  (
    .i0(data_rd[60]),
    .i1(data_rd[61]),
    .sel(ex_size[2]),
    .o(\exu/n54 [29]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b3  (
    .i0(data_rd[34]),
    .i1(data_rd[35]),
    .sel(ex_size[2]),
    .o(\exu/n54 [3]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b30  (
    .i0(data_rd[61]),
    .i1(data_rd[62]),
    .sel(ex_size[2]),
    .o(\exu/n54 [30]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b31  (
    .i0(data_rd[62]),
    .i1(data_rd[63]),
    .sel(ex_size[2]),
    .o(\exu/n54 [31]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b4  (
    .i0(data_rd[35]),
    .i1(data_rd[36]),
    .sel(ex_size[2]),
    .o(\exu/n54 [4]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b5  (
    .i0(data_rd[36]),
    .i1(data_rd[37]),
    .sel(ex_size[2]),
    .o(\exu/n54 [5]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b6  (
    .i0(data_rd[37]),
    .i1(data_rd[38]),
    .sel(ex_size[2]),
    .o(\exu/n54 [6]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b7  (
    .i0(data_rd[38]),
    .i1(data_rd[39]),
    .sel(ex_size[2]),
    .o(\exu/n54 [7]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b8  (
    .i0(data_rd[39]),
    .i1(data_rd[40]),
    .sel(ex_size[2]),
    .o(\exu/n54 [8]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux25_b9  (
    .i0(data_rd[40]),
    .i1(data_rd[41]),
    .sel(ex_size[2]),
    .o(\exu/n54 [9]));  // ../../RTL/CPU/EX/exu.v(303)
  binary_mux_s1_w1 \exu/mux26_b0  (
    .i0(data_rd[32]),
    .i1(1'b0),
    .sel(ex_size[2]),
    .o(\exu/n55 [0]));  // ../../RTL/CPU/EX/exu.v(310)
  binary_mux_s1_w1 \exu/mux26_b33  (
    .i0(data_rd[32]),
    .i1(data_rd[31]),
    .sel(ex_size[2]),
    .o(\exu/n55 [33]));  // ../../RTL/CPU/EX/exu.v(310)
  binary_mux_s1_w1 \exu/mux27_b0  (
    .i0(data_rd[0]),
    .i1(data_rd[1]),
    .sel(shift_r),
    .o(\exu/n57 [0]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b1  (
    .i0(data_rd[1]),
    .i1(data_rd[2]),
    .sel(shift_r),
    .o(\exu/n57 [1]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b10  (
    .i0(data_rd[10]),
    .i1(data_rd[11]),
    .sel(shift_r),
    .o(\exu/n57 [10]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b11  (
    .i0(data_rd[11]),
    .i1(data_rd[12]),
    .sel(shift_r),
    .o(\exu/n57 [11]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b12  (
    .i0(data_rd[12]),
    .i1(data_rd[13]),
    .sel(shift_r),
    .o(\exu/n57 [12]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b13  (
    .i0(data_rd[13]),
    .i1(data_rd[14]),
    .sel(shift_r),
    .o(\exu/n57 [13]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b14  (
    .i0(data_rd[14]),
    .i1(data_rd[15]),
    .sel(shift_r),
    .o(\exu/n57 [14]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b15  (
    .i0(data_rd[15]),
    .i1(data_rd[16]),
    .sel(shift_r),
    .o(\exu/n57 [15]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b16  (
    .i0(data_rd[16]),
    .i1(data_rd[17]),
    .sel(shift_r),
    .o(\exu/n57 [16]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b17  (
    .i0(data_rd[17]),
    .i1(data_rd[18]),
    .sel(shift_r),
    .o(\exu/n57 [17]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b18  (
    .i0(data_rd[18]),
    .i1(data_rd[19]),
    .sel(shift_r),
    .o(\exu/n57 [18]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b19  (
    .i0(data_rd[19]),
    .i1(data_rd[20]),
    .sel(shift_r),
    .o(\exu/n57 [19]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b2  (
    .i0(data_rd[2]),
    .i1(data_rd[3]),
    .sel(shift_r),
    .o(\exu/n57 [2]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b20  (
    .i0(data_rd[20]),
    .i1(data_rd[21]),
    .sel(shift_r),
    .o(\exu/n57 [20]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b21  (
    .i0(data_rd[21]),
    .i1(data_rd[22]),
    .sel(shift_r),
    .o(\exu/n57 [21]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b22  (
    .i0(data_rd[22]),
    .i1(data_rd[23]),
    .sel(shift_r),
    .o(\exu/n57 [22]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b23  (
    .i0(data_rd[23]),
    .i1(data_rd[24]),
    .sel(shift_r),
    .o(\exu/n57 [23]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b24  (
    .i0(data_rd[24]),
    .i1(data_rd[25]),
    .sel(shift_r),
    .o(\exu/n57 [24]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b25  (
    .i0(data_rd[25]),
    .i1(data_rd[26]),
    .sel(shift_r),
    .o(\exu/n57 [25]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b26  (
    .i0(data_rd[26]),
    .i1(data_rd[27]),
    .sel(shift_r),
    .o(\exu/n57 [26]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b27  (
    .i0(data_rd[27]),
    .i1(data_rd[28]),
    .sel(shift_r),
    .o(\exu/n57 [27]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b28  (
    .i0(data_rd[28]),
    .i1(data_rd[29]),
    .sel(shift_r),
    .o(\exu/n57 [28]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b29  (
    .i0(data_rd[29]),
    .i1(data_rd[30]),
    .sel(shift_r),
    .o(\exu/n57 [29]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b3  (
    .i0(data_rd[3]),
    .i1(data_rd[4]),
    .sel(shift_r),
    .o(\exu/n57 [3]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b30  (
    .i0(data_rd[30]),
    .i1(data_rd[31]),
    .sel(shift_r),
    .o(\exu/n57 [30]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b31  (
    .i0(data_rd[31]),
    .i1(\exu/n56 [0]),
    .sel(shift_r),
    .o(\exu/n57 [31]));  // ../../RTL/CPU/EX/exu.v(312)
  AL_MUX \exu/mux27_b32  (
    .i0(data_rd[32]),
    .i1(data_rd[33]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [32]));
  and \exu/mux27_b32_sel_is_1  (\exu/mux27_b32_sel_is_1_o , shift_r, \ex_size[2]_neg );
  AL_MUX \exu/mux27_b33  (
    .i0(data_rd[33]),
    .i1(data_rd[34]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [33]));
  AL_MUX \exu/mux27_b34  (
    .i0(data_rd[34]),
    .i1(data_rd[35]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [34]));
  AL_MUX \exu/mux27_b35  (
    .i0(data_rd[35]),
    .i1(data_rd[36]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [35]));
  AL_MUX \exu/mux27_b36  (
    .i0(data_rd[36]),
    .i1(data_rd[37]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [36]));
  AL_MUX \exu/mux27_b37  (
    .i0(data_rd[37]),
    .i1(data_rd[38]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [37]));
  AL_MUX \exu/mux27_b38  (
    .i0(data_rd[38]),
    .i1(data_rd[39]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [38]));
  AL_MUX \exu/mux27_b39  (
    .i0(data_rd[39]),
    .i1(data_rd[40]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [39]));
  binary_mux_s1_w1 \exu/mux27_b4  (
    .i0(data_rd[4]),
    .i1(data_rd[5]),
    .sel(shift_r),
    .o(\exu/n57 [4]));  // ../../RTL/CPU/EX/exu.v(312)
  AL_MUX \exu/mux27_b40  (
    .i0(data_rd[40]),
    .i1(data_rd[41]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [40]));
  AL_MUX \exu/mux27_b41  (
    .i0(data_rd[41]),
    .i1(data_rd[42]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [41]));
  AL_MUX \exu/mux27_b42  (
    .i0(data_rd[42]),
    .i1(data_rd[43]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [42]));
  AL_MUX \exu/mux27_b43  (
    .i0(data_rd[43]),
    .i1(data_rd[44]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [43]));
  AL_MUX \exu/mux27_b44  (
    .i0(data_rd[44]),
    .i1(data_rd[45]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [44]));
  AL_MUX \exu/mux27_b45  (
    .i0(data_rd[45]),
    .i1(data_rd[46]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [45]));
  AL_MUX \exu/mux27_b46  (
    .i0(data_rd[46]),
    .i1(data_rd[47]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [46]));
  AL_MUX \exu/mux27_b47  (
    .i0(data_rd[47]),
    .i1(data_rd[48]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [47]));
  AL_MUX \exu/mux27_b48  (
    .i0(data_rd[48]),
    .i1(data_rd[49]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [48]));
  AL_MUX \exu/mux27_b49  (
    .i0(data_rd[49]),
    .i1(data_rd[50]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [49]));
  binary_mux_s1_w1 \exu/mux27_b5  (
    .i0(data_rd[5]),
    .i1(data_rd[6]),
    .sel(shift_r),
    .o(\exu/n57 [5]));  // ../../RTL/CPU/EX/exu.v(312)
  AL_MUX \exu/mux27_b50  (
    .i0(data_rd[50]),
    .i1(data_rd[51]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [50]));
  AL_MUX \exu/mux27_b51  (
    .i0(data_rd[51]),
    .i1(data_rd[52]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [51]));
  AL_MUX \exu/mux27_b52  (
    .i0(data_rd[52]),
    .i1(data_rd[53]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [52]));
  AL_MUX \exu/mux27_b53  (
    .i0(data_rd[53]),
    .i1(data_rd[54]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [53]));
  AL_MUX \exu/mux27_b54  (
    .i0(data_rd[54]),
    .i1(data_rd[55]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [54]));
  AL_MUX \exu/mux27_b55  (
    .i0(data_rd[55]),
    .i1(data_rd[56]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [55]));
  AL_MUX \exu/mux27_b56  (
    .i0(data_rd[56]),
    .i1(data_rd[57]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [56]));
  AL_MUX \exu/mux27_b57  (
    .i0(data_rd[57]),
    .i1(data_rd[58]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [57]));
  AL_MUX \exu/mux27_b58  (
    .i0(data_rd[58]),
    .i1(data_rd[59]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [58]));
  AL_MUX \exu/mux27_b59  (
    .i0(data_rd[59]),
    .i1(data_rd[60]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [59]));
  binary_mux_s1_w1 \exu/mux27_b6  (
    .i0(data_rd[6]),
    .i1(data_rd[7]),
    .sel(shift_r),
    .o(\exu/n57 [6]));  // ../../RTL/CPU/EX/exu.v(312)
  AL_MUX \exu/mux27_b60  (
    .i0(data_rd[60]),
    .i1(data_rd[61]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [60]));
  AL_MUX \exu/mux27_b61  (
    .i0(data_rd[61]),
    .i1(data_rd[62]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [61]));
  AL_MUX \exu/mux27_b62  (
    .i0(data_rd[62]),
    .i1(data_rd[63]),
    .sel(\exu/mux27_b32_sel_is_1_o ),
    .o(\exu/n57 [62]));
  AL_MUX \exu/mux27_b63  (
    .i0(data_rd[63]),
    .i1(1'b0),
    .sel(\exu/mux27_b63_sel_is_3_o ),
    .o(\exu/n57 [63]));
  and \exu/mux27_b63_sel_is_3  (\exu/mux27_b63_sel_is_3_o , shift_r, \exu/mux48_b32_sel_is_1_o );
  binary_mux_s1_w1 \exu/mux27_b7  (
    .i0(data_rd[7]),
    .i1(data_rd[8]),
    .sel(shift_r),
    .o(\exu/n57 [7]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b8  (
    .i0(data_rd[8]),
    .i1(data_rd[9]),
    .sel(shift_r),
    .o(\exu/n57 [8]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux27_b9  (
    .i0(data_rd[9]),
    .i1(data_rd[10]),
    .sel(shift_r),
    .o(\exu/n57 [9]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b0  (
    .i0(\exu/n57 [0]),
    .i1(1'b0),
    .sel(shift_l),
    .o(\exu/n58 [0]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b1  (
    .i0(\exu/n57 [1]),
    .i1(data_rd[0]),
    .sel(shift_l),
    .o(\exu/n58 [1]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b10  (
    .i0(\exu/n57 [10]),
    .i1(data_rd[9]),
    .sel(shift_l),
    .o(\exu/n58 [10]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b11  (
    .i0(\exu/n57 [11]),
    .i1(data_rd[10]),
    .sel(shift_l),
    .o(\exu/n58 [11]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b12  (
    .i0(\exu/n57 [12]),
    .i1(data_rd[11]),
    .sel(shift_l),
    .o(\exu/n58 [12]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b13  (
    .i0(\exu/n57 [13]),
    .i1(data_rd[12]),
    .sel(shift_l),
    .o(\exu/n58 [13]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b14  (
    .i0(\exu/n57 [14]),
    .i1(data_rd[13]),
    .sel(shift_l),
    .o(\exu/n58 [14]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b15  (
    .i0(\exu/n57 [15]),
    .i1(data_rd[14]),
    .sel(shift_l),
    .o(\exu/n58 [15]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b16  (
    .i0(\exu/n57 [16]),
    .i1(data_rd[15]),
    .sel(shift_l),
    .o(\exu/n58 [16]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b17  (
    .i0(\exu/n57 [17]),
    .i1(data_rd[16]),
    .sel(shift_l),
    .o(\exu/n58 [17]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b18  (
    .i0(\exu/n57 [18]),
    .i1(data_rd[17]),
    .sel(shift_l),
    .o(\exu/n58 [18]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b19  (
    .i0(\exu/n57 [19]),
    .i1(data_rd[18]),
    .sel(shift_l),
    .o(\exu/n58 [19]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b2  (
    .i0(\exu/n57 [2]),
    .i1(data_rd[1]),
    .sel(shift_l),
    .o(\exu/n58 [2]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b20  (
    .i0(\exu/n57 [20]),
    .i1(data_rd[19]),
    .sel(shift_l),
    .o(\exu/n58 [20]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b21  (
    .i0(\exu/n57 [21]),
    .i1(data_rd[20]),
    .sel(shift_l),
    .o(\exu/n58 [21]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b22  (
    .i0(\exu/n57 [22]),
    .i1(data_rd[21]),
    .sel(shift_l),
    .o(\exu/n58 [22]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b23  (
    .i0(\exu/n57 [23]),
    .i1(data_rd[22]),
    .sel(shift_l),
    .o(\exu/n58 [23]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b24  (
    .i0(\exu/n57 [24]),
    .i1(data_rd[23]),
    .sel(shift_l),
    .o(\exu/n58 [24]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b25  (
    .i0(\exu/n57 [25]),
    .i1(data_rd[24]),
    .sel(shift_l),
    .o(\exu/n58 [25]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b26  (
    .i0(\exu/n57 [26]),
    .i1(data_rd[25]),
    .sel(shift_l),
    .o(\exu/n58 [26]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b27  (
    .i0(\exu/n57 [27]),
    .i1(data_rd[26]),
    .sel(shift_l),
    .o(\exu/n58 [27]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b28  (
    .i0(\exu/n57 [28]),
    .i1(data_rd[27]),
    .sel(shift_l),
    .o(\exu/n58 [28]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b29  (
    .i0(\exu/n57 [29]),
    .i1(data_rd[28]),
    .sel(shift_l),
    .o(\exu/n58 [29]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b3  (
    .i0(\exu/n57 [3]),
    .i1(data_rd[2]),
    .sel(shift_l),
    .o(\exu/n58 [3]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b30  (
    .i0(\exu/n57 [30]),
    .i1(data_rd[29]),
    .sel(shift_l),
    .o(\exu/n58 [30]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b31  (
    .i0(\exu/n57 [31]),
    .i1(data_rd[30]),
    .sel(shift_l),
    .o(\exu/n58 [31]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b32  (
    .i0(\exu/n57 [32]),
    .i1(\exu/n54 [0]),
    .sel(shift_l),
    .o(\exu/n58 [32]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b33  (
    .i0(\exu/n57 [33]),
    .i1(\exu/n54 [1]),
    .sel(shift_l),
    .o(\exu/n58 [33]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b34  (
    .i0(\exu/n57 [34]),
    .i1(\exu/n54 [2]),
    .sel(shift_l),
    .o(\exu/n58 [34]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b35  (
    .i0(\exu/n57 [35]),
    .i1(\exu/n54 [3]),
    .sel(shift_l),
    .o(\exu/n58 [35]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b36  (
    .i0(\exu/n57 [36]),
    .i1(\exu/n54 [4]),
    .sel(shift_l),
    .o(\exu/n58 [36]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b37  (
    .i0(\exu/n57 [37]),
    .i1(\exu/n54 [5]),
    .sel(shift_l),
    .o(\exu/n58 [37]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b38  (
    .i0(\exu/n57 [38]),
    .i1(\exu/n54 [6]),
    .sel(shift_l),
    .o(\exu/n58 [38]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b39  (
    .i0(\exu/n57 [39]),
    .i1(\exu/n54 [7]),
    .sel(shift_l),
    .o(\exu/n58 [39]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b4  (
    .i0(\exu/n57 [4]),
    .i1(data_rd[3]),
    .sel(shift_l),
    .o(\exu/n58 [4]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b40  (
    .i0(\exu/n57 [40]),
    .i1(\exu/n54 [8]),
    .sel(shift_l),
    .o(\exu/n58 [40]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b41  (
    .i0(\exu/n57 [41]),
    .i1(\exu/n54 [9]),
    .sel(shift_l),
    .o(\exu/n58 [41]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b42  (
    .i0(\exu/n57 [42]),
    .i1(\exu/n54 [10]),
    .sel(shift_l),
    .o(\exu/n58 [42]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b43  (
    .i0(\exu/n57 [43]),
    .i1(\exu/n54 [11]),
    .sel(shift_l),
    .o(\exu/n58 [43]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b44  (
    .i0(\exu/n57 [44]),
    .i1(\exu/n54 [12]),
    .sel(shift_l),
    .o(\exu/n58 [44]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b45  (
    .i0(\exu/n57 [45]),
    .i1(\exu/n54 [13]),
    .sel(shift_l),
    .o(\exu/n58 [45]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b46  (
    .i0(\exu/n57 [46]),
    .i1(\exu/n54 [14]),
    .sel(shift_l),
    .o(\exu/n58 [46]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b47  (
    .i0(\exu/n57 [47]),
    .i1(\exu/n54 [15]),
    .sel(shift_l),
    .o(\exu/n58 [47]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b48  (
    .i0(\exu/n57 [48]),
    .i1(\exu/n54 [16]),
    .sel(shift_l),
    .o(\exu/n58 [48]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b49  (
    .i0(\exu/n57 [49]),
    .i1(\exu/n54 [17]),
    .sel(shift_l),
    .o(\exu/n58 [49]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b5  (
    .i0(\exu/n57 [5]),
    .i1(data_rd[4]),
    .sel(shift_l),
    .o(\exu/n58 [5]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b50  (
    .i0(\exu/n57 [50]),
    .i1(\exu/n54 [18]),
    .sel(shift_l),
    .o(\exu/n58 [50]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b51  (
    .i0(\exu/n57 [51]),
    .i1(\exu/n54 [19]),
    .sel(shift_l),
    .o(\exu/n58 [51]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b52  (
    .i0(\exu/n57 [52]),
    .i1(\exu/n54 [20]),
    .sel(shift_l),
    .o(\exu/n58 [52]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b53  (
    .i0(\exu/n57 [53]),
    .i1(\exu/n54 [21]),
    .sel(shift_l),
    .o(\exu/n58 [53]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b54  (
    .i0(\exu/n57 [54]),
    .i1(\exu/n54 [22]),
    .sel(shift_l),
    .o(\exu/n58 [54]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b55  (
    .i0(\exu/n57 [55]),
    .i1(\exu/n54 [23]),
    .sel(shift_l),
    .o(\exu/n58 [55]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b56  (
    .i0(\exu/n57 [56]),
    .i1(\exu/n54 [24]),
    .sel(shift_l),
    .o(\exu/n58 [56]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b57  (
    .i0(\exu/n57 [57]),
    .i1(\exu/n54 [25]),
    .sel(shift_l),
    .o(\exu/n58 [57]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b58  (
    .i0(\exu/n57 [58]),
    .i1(\exu/n54 [26]),
    .sel(shift_l),
    .o(\exu/n58 [58]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b59  (
    .i0(\exu/n57 [59]),
    .i1(\exu/n54 [27]),
    .sel(shift_l),
    .o(\exu/n58 [59]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b6  (
    .i0(\exu/n57 [6]),
    .i1(data_rd[5]),
    .sel(shift_l),
    .o(\exu/n58 [6]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b60  (
    .i0(\exu/n57 [60]),
    .i1(\exu/n54 [28]),
    .sel(shift_l),
    .o(\exu/n58 [60]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b61  (
    .i0(\exu/n57 [61]),
    .i1(\exu/n54 [29]),
    .sel(shift_l),
    .o(\exu/n58 [61]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b62  (
    .i0(\exu/n57 [62]),
    .i1(\exu/n54 [30]),
    .sel(shift_l),
    .o(\exu/n58 [62]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b63  (
    .i0(\exu/n57 [63]),
    .i1(\exu/n54 [31]),
    .sel(shift_l),
    .o(\exu/n58 [63]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b7  (
    .i0(\exu/n57 [7]),
    .i1(data_rd[6]),
    .sel(shift_l),
    .o(\exu/n58 [7]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b8  (
    .i0(\exu/n57 [8]),
    .i1(data_rd[7]),
    .sel(shift_l),
    .o(\exu/n58 [8]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux28_b9  (
    .i0(\exu/n57 [9]),
    .i1(data_rd[8]),
    .sel(shift_l),
    .o(\exu/n58 [9]));  // ../../RTL/CPU/EX/exu.v(312)
  binary_mux_s1_w1 \exu/mux29_b0  (
    .i0(data_rd[0]),
    .i1(\exu/data_lsu_cache [0]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [0]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b1  (
    .i0(data_rd[1]),
    .i1(\exu/data_lsu_cache [1]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [1]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b10  (
    .i0(data_rd[10]),
    .i1(\exu/data_lsu_cache [10]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [10]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b11  (
    .i0(data_rd[11]),
    .i1(\exu/data_lsu_cache [11]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [11]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b12  (
    .i0(data_rd[12]),
    .i1(\exu/data_lsu_cache [12]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [12]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b13  (
    .i0(data_rd[13]),
    .i1(\exu/data_lsu_cache [13]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [13]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b14  (
    .i0(data_rd[14]),
    .i1(\exu/data_lsu_cache [14]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [14]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b15  (
    .i0(data_rd[15]),
    .i1(\exu/data_lsu_cache [15]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [15]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b16  (
    .i0(data_rd[16]),
    .i1(\exu/data_lsu_cache [16]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [16]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b17  (
    .i0(data_rd[17]),
    .i1(\exu/data_lsu_cache [17]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [17]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b18  (
    .i0(data_rd[18]),
    .i1(\exu/data_lsu_cache [18]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [18]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b19  (
    .i0(data_rd[19]),
    .i1(\exu/data_lsu_cache [19]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [19]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b2  (
    .i0(data_rd[2]),
    .i1(\exu/data_lsu_cache [2]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [2]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b20  (
    .i0(data_rd[20]),
    .i1(\exu/data_lsu_cache [20]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [20]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b21  (
    .i0(data_rd[21]),
    .i1(\exu/data_lsu_cache [21]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [21]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b22  (
    .i0(data_rd[22]),
    .i1(\exu/data_lsu_cache [22]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [22]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b23  (
    .i0(data_rd[23]),
    .i1(\exu/data_lsu_cache [23]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [23]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b24  (
    .i0(data_rd[24]),
    .i1(\exu/data_lsu_cache [24]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [24]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b25  (
    .i0(data_rd[25]),
    .i1(\exu/data_lsu_cache [25]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [25]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b26  (
    .i0(data_rd[26]),
    .i1(\exu/data_lsu_cache [26]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [26]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b27  (
    .i0(data_rd[27]),
    .i1(\exu/data_lsu_cache [27]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [27]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b28  (
    .i0(data_rd[28]),
    .i1(\exu/data_lsu_cache [28]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [28]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b29  (
    .i0(data_rd[29]),
    .i1(\exu/data_lsu_cache [29]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [29]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b3  (
    .i0(data_rd[3]),
    .i1(\exu/data_lsu_cache [3]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [3]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b30  (
    .i0(data_rd[30]),
    .i1(\exu/data_lsu_cache [30]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [30]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b31  (
    .i0(data_rd[31]),
    .i1(\exu/data_lsu_cache [31]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [31]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b32  (
    .i0(data_rd[32]),
    .i1(\exu/data_lsu_cache [32]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [32]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b33  (
    .i0(data_rd[33]),
    .i1(\exu/data_lsu_cache [33]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [33]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b34  (
    .i0(data_rd[34]),
    .i1(\exu/data_lsu_cache [34]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [34]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b35  (
    .i0(data_rd[35]),
    .i1(\exu/data_lsu_cache [35]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [35]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b36  (
    .i0(data_rd[36]),
    .i1(\exu/data_lsu_cache [36]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [36]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b37  (
    .i0(data_rd[37]),
    .i1(\exu/data_lsu_cache [37]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [37]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b38  (
    .i0(data_rd[38]),
    .i1(\exu/data_lsu_cache [38]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [38]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b39  (
    .i0(data_rd[39]),
    .i1(\exu/data_lsu_cache [39]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [39]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b4  (
    .i0(data_rd[4]),
    .i1(\exu/data_lsu_cache [4]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [4]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b40  (
    .i0(data_rd[40]),
    .i1(\exu/data_lsu_cache [40]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [40]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b41  (
    .i0(data_rd[41]),
    .i1(\exu/data_lsu_cache [41]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [41]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b42  (
    .i0(data_rd[42]),
    .i1(\exu/data_lsu_cache [42]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [42]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b43  (
    .i0(data_rd[43]),
    .i1(\exu/data_lsu_cache [43]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [43]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b44  (
    .i0(data_rd[44]),
    .i1(\exu/data_lsu_cache [44]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [44]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b45  (
    .i0(data_rd[45]),
    .i1(\exu/data_lsu_cache [45]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [45]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b46  (
    .i0(data_rd[46]),
    .i1(\exu/data_lsu_cache [46]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [46]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b47  (
    .i0(data_rd[47]),
    .i1(\exu/data_lsu_cache [47]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [47]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b48  (
    .i0(data_rd[48]),
    .i1(\exu/data_lsu_cache [48]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [48]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b49  (
    .i0(data_rd[49]),
    .i1(\exu/data_lsu_cache [49]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [49]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b5  (
    .i0(data_rd[5]),
    .i1(\exu/data_lsu_cache [5]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [5]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b50  (
    .i0(data_rd[50]),
    .i1(\exu/data_lsu_cache [50]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [50]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b51  (
    .i0(data_rd[51]),
    .i1(\exu/data_lsu_cache [51]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [51]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b52  (
    .i0(data_rd[52]),
    .i1(\exu/data_lsu_cache [52]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [52]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b53  (
    .i0(data_rd[53]),
    .i1(\exu/data_lsu_cache [53]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [53]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b54  (
    .i0(data_rd[54]),
    .i1(\exu/data_lsu_cache [54]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [54]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b55  (
    .i0(data_rd[55]),
    .i1(\exu/data_lsu_cache [55]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [55]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b56  (
    .i0(data_rd[56]),
    .i1(\exu/data_lsu_cache [56]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [56]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b57  (
    .i0(data_rd[57]),
    .i1(\exu/data_lsu_cache [57]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [57]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b58  (
    .i0(data_rd[58]),
    .i1(\exu/data_lsu_cache [58]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [58]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b59  (
    .i0(data_rd[59]),
    .i1(\exu/data_lsu_cache [59]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [59]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b6  (
    .i0(data_rd[6]),
    .i1(\exu/data_lsu_cache [6]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [6]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b60  (
    .i0(data_rd[60]),
    .i1(\exu/data_lsu_cache [60]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [60]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b61  (
    .i0(data_rd[61]),
    .i1(\exu/data_lsu_cache [61]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [61]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b62  (
    .i0(data_rd[62]),
    .i1(\exu/data_lsu_cache [62]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [62]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b63  (
    .i0(data_rd[63]),
    .i1(\exu/data_lsu_cache [63]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [63]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b7  (
    .i0(data_rd[7]),
    .i1(\exu/data_lsu_cache [7]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [7]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b8  (
    .i0(data_rd[8]),
    .i1(\exu/data_lsu_cache [8]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [8]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux29_b9  (
    .i0(data_rd[9]),
    .i1(\exu/data_lsu_cache [9]),
    .sel(\exu/n60 ),
    .o(\exu/n61 [9]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux2_b0  (
    .i0(\exu/n23 [0]),
    .i1(1'b1),
    .sel(\exu/n20 ),
    .o(\exu/n24 [0]));  // ../../RTL/CPU/EX/exu.v(240)
  and \exu/mux2_b1_sel_is_2  (\exu/mux2_b1_sel_is_2_o , \exu/n20_neg , \exu/mux1_b0_sel_is_0_o );
  AL_MUX \exu/mux2_b2  (
    .i0(1'b0),
    .i1(\exu/n22 [2]),
    .sel(\exu/mux2_b2_sel_is_0_o ),
    .o(\exu/n24 [2]));
  and \exu/mux2_b2_sel_is_0  (\exu/mux2_b2_sel_is_0_o , \exu/n20_neg , amo_neg);
  binary_mux_s1_w1 \exu/mux30_b0  (
    .i0(\exu/n61 [0]),
    .i1(\exu/data_lsu_uncache [0]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [0]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b1  (
    .i0(\exu/n61 [1]),
    .i1(\exu/data_lsu_uncache [1]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [1]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b10  (
    .i0(\exu/n61 [10]),
    .i1(\exu/data_lsu_uncache [10]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [10]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b11  (
    .i0(\exu/n61 [11]),
    .i1(\exu/data_lsu_uncache [11]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [11]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b12  (
    .i0(\exu/n61 [12]),
    .i1(\exu/data_lsu_uncache [12]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [12]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b13  (
    .i0(\exu/n61 [13]),
    .i1(\exu/data_lsu_uncache [13]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [13]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b14  (
    .i0(\exu/n61 [14]),
    .i1(\exu/data_lsu_uncache [14]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [14]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b15  (
    .i0(\exu/n61 [15]),
    .i1(\exu/data_lsu_uncache [15]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [15]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b16  (
    .i0(\exu/n61 [16]),
    .i1(\exu/data_lsu_uncache [16]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [16]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b17  (
    .i0(\exu/n61 [17]),
    .i1(\exu/data_lsu_uncache [17]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [17]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b18  (
    .i0(\exu/n61 [18]),
    .i1(\exu/data_lsu_uncache [18]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [18]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b19  (
    .i0(\exu/n61 [19]),
    .i1(\exu/data_lsu_uncache [19]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [19]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b2  (
    .i0(\exu/n61 [2]),
    .i1(\exu/data_lsu_uncache [2]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [2]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b20  (
    .i0(\exu/n61 [20]),
    .i1(\exu/data_lsu_uncache [20]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [20]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b21  (
    .i0(\exu/n61 [21]),
    .i1(\exu/data_lsu_uncache [21]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [21]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b22  (
    .i0(\exu/n61 [22]),
    .i1(\exu/data_lsu_uncache [22]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [22]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b23  (
    .i0(\exu/n61 [23]),
    .i1(\exu/data_lsu_uncache [23]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [23]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b24  (
    .i0(\exu/n61 [24]),
    .i1(\exu/data_lsu_uncache [24]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [24]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b25  (
    .i0(\exu/n61 [25]),
    .i1(\exu/data_lsu_uncache [25]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [25]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b26  (
    .i0(\exu/n61 [26]),
    .i1(\exu/data_lsu_uncache [26]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [26]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b27  (
    .i0(\exu/n61 [27]),
    .i1(\exu/data_lsu_uncache [27]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [27]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b28  (
    .i0(\exu/n61 [28]),
    .i1(\exu/data_lsu_uncache [28]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [28]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b29  (
    .i0(\exu/n61 [29]),
    .i1(\exu/data_lsu_uncache [29]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [29]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b3  (
    .i0(\exu/n61 [3]),
    .i1(\exu/data_lsu_uncache [3]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [3]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b30  (
    .i0(\exu/n61 [30]),
    .i1(\exu/data_lsu_uncache [30]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [30]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b31  (
    .i0(\exu/n61 [31]),
    .i1(\exu/data_lsu_uncache [31]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [31]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b32  (
    .i0(\exu/n61 [32]),
    .i1(\exu/data_lsu_uncache [32]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [32]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b33  (
    .i0(\exu/n61 [33]),
    .i1(\exu/data_lsu_uncache [33]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [33]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b34  (
    .i0(\exu/n61 [34]),
    .i1(\exu/data_lsu_uncache [34]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [34]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b35  (
    .i0(\exu/n61 [35]),
    .i1(\exu/data_lsu_uncache [35]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [35]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b36  (
    .i0(\exu/n61 [36]),
    .i1(\exu/data_lsu_uncache [36]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [36]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b37  (
    .i0(\exu/n61 [37]),
    .i1(\exu/data_lsu_uncache [37]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [37]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b38  (
    .i0(\exu/n61 [38]),
    .i1(\exu/data_lsu_uncache [38]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [38]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b39  (
    .i0(\exu/n61 [39]),
    .i1(\exu/data_lsu_uncache [39]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [39]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b4  (
    .i0(\exu/n61 [4]),
    .i1(\exu/data_lsu_uncache [4]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [4]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b40  (
    .i0(\exu/n61 [40]),
    .i1(\exu/data_lsu_uncache [40]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [40]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b41  (
    .i0(\exu/n61 [41]),
    .i1(\exu/data_lsu_uncache [41]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [41]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b42  (
    .i0(\exu/n61 [42]),
    .i1(\exu/data_lsu_uncache [42]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [42]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b43  (
    .i0(\exu/n61 [43]),
    .i1(\exu/data_lsu_uncache [43]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [43]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b44  (
    .i0(\exu/n61 [44]),
    .i1(\exu/data_lsu_uncache [44]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [44]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b45  (
    .i0(\exu/n61 [45]),
    .i1(\exu/data_lsu_uncache [45]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [45]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b46  (
    .i0(\exu/n61 [46]),
    .i1(\exu/data_lsu_uncache [46]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [46]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b47  (
    .i0(\exu/n61 [47]),
    .i1(\exu/data_lsu_uncache [47]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [47]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b48  (
    .i0(\exu/n61 [48]),
    .i1(\exu/data_lsu_uncache [48]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [48]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b49  (
    .i0(\exu/n61 [49]),
    .i1(\exu/data_lsu_uncache [49]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [49]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b5  (
    .i0(\exu/n61 [5]),
    .i1(\exu/data_lsu_uncache [5]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [5]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b50  (
    .i0(\exu/n61 [50]),
    .i1(\exu/data_lsu_uncache [50]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [50]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b51  (
    .i0(\exu/n61 [51]),
    .i1(\exu/data_lsu_uncache [51]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [51]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b52  (
    .i0(\exu/n61 [52]),
    .i1(\exu/data_lsu_uncache [52]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [52]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b53  (
    .i0(\exu/n61 [53]),
    .i1(\exu/data_lsu_uncache [53]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [53]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b54  (
    .i0(\exu/n61 [54]),
    .i1(\exu/data_lsu_uncache [54]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [54]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b55  (
    .i0(\exu/n61 [55]),
    .i1(\exu/data_lsu_uncache [55]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [55]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b56  (
    .i0(\exu/n61 [56]),
    .i1(\exu/data_lsu_uncache [56]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [56]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b57  (
    .i0(\exu/n61 [57]),
    .i1(\exu/data_lsu_uncache [57]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [57]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b58  (
    .i0(\exu/n61 [58]),
    .i1(\exu/data_lsu_uncache [58]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [58]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b59  (
    .i0(\exu/n61 [59]),
    .i1(\exu/data_lsu_uncache [59]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [59]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b6  (
    .i0(\exu/n61 [6]),
    .i1(\exu/data_lsu_uncache [6]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [6]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b60  (
    .i0(\exu/n61 [60]),
    .i1(\exu/data_lsu_uncache [60]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [60]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b61  (
    .i0(\exu/n61 [61]),
    .i1(\exu/data_lsu_uncache [61]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [61]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b62  (
    .i0(\exu/n61 [62]),
    .i1(\exu/data_lsu_uncache [62]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [62]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b63  (
    .i0(\exu/n61 [63]),
    .i1(\exu/data_lsu_uncache [63]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [63]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b7  (
    .i0(\exu/n61 [7]),
    .i1(\exu/data_lsu_uncache [7]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [7]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b8  (
    .i0(\exu/n61 [8]),
    .i1(\exu/data_lsu_uncache [8]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [8]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux30_b9  (
    .i0(\exu/n61 [9]),
    .i1(\exu/data_lsu_uncache [9]),
    .sel(\exu/n59 ),
    .o(\exu/n62 [9]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b0  (
    .i0(\exu/n62 [0]),
    .i1(\exu/alu_au/n40 [0]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [0]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b1  (
    .i0(\exu/n62 [1]),
    .i1(\exu/alu_au/n38 [1]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [1]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b10  (
    .i0(\exu/n62 [10]),
    .i1(\exu/alu_au/n38 [10]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [10]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b11  (
    .i0(\exu/n62 [11]),
    .i1(\exu/alu_au/n38 [11]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [11]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b12  (
    .i0(\exu/n62 [12]),
    .i1(\exu/alu_au/n38 [12]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [12]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b13  (
    .i0(\exu/n62 [13]),
    .i1(\exu/alu_au/n38 [13]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [13]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b14  (
    .i0(\exu/n62 [14]),
    .i1(\exu/alu_au/n38 [14]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [14]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b15  (
    .i0(\exu/n62 [15]),
    .i1(\exu/alu_au/n38 [15]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [15]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b16  (
    .i0(\exu/n62 [16]),
    .i1(\exu/alu_au/n38 [16]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [16]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b17  (
    .i0(\exu/n62 [17]),
    .i1(\exu/alu_au/n38 [17]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [17]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b18  (
    .i0(\exu/n62 [18]),
    .i1(\exu/alu_au/n38 [18]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [18]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b19  (
    .i0(\exu/n62 [19]),
    .i1(\exu/alu_au/n38 [19]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [19]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b2  (
    .i0(\exu/n62 [2]),
    .i1(\exu/alu_au/n38 [2]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [2]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b20  (
    .i0(\exu/n62 [20]),
    .i1(\exu/alu_au/n38 [20]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [20]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b21  (
    .i0(\exu/n62 [21]),
    .i1(\exu/alu_au/n38 [21]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [21]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b22  (
    .i0(\exu/n62 [22]),
    .i1(\exu/alu_au/n38 [22]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [22]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b23  (
    .i0(\exu/n62 [23]),
    .i1(\exu/alu_au/n38 [23]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [23]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b24  (
    .i0(\exu/n62 [24]),
    .i1(\exu/alu_au/n38 [24]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [24]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b25  (
    .i0(\exu/n62 [25]),
    .i1(\exu/alu_au/n38 [25]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [25]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b26  (
    .i0(\exu/n62 [26]),
    .i1(\exu/alu_au/n38 [26]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [26]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b27  (
    .i0(\exu/n62 [27]),
    .i1(\exu/alu_au/n38 [27]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [27]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b28  (
    .i0(\exu/n62 [28]),
    .i1(\exu/alu_au/n38 [28]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [28]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b29  (
    .i0(\exu/n62 [29]),
    .i1(\exu/alu_au/n38 [29]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [29]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b3  (
    .i0(\exu/n62 [3]),
    .i1(\exu/alu_au/n38 [3]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [3]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b30  (
    .i0(\exu/n62 [30]),
    .i1(\exu/alu_au/n38 [30]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [30]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b31  (
    .i0(\exu/n62 [31]),
    .i1(\exu/alu_au/n38 [31]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [31]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b32  (
    .i0(\exu/n62 [32]),
    .i1(\exu/alu_au/n38 [32]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [32]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b33  (
    .i0(\exu/n62 [33]),
    .i1(\exu/alu_au/n38 [33]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [33]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b34  (
    .i0(\exu/n62 [34]),
    .i1(\exu/alu_au/n38 [34]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [34]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b35  (
    .i0(\exu/n62 [35]),
    .i1(\exu/alu_au/n38 [35]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [35]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b36  (
    .i0(\exu/n62 [36]),
    .i1(\exu/alu_au/n38 [36]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [36]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b37  (
    .i0(\exu/n62 [37]),
    .i1(\exu/alu_au/n38 [37]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [37]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b38  (
    .i0(\exu/n62 [38]),
    .i1(\exu/alu_au/n38 [38]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [38]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b39  (
    .i0(\exu/n62 [39]),
    .i1(\exu/alu_au/n38 [39]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [39]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b4  (
    .i0(\exu/n62 [4]),
    .i1(\exu/alu_au/n38 [4]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [4]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b40  (
    .i0(\exu/n62 [40]),
    .i1(\exu/alu_au/n38 [40]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [40]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b41  (
    .i0(\exu/n62 [41]),
    .i1(\exu/alu_au/n38 [41]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [41]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b42  (
    .i0(\exu/n62 [42]),
    .i1(\exu/alu_au/n38 [42]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [42]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b43  (
    .i0(\exu/n62 [43]),
    .i1(\exu/alu_au/n38 [43]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [43]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b44  (
    .i0(\exu/n62 [44]),
    .i1(\exu/alu_au/n38 [44]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [44]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b45  (
    .i0(\exu/n62 [45]),
    .i1(\exu/alu_au/n38 [45]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [45]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b46  (
    .i0(\exu/n62 [46]),
    .i1(\exu/alu_au/n38 [46]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [46]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b47  (
    .i0(\exu/n62 [47]),
    .i1(\exu/alu_au/n38 [47]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [47]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b48  (
    .i0(\exu/n62 [48]),
    .i1(\exu/alu_au/n38 [48]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [48]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b49  (
    .i0(\exu/n62 [49]),
    .i1(\exu/alu_au/n38 [49]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [49]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b5  (
    .i0(\exu/n62 [5]),
    .i1(\exu/alu_au/n38 [5]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [5]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b50  (
    .i0(\exu/n62 [50]),
    .i1(\exu/alu_au/n38 [50]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [50]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b51  (
    .i0(\exu/n62 [51]),
    .i1(\exu/alu_au/n38 [51]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [51]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b52  (
    .i0(\exu/n62 [52]),
    .i1(\exu/alu_au/n38 [52]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [52]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b53  (
    .i0(\exu/n62 [53]),
    .i1(\exu/alu_au/n38 [53]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [53]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b54  (
    .i0(\exu/n62 [54]),
    .i1(\exu/alu_au/n38 [54]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [54]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b55  (
    .i0(\exu/n62 [55]),
    .i1(\exu/alu_au/n38 [55]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [55]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b56  (
    .i0(\exu/n62 [56]),
    .i1(\exu/alu_au/n38 [56]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [56]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b57  (
    .i0(\exu/n62 [57]),
    .i1(\exu/alu_au/n38 [57]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [57]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b58  (
    .i0(\exu/n62 [58]),
    .i1(\exu/alu_au/n38 [58]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [58]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b59  (
    .i0(\exu/n62 [59]),
    .i1(\exu/alu_au/n38 [59]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [59]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b6  (
    .i0(\exu/n62 [6]),
    .i1(\exu/alu_au/n38 [6]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [6]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b60  (
    .i0(\exu/n62 [60]),
    .i1(\exu/alu_au/n38 [60]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [60]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b61  (
    .i0(\exu/n62 [61]),
    .i1(\exu/alu_au/n38 [61]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [61]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b62  (
    .i0(\exu/n62 [62]),
    .i1(\exu/alu_au/n38 [62]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [62]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b63  (
    .i0(\exu/n62 [63]),
    .i1(\exu/alu_au/n38 [63]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [63]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b7  (
    .i0(\exu/n62 [7]),
    .i1(\exu/alu_au/n38 [7]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [7]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b8  (
    .i0(\exu/n62 [8]),
    .i1(\exu/alu_au/n38 [8]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [8]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux31_b9  (
    .i0(\exu/n62 [9]),
    .i1(\exu/alu_au/n38 [9]),
    .sel(\exu/c_stb ),
    .o(\exu/n63 [9]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b0  (
    .i0(\exu/n63 [0]),
    .i1(\exu/n58 [0]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [0]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b1  (
    .i0(\exu/n63 [1]),
    .i1(\exu/n58 [1]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [1]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b10  (
    .i0(\exu/n63 [10]),
    .i1(\exu/n58 [10]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [10]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b11  (
    .i0(\exu/n63 [11]),
    .i1(\exu/n58 [11]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [11]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b12  (
    .i0(\exu/n63 [12]),
    .i1(\exu/n58 [12]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [12]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b13  (
    .i0(\exu/n63 [13]),
    .i1(\exu/n58 [13]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [13]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b14  (
    .i0(\exu/n63 [14]),
    .i1(\exu/n58 [14]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [14]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b15  (
    .i0(\exu/n63 [15]),
    .i1(\exu/n58 [15]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [15]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b16  (
    .i0(\exu/n63 [16]),
    .i1(\exu/n58 [16]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [16]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b17  (
    .i0(\exu/n63 [17]),
    .i1(\exu/n58 [17]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [17]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b18  (
    .i0(\exu/n63 [18]),
    .i1(\exu/n58 [18]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [18]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b19  (
    .i0(\exu/n63 [19]),
    .i1(\exu/n58 [19]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [19]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b2  (
    .i0(\exu/n63 [2]),
    .i1(\exu/n58 [2]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [2]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b20  (
    .i0(\exu/n63 [20]),
    .i1(\exu/n58 [20]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [20]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b21  (
    .i0(\exu/n63 [21]),
    .i1(\exu/n58 [21]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [21]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b22  (
    .i0(\exu/n63 [22]),
    .i1(\exu/n58 [22]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [22]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b23  (
    .i0(\exu/n63 [23]),
    .i1(\exu/n58 [23]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [23]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b24  (
    .i0(\exu/n63 [24]),
    .i1(\exu/n58 [24]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [24]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b25  (
    .i0(\exu/n63 [25]),
    .i1(\exu/n58 [25]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [25]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b26  (
    .i0(\exu/n63 [26]),
    .i1(\exu/n58 [26]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [26]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b27  (
    .i0(\exu/n63 [27]),
    .i1(\exu/n58 [27]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [27]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b28  (
    .i0(\exu/n63 [28]),
    .i1(\exu/n58 [28]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [28]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b29  (
    .i0(\exu/n63 [29]),
    .i1(\exu/n58 [29]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [29]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b3  (
    .i0(\exu/n63 [3]),
    .i1(\exu/n58 [3]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [3]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b30  (
    .i0(\exu/n63 [30]),
    .i1(\exu/n58 [30]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [30]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b31  (
    .i0(\exu/n63 [31]),
    .i1(\exu/n58 [31]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [31]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b32  (
    .i0(\exu/n63 [32]),
    .i1(\exu/n58 [32]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [32]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b33  (
    .i0(\exu/n63 [33]),
    .i1(\exu/n58 [33]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [33]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b34  (
    .i0(\exu/n63 [34]),
    .i1(\exu/n58 [34]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [34]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b35  (
    .i0(\exu/n63 [35]),
    .i1(\exu/n58 [35]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [35]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b36  (
    .i0(\exu/n63 [36]),
    .i1(\exu/n58 [36]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [36]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b37  (
    .i0(\exu/n63 [37]),
    .i1(\exu/n58 [37]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [37]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b38  (
    .i0(\exu/n63 [38]),
    .i1(\exu/n58 [38]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [38]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b39  (
    .i0(\exu/n63 [39]),
    .i1(\exu/n58 [39]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [39]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b4  (
    .i0(\exu/n63 [4]),
    .i1(\exu/n58 [4]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [4]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b40  (
    .i0(\exu/n63 [40]),
    .i1(\exu/n58 [40]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [40]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b41  (
    .i0(\exu/n63 [41]),
    .i1(\exu/n58 [41]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [41]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b42  (
    .i0(\exu/n63 [42]),
    .i1(\exu/n58 [42]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [42]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b43  (
    .i0(\exu/n63 [43]),
    .i1(\exu/n58 [43]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [43]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b44  (
    .i0(\exu/n63 [44]),
    .i1(\exu/n58 [44]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [44]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b45  (
    .i0(\exu/n63 [45]),
    .i1(\exu/n58 [45]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [45]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b46  (
    .i0(\exu/n63 [46]),
    .i1(\exu/n58 [46]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [46]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b47  (
    .i0(\exu/n63 [47]),
    .i1(\exu/n58 [47]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [47]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b48  (
    .i0(\exu/n63 [48]),
    .i1(\exu/n58 [48]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [48]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b49  (
    .i0(\exu/n63 [49]),
    .i1(\exu/n58 [49]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [49]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b5  (
    .i0(\exu/n63 [5]),
    .i1(\exu/n58 [5]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [5]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b50  (
    .i0(\exu/n63 [50]),
    .i1(\exu/n58 [50]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [50]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b51  (
    .i0(\exu/n63 [51]),
    .i1(\exu/n58 [51]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [51]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b52  (
    .i0(\exu/n63 [52]),
    .i1(\exu/n58 [52]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [52]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b53  (
    .i0(\exu/n63 [53]),
    .i1(\exu/n58 [53]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [53]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b54  (
    .i0(\exu/n63 [54]),
    .i1(\exu/n58 [54]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [54]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b55  (
    .i0(\exu/n63 [55]),
    .i1(\exu/n58 [55]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [55]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b56  (
    .i0(\exu/n63 [56]),
    .i1(\exu/n58 [56]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [56]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b57  (
    .i0(\exu/n63 [57]),
    .i1(\exu/n58 [57]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [57]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b58  (
    .i0(\exu/n63 [58]),
    .i1(\exu/n58 [58]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [58]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b59  (
    .i0(\exu/n63 [59]),
    .i1(\exu/n58 [59]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [59]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b6  (
    .i0(\exu/n63 [6]),
    .i1(\exu/n58 [6]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [6]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b60  (
    .i0(\exu/n63 [60]),
    .i1(\exu/n58 [60]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [60]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b61  (
    .i0(\exu/n63 [61]),
    .i1(\exu/n58 [61]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [61]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b62  (
    .i0(\exu/n63 [62]),
    .i1(\exu/n58 [62]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [62]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b63  (
    .i0(\exu/n63 [63]),
    .i1(\exu/n58 [63]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [63]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b7  (
    .i0(\exu/n63 [7]),
    .i1(\exu/n58 [7]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [7]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b8  (
    .i0(\exu/n63 [8]),
    .i1(\exu/n58 [8]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [8]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux32_b9  (
    .i0(\exu/n63 [9]),
    .i1(\exu/n58 [9]),
    .sel(\exu/c_shift ),
    .o(\exu/n64 [9]));  // ../../RTL/CPU/EX/exu.v(326)
  binary_mux_s1_w1 \exu/mux39_b0  (
    .i0(ex_exc_code[0]),
    .i1(addr_ex[0]),
    .sel(ex_more_exception),
    .o(\exu/n71 [0]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b1  (
    .i0(ex_exc_code[1]),
    .i1(addr_ex[1]),
    .sel(ex_more_exception),
    .o(\exu/n71 [1]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b10  (
    .i0(ex_exc_code[10]),
    .i1(addr_ex[10]),
    .sel(ex_more_exception),
    .o(\exu/n71 [10]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b11  (
    .i0(ex_exc_code[11]),
    .i1(addr_ex[11]),
    .sel(ex_more_exception),
    .o(\exu/n71 [11]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b12  (
    .i0(ex_exc_code[12]),
    .i1(addr_ex[12]),
    .sel(ex_more_exception),
    .o(\exu/n71 [12]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b13  (
    .i0(ex_exc_code[13]),
    .i1(addr_ex[13]),
    .sel(ex_more_exception),
    .o(\exu/n71 [13]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b14  (
    .i0(ex_exc_code[14]),
    .i1(addr_ex[14]),
    .sel(ex_more_exception),
    .o(\exu/n71 [14]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b15  (
    .i0(ex_exc_code[15]),
    .i1(addr_ex[15]),
    .sel(ex_more_exception),
    .o(\exu/n71 [15]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b16  (
    .i0(ex_exc_code[16]),
    .i1(addr_ex[16]),
    .sel(ex_more_exception),
    .o(\exu/n71 [16]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b17  (
    .i0(ex_exc_code[17]),
    .i1(addr_ex[17]),
    .sel(ex_more_exception),
    .o(\exu/n71 [17]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b18  (
    .i0(ex_exc_code[18]),
    .i1(addr_ex[18]),
    .sel(ex_more_exception),
    .o(\exu/n71 [18]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b19  (
    .i0(ex_exc_code[19]),
    .i1(addr_ex[19]),
    .sel(ex_more_exception),
    .o(\exu/n71 [19]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b2  (
    .i0(ex_exc_code[2]),
    .i1(addr_ex[2]),
    .sel(ex_more_exception),
    .o(\exu/n71 [2]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b20  (
    .i0(ex_exc_code[20]),
    .i1(addr_ex[20]),
    .sel(ex_more_exception),
    .o(\exu/n71 [20]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b21  (
    .i0(ex_exc_code[21]),
    .i1(addr_ex[21]),
    .sel(ex_more_exception),
    .o(\exu/n71 [21]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b22  (
    .i0(ex_exc_code[22]),
    .i1(addr_ex[22]),
    .sel(ex_more_exception),
    .o(\exu/n71 [22]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b23  (
    .i0(ex_exc_code[23]),
    .i1(addr_ex[23]),
    .sel(ex_more_exception),
    .o(\exu/n71 [23]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b24  (
    .i0(ex_exc_code[24]),
    .i1(addr_ex[24]),
    .sel(ex_more_exception),
    .o(\exu/n71 [24]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b25  (
    .i0(ex_exc_code[25]),
    .i1(addr_ex[25]),
    .sel(ex_more_exception),
    .o(\exu/n71 [25]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b26  (
    .i0(ex_exc_code[26]),
    .i1(addr_ex[26]),
    .sel(ex_more_exception),
    .o(\exu/n71 [26]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b27  (
    .i0(ex_exc_code[27]),
    .i1(addr_ex[27]),
    .sel(ex_more_exception),
    .o(\exu/n71 [27]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b28  (
    .i0(ex_exc_code[28]),
    .i1(addr_ex[28]),
    .sel(ex_more_exception),
    .o(\exu/n71 [28]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b29  (
    .i0(ex_exc_code[29]),
    .i1(addr_ex[29]),
    .sel(ex_more_exception),
    .o(\exu/n71 [29]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b3  (
    .i0(ex_exc_code[3]),
    .i1(addr_ex[3]),
    .sel(ex_more_exception),
    .o(\exu/n71 [3]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b30  (
    .i0(ex_exc_code[30]),
    .i1(addr_ex[30]),
    .sel(ex_more_exception),
    .o(\exu/n71 [30]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b31  (
    .i0(ex_exc_code[31]),
    .i1(addr_ex[31]),
    .sel(ex_more_exception),
    .o(\exu/n71 [31]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b32  (
    .i0(1'b0),
    .i1(addr_ex[32]),
    .sel(ex_more_exception),
    .o(\exu/n71 [32]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b33  (
    .i0(1'b0),
    .i1(addr_ex[33]),
    .sel(ex_more_exception),
    .o(\exu/n71 [33]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b34  (
    .i0(1'b0),
    .i1(addr_ex[34]),
    .sel(ex_more_exception),
    .o(\exu/n71 [34]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b35  (
    .i0(1'b0),
    .i1(addr_ex[35]),
    .sel(ex_more_exception),
    .o(\exu/n71 [35]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b36  (
    .i0(1'b0),
    .i1(addr_ex[36]),
    .sel(ex_more_exception),
    .o(\exu/n71 [36]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b37  (
    .i0(1'b0),
    .i1(addr_ex[37]),
    .sel(ex_more_exception),
    .o(\exu/n71 [37]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b38  (
    .i0(1'b0),
    .i1(addr_ex[38]),
    .sel(ex_more_exception),
    .o(\exu/n71 [38]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b39  (
    .i0(1'b0),
    .i1(addr_ex[39]),
    .sel(ex_more_exception),
    .o(\exu/n71 [39]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b4  (
    .i0(ex_exc_code[4]),
    .i1(addr_ex[4]),
    .sel(ex_more_exception),
    .o(\exu/n71 [4]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b40  (
    .i0(1'b0),
    .i1(addr_ex[40]),
    .sel(ex_more_exception),
    .o(\exu/n71 [40]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b41  (
    .i0(1'b0),
    .i1(addr_ex[41]),
    .sel(ex_more_exception),
    .o(\exu/n71 [41]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b42  (
    .i0(1'b0),
    .i1(addr_ex[42]),
    .sel(ex_more_exception),
    .o(\exu/n71 [42]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b43  (
    .i0(1'b0),
    .i1(addr_ex[43]),
    .sel(ex_more_exception),
    .o(\exu/n71 [43]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b44  (
    .i0(1'b0),
    .i1(addr_ex[44]),
    .sel(ex_more_exception),
    .o(\exu/n71 [44]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b45  (
    .i0(1'b0),
    .i1(addr_ex[45]),
    .sel(ex_more_exception),
    .o(\exu/n71 [45]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b46  (
    .i0(1'b0),
    .i1(addr_ex[46]),
    .sel(ex_more_exception),
    .o(\exu/n71 [46]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b47  (
    .i0(1'b0),
    .i1(addr_ex[47]),
    .sel(ex_more_exception),
    .o(\exu/n71 [47]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b48  (
    .i0(1'b0),
    .i1(addr_ex[48]),
    .sel(ex_more_exception),
    .o(\exu/n71 [48]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b49  (
    .i0(1'b0),
    .i1(addr_ex[49]),
    .sel(ex_more_exception),
    .o(\exu/n71 [49]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b5  (
    .i0(ex_exc_code[5]),
    .i1(addr_ex[5]),
    .sel(ex_more_exception),
    .o(\exu/n71 [5]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b50  (
    .i0(1'b0),
    .i1(addr_ex[50]),
    .sel(ex_more_exception),
    .o(\exu/n71 [50]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b51  (
    .i0(1'b0),
    .i1(addr_ex[51]),
    .sel(ex_more_exception),
    .o(\exu/n71 [51]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b52  (
    .i0(1'b0),
    .i1(addr_ex[52]),
    .sel(ex_more_exception),
    .o(\exu/n71 [52]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b53  (
    .i0(1'b0),
    .i1(addr_ex[53]),
    .sel(ex_more_exception),
    .o(\exu/n71 [53]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b54  (
    .i0(1'b0),
    .i1(addr_ex[54]),
    .sel(ex_more_exception),
    .o(\exu/n71 [54]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b55  (
    .i0(1'b0),
    .i1(addr_ex[55]),
    .sel(ex_more_exception),
    .o(\exu/n71 [55]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b56  (
    .i0(1'b0),
    .i1(addr_ex[56]),
    .sel(ex_more_exception),
    .o(\exu/n71 [56]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b57  (
    .i0(1'b0),
    .i1(addr_ex[57]),
    .sel(ex_more_exception),
    .o(\exu/n71 [57]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b58  (
    .i0(1'b0),
    .i1(addr_ex[58]),
    .sel(ex_more_exception),
    .o(\exu/n71 [58]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b59  (
    .i0(1'b0),
    .i1(addr_ex[59]),
    .sel(ex_more_exception),
    .o(\exu/n71 [59]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b6  (
    .i0(ex_exc_code[6]),
    .i1(addr_ex[6]),
    .sel(ex_more_exception),
    .o(\exu/n71 [6]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b60  (
    .i0(1'b0),
    .i1(addr_ex[60]),
    .sel(ex_more_exception),
    .o(\exu/n71 [60]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b61  (
    .i0(1'b0),
    .i1(addr_ex[61]),
    .sel(ex_more_exception),
    .o(\exu/n71 [61]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b62  (
    .i0(1'b0),
    .i1(addr_ex[62]),
    .sel(ex_more_exception),
    .o(\exu/n71 [62]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b63  (
    .i0(1'b0),
    .i1(addr_ex[63]),
    .sel(ex_more_exception),
    .o(\exu/n71 [63]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b7  (
    .i0(ex_exc_code[7]),
    .i1(addr_ex[7]),
    .sel(ex_more_exception),
    .o(\exu/n71 [7]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b8  (
    .i0(ex_exc_code[8]),
    .i1(addr_ex[8]),
    .sel(ex_more_exception),
    .o(\exu/n71 [8]));  // ../../RTL/CPU/EX/exu.v(356)
  binary_mux_s1_w1 \exu/mux39_b9  (
    .i0(ex_exc_code[9]),
    .i1(addr_ex[9]),
    .sel(ex_more_exception),
    .o(\exu/n71 [9]));  // ../../RTL/CPU/EX/exu.v(356)
  AL_MUX \exu/mux3_b1  (
    .i0(1'b0),
    .i1(\exu/main_state [1]),
    .sel(\exu/mux3_b1_sel_is_2_o ),
    .o(\exu/n25 [1]));
  and \exu/mux3_b1_sel_is_2  (\exu/mux3_b1_sel_is_2_o , store_neg, \exu/mux2_b1_sel_is_2_o );
  binary_mux_s1_w1 \exu/mux3_b2  (
    .i0(\exu/n24 [2]),
    .i1(1'b1),
    .sel(store),
    .o(\exu/n25 [2]));  // ../../RTL/CPU/EX/exu.v(240)
  and \exu/mux3_b3_sel_is_0  (\exu/mux3_b3_sel_is_0_o , store_neg, \exu/n20_neg );
  binary_mux_s1_w1 \exu/mux48_b0  (
    .i0(\exu/n55 [33]),
    .i1(\exu/n55 [0]),
    .sel(unsign),
    .o(\exu/n56 [0]));  // ../../RTL/CPU/EX/exu.v(311)
  and \exu/mux48_b32_sel_is_1  (\exu/mux48_b32_sel_is_1_o , unsign, \ex_size[2]_neg );
  binary_mux_s1_w1 \exu/mux49_b0  (
    .i0(priv[0]),
    .i1(mod_priv[0]),
    .sel(unpage),
    .o(ex_priv[0]));  // ../../RTL/CPU/EX/exu.v(507)
  binary_mux_s1_w1 \exu/mux49_b1  (
    .i0(priv[1]),
    .i1(mod_priv[1]),
    .sel(unpage),
    .o(ex_priv[1]));  // ../../RTL/CPU/EX/exu.v(507)
  binary_mux_s1_w1 \exu/mux49_b3  (
    .i0(priv[3]),
    .i1(mod_priv[3]),
    .sel(unpage),
    .o(ex_priv[3]));  // ../../RTL/CPU/EX/exu.v(507)
  AL_MUX \exu/mux4_b0  (
    .i0(1'b0),
    .i1(\exu/n24 [0]),
    .sel(\exu/mux4_b0_sel_is_0_o ),
    .o(\exu/n26 [0]));
  and \exu/mux4_b0_sel_is_0  (\exu/mux4_b0_sel_is_0_o , load_neg, store_neg);
  binary_mux_s1_w1 \exu/mux4_b1  (
    .i0(\exu/n25 [1]),
    .i1(1'b1),
    .sel(load),
    .o(\exu/n26 [1]));  // ../../RTL/CPU/EX/exu.v(240)
  binary_mux_s1_w1 \exu/mux4_b2  (
    .i0(\exu/n25 [2]),
    .i1(1'b0),
    .sel(load),
    .o(\exu/n26 [2]));  // ../../RTL/CPU/EX/exu.v(240)
  AL_MUX \exu/mux4_b3  (
    .i0(1'b0),
    .i1(\exu/n23 [3]),
    .sel(\exu/mux4_b3_sel_is_2_o ),
    .o(\exu/n26 [3]));
  and \exu/mux4_b3_sel_is_2  (\exu/mux4_b3_sel_is_2_o , load_neg, \exu/mux3_b3_sel_is_0_o );
  binary_mux_s1_w1 \exu/mux5_b0  (
    .i0(cache_ready_ex),
    .i1(1'b0),
    .sel(uncache_data_rdy),
    .o(\exu/n27 [0]));  // ../../RTL/CPU/EX/exu.v(244)
  binary_mux_s1_w1 \exu/mux5_b1  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(uncache_data_rdy),
    .o(\exu/n27 [1]));  // ../../RTL/CPU/EX/exu.v(244)
  binary_mux_s1_w1 \exu/mux8_b0  (
    .i0(\exu/n27 [0]),
    .i1(1'b0),
    .sel(ex_more_exception),
    .o(\exu/n33 [0]));  // ../../RTL/CPU/EX/exu.v(253)
  AL_MUX \exu/mux8_b1  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\exu/mux8_b1_sel_is_2_o ),
    .o(\exu/n33 [1]));
  and \exu/mux8_b1_sel_is_2  (\exu/mux8_b1_sel_is_2_o , ex_more_exception_neg, uncache_data_rdy);
  binary_mux_s1_w1 \exu/mux8_b3  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(ex_more_exception),
    .o(\exu/n33 [3]));  // ../../RTL/CPU/EX/exu.v(253)
  not \exu/n20_inv  (\exu/n20_neg , \exu/n20 );
  not \exu/n21_inv  (\exu/n21_neg , \exu/n21 );
  not \exu/n35_inv  (\exu/n35_neg , \exu/n35 );
  ne_w2 \exu/neq0  (
    .i0(addr_ex[1:0]),
    .i1(2'b00),
    .o(\exu/n3 ));  // ../../RTL/CPU/EX/exu.v(211)
  ne_w3 \exu/neq1  (
    .i0(addr_ex[2:0]),
    .i1(3'b000),
    .o(\exu/n6 ));  // ../../RTL/CPU/EX/exu.v(211)
  reg_sr_as_w1 \exu/pc_jmp_reg  (
    .clk(clk),
    .d(jmp),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(pc_jmp));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg0_b0  (
    .clk(clk),
    .d(\exu/n52 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\exu/shift_count [0]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b1  (
    .clk(clk),
    .d(\exu/n52 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\exu/shift_count [1]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b2  (
    .clk(clk),
    .d(\exu/n52 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\exu/shift_count [2]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b3  (
    .clk(clk),
    .d(\exu/n52 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\exu/shift_count [3]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b4  (
    .clk(clk),
    .d(\exu/n52 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\exu/shift_count [4]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b5  (
    .clk(clk),
    .d(\exu/n52 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\exu/shift_count [5]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b6  (
    .clk(clk),
    .d(\exu/n52 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\exu/shift_count [6]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg0_b7  (
    .clk(clk),
    .d(\exu/n52 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(\exu/shift_count [7]));  // ../../RTL/CPU/EX/exu.v(290)
  reg_sr_as_w1 \exu/reg1_b0  (
    .clk(clk),
    .d(\exu/n64 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[0]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b1  (
    .clk(clk),
    .d(\exu/n64 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[1]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b10  (
    .clk(clk),
    .d(\exu/n64 [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[10]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b11  (
    .clk(clk),
    .d(\exu/n64 [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[11]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b12  (
    .clk(clk),
    .d(\exu/n64 [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[12]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b13  (
    .clk(clk),
    .d(\exu/n64 [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[13]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b14  (
    .clk(clk),
    .d(\exu/n64 [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[14]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b15  (
    .clk(clk),
    .d(\exu/n64 [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[15]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b16  (
    .clk(clk),
    .d(\exu/n64 [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[16]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b17  (
    .clk(clk),
    .d(\exu/n64 [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[17]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b18  (
    .clk(clk),
    .d(\exu/n64 [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[18]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b19  (
    .clk(clk),
    .d(\exu/n64 [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[19]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b2  (
    .clk(clk),
    .d(\exu/n64 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[2]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b20  (
    .clk(clk),
    .d(\exu/n64 [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[20]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b21  (
    .clk(clk),
    .d(\exu/n64 [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[21]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b22  (
    .clk(clk),
    .d(\exu/n64 [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[22]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b23  (
    .clk(clk),
    .d(\exu/n64 [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[23]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b24  (
    .clk(clk),
    .d(\exu/n64 [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[24]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b25  (
    .clk(clk),
    .d(\exu/n64 [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[25]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b26  (
    .clk(clk),
    .d(\exu/n64 [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[26]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b27  (
    .clk(clk),
    .d(\exu/n64 [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[27]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b28  (
    .clk(clk),
    .d(\exu/n64 [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[28]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b29  (
    .clk(clk),
    .d(\exu/n64 [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[29]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b3  (
    .clk(clk),
    .d(\exu/n64 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[3]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b30  (
    .clk(clk),
    .d(\exu/n64 [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[30]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b31  (
    .clk(clk),
    .d(\exu/n64 [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[31]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b32  (
    .clk(clk),
    .d(\exu/n64 [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[32]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b33  (
    .clk(clk),
    .d(\exu/n64 [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[33]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b34  (
    .clk(clk),
    .d(\exu/n64 [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[34]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b35  (
    .clk(clk),
    .d(\exu/n64 [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[35]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b36  (
    .clk(clk),
    .d(\exu/n64 [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[36]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b37  (
    .clk(clk),
    .d(\exu/n64 [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[37]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b38  (
    .clk(clk),
    .d(\exu/n64 [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[38]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b39  (
    .clk(clk),
    .d(\exu/n64 [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[39]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b4  (
    .clk(clk),
    .d(\exu/n64 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[4]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b40  (
    .clk(clk),
    .d(\exu/n64 [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[40]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b41  (
    .clk(clk),
    .d(\exu/n64 [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[41]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b42  (
    .clk(clk),
    .d(\exu/n64 [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[42]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b43  (
    .clk(clk),
    .d(\exu/n64 [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[43]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b44  (
    .clk(clk),
    .d(\exu/n64 [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[44]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b45  (
    .clk(clk),
    .d(\exu/n64 [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[45]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b46  (
    .clk(clk),
    .d(\exu/n64 [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[46]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b47  (
    .clk(clk),
    .d(\exu/n64 [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[47]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b48  (
    .clk(clk),
    .d(\exu/n64 [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[48]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b49  (
    .clk(clk),
    .d(\exu/n64 [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[49]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b5  (
    .clk(clk),
    .d(\exu/n64 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[5]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b50  (
    .clk(clk),
    .d(\exu/n64 [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[50]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b51  (
    .clk(clk),
    .d(\exu/n64 [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[51]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b52  (
    .clk(clk),
    .d(\exu/n64 [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[52]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b53  (
    .clk(clk),
    .d(\exu/n64 [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[53]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b54  (
    .clk(clk),
    .d(\exu/n64 [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[54]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b55  (
    .clk(clk),
    .d(\exu/n64 [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[55]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b56  (
    .clk(clk),
    .d(\exu/n64 [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[56]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b57  (
    .clk(clk),
    .d(\exu/n64 [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[57]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b58  (
    .clk(clk),
    .d(\exu/n64 [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[58]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b59  (
    .clk(clk),
    .d(\exu/n64 [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[59]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b6  (
    .clk(clk),
    .d(\exu/n64 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[6]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b60  (
    .clk(clk),
    .d(\exu/n64 [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[60]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b61  (
    .clk(clk),
    .d(\exu/n64 [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[61]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b62  (
    .clk(clk),
    .d(\exu/n64 [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[62]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b63  (
    .clk(clk),
    .d(\exu/n64 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[63]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b7  (
    .clk(clk),
    .d(\exu/n64 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[7]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b8  (
    .clk(clk),
    .d(\exu/n64 [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[8]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg1_b9  (
    .clk(clk),
    .d(\exu/n64 [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_rd[9]));  // ../../RTL/CPU/EX/exu.v(327)
  reg_sr_as_w1 \exu/reg2_b0  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[0]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b1  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[1]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b10  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[10]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b11  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[11]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b12  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[12]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b13  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[13]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b14  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[14]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b15  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[15]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b16  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[16]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b17  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[17]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b18  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[18]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b19  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[19]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b2  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[2]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b20  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[20]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b21  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[21]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b22  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[22]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b23  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[23]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b24  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[24]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b25  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[25]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b26  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[26]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b27  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[27]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b28  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[28]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b29  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[29]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b3  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[3]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b30  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[30]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b31  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[31]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b32  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[32]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b33  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[33]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b34  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[34]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b35  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[35]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b36  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[36]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b37  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[37]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b38  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[38]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b39  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[39]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b4  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[4]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b40  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[40]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b41  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[41]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b42  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[42]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b43  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[43]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b44  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[44]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b45  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[45]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b46  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[46]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b47  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[47]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b48  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[48]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b49  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[49]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b5  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[5]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b50  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[50]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b51  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[51]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b52  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[52]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b53  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[53]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b54  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[54]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b55  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[55]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b56  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[56]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b57  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[57]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b58  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[58]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b59  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[59]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b6  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[6]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b60  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[60]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b61  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[61]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b62  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[62]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b63  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[63]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b7  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[7]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b8  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[8]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg2_b9  (
    .clk(clk),
    .d(\exu/alu_data_mem_csr [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(data_csr[9]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b0  (
    .clk(clk),
    .d(addr_ex[0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[0]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b1  (
    .clk(clk),
    .d(addr_ex[1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[1]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b10  (
    .clk(clk),
    .d(addr_ex[10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[10]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b11  (
    .clk(clk),
    .d(addr_ex[11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[11]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b12  (
    .clk(clk),
    .d(addr_ex[12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[12]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b13  (
    .clk(clk),
    .d(addr_ex[13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[13]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b14  (
    .clk(clk),
    .d(addr_ex[14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[14]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b15  (
    .clk(clk),
    .d(addr_ex[15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[15]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b16  (
    .clk(clk),
    .d(addr_ex[16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[16]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b17  (
    .clk(clk),
    .d(addr_ex[17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[17]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b18  (
    .clk(clk),
    .d(addr_ex[18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[18]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b19  (
    .clk(clk),
    .d(addr_ex[19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[19]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b2  (
    .clk(clk),
    .d(addr_ex[2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[2]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b20  (
    .clk(clk),
    .d(addr_ex[20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[20]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b21  (
    .clk(clk),
    .d(addr_ex[21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[21]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b22  (
    .clk(clk),
    .d(addr_ex[22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[22]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b23  (
    .clk(clk),
    .d(addr_ex[23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[23]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b24  (
    .clk(clk),
    .d(addr_ex[24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[24]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b25  (
    .clk(clk),
    .d(addr_ex[25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[25]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b26  (
    .clk(clk),
    .d(addr_ex[26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[26]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b27  (
    .clk(clk),
    .d(addr_ex[27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[27]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b28  (
    .clk(clk),
    .d(addr_ex[28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[28]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b29  (
    .clk(clk),
    .d(addr_ex[29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[29]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b3  (
    .clk(clk),
    .d(addr_ex[3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[3]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b30  (
    .clk(clk),
    .d(addr_ex[30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[30]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b31  (
    .clk(clk),
    .d(addr_ex[31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[31]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b32  (
    .clk(clk),
    .d(addr_ex[32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[32]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b33  (
    .clk(clk),
    .d(addr_ex[33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[33]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b34  (
    .clk(clk),
    .d(addr_ex[34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[34]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b35  (
    .clk(clk),
    .d(addr_ex[35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[35]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b36  (
    .clk(clk),
    .d(addr_ex[36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[36]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b37  (
    .clk(clk),
    .d(addr_ex[37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[37]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b38  (
    .clk(clk),
    .d(addr_ex[38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[38]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b39  (
    .clk(clk),
    .d(addr_ex[39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[39]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b4  (
    .clk(clk),
    .d(addr_ex[4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[4]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b40  (
    .clk(clk),
    .d(addr_ex[40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[40]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b41  (
    .clk(clk),
    .d(addr_ex[41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[41]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b42  (
    .clk(clk),
    .d(addr_ex[42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[42]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b43  (
    .clk(clk),
    .d(addr_ex[43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[43]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b44  (
    .clk(clk),
    .d(addr_ex[44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[44]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b45  (
    .clk(clk),
    .d(addr_ex[45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[45]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b46  (
    .clk(clk),
    .d(addr_ex[46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[46]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b47  (
    .clk(clk),
    .d(addr_ex[47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[47]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b48  (
    .clk(clk),
    .d(addr_ex[48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[48]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b49  (
    .clk(clk),
    .d(addr_ex[49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[49]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b5  (
    .clk(clk),
    .d(addr_ex[5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[5]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b50  (
    .clk(clk),
    .d(addr_ex[50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[50]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b51  (
    .clk(clk),
    .d(addr_ex[51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[51]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b52  (
    .clk(clk),
    .d(addr_ex[52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[52]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b53  (
    .clk(clk),
    .d(addr_ex[53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[53]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b54  (
    .clk(clk),
    .d(addr_ex[54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[54]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b55  (
    .clk(clk),
    .d(addr_ex[55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[55]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b56  (
    .clk(clk),
    .d(addr_ex[56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[56]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b57  (
    .clk(clk),
    .d(addr_ex[57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[57]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b58  (
    .clk(clk),
    .d(addr_ex[58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[58]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b59  (
    .clk(clk),
    .d(addr_ex[59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[59]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b6  (
    .clk(clk),
    .d(addr_ex[6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[6]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b60  (
    .clk(clk),
    .d(addr_ex[60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[60]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b61  (
    .clk(clk),
    .d(addr_ex[61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[61]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b62  (
    .clk(clk),
    .d(addr_ex[62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[62]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b63  (
    .clk(clk),
    .d(addr_ex[63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[63]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b7  (
    .clk(clk),
    .d(addr_ex[7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[7]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b8  (
    .clk(clk),
    .d(addr_ex[8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[8]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg3_b9  (
    .clk(clk),
    .d(addr_ex[9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(new_pc[9]));  // ../../RTL/CPU/EX/exu.v(342)
  reg_sr_as_w1 \exu/reg4_b0  (
    .clk(clk),
    .d(ex_ins_pc[0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[0]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b1  (
    .clk(clk),
    .d(ex_ins_pc[1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[1]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b10  (
    .clk(clk),
    .d(ex_ins_pc[10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[10]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b11  (
    .clk(clk),
    .d(ex_ins_pc[11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[11]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b12  (
    .clk(clk),
    .d(ex_ins_pc[12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[12]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b13  (
    .clk(clk),
    .d(ex_ins_pc[13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[13]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b14  (
    .clk(clk),
    .d(ex_ins_pc[14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[14]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b15  (
    .clk(clk),
    .d(ex_ins_pc[15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[15]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b16  (
    .clk(clk),
    .d(ex_ins_pc[16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[16]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b17  (
    .clk(clk),
    .d(ex_ins_pc[17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[17]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b18  (
    .clk(clk),
    .d(ex_ins_pc[18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[18]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b19  (
    .clk(clk),
    .d(ex_ins_pc[19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[19]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b2  (
    .clk(clk),
    .d(ex_ins_pc[2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[2]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b20  (
    .clk(clk),
    .d(ex_ins_pc[20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[20]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b21  (
    .clk(clk),
    .d(ex_ins_pc[21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[21]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b22  (
    .clk(clk),
    .d(ex_ins_pc[22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[22]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b23  (
    .clk(clk),
    .d(ex_ins_pc[23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[23]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b24  (
    .clk(clk),
    .d(ex_ins_pc[24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[24]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b25  (
    .clk(clk),
    .d(ex_ins_pc[25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[25]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b26  (
    .clk(clk),
    .d(ex_ins_pc[26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[26]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b27  (
    .clk(clk),
    .d(ex_ins_pc[27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[27]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b28  (
    .clk(clk),
    .d(ex_ins_pc[28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[28]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b29  (
    .clk(clk),
    .d(ex_ins_pc[29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[29]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b3  (
    .clk(clk),
    .d(ex_ins_pc[3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[3]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b30  (
    .clk(clk),
    .d(ex_ins_pc[30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[30]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b31  (
    .clk(clk),
    .d(ex_ins_pc[31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[31]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b32  (
    .clk(clk),
    .d(ex_ins_pc[32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[32]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b33  (
    .clk(clk),
    .d(ex_ins_pc[33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[33]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b34  (
    .clk(clk),
    .d(ex_ins_pc[34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[34]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b35  (
    .clk(clk),
    .d(ex_ins_pc[35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[35]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b36  (
    .clk(clk),
    .d(ex_ins_pc[36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[36]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b37  (
    .clk(clk),
    .d(ex_ins_pc[37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[37]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b38  (
    .clk(clk),
    .d(ex_ins_pc[38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[38]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b39  (
    .clk(clk),
    .d(ex_ins_pc[39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[39]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b4  (
    .clk(clk),
    .d(ex_ins_pc[4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[4]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b40  (
    .clk(clk),
    .d(ex_ins_pc[40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[40]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b41  (
    .clk(clk),
    .d(ex_ins_pc[41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[41]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b42  (
    .clk(clk),
    .d(ex_ins_pc[42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[42]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b43  (
    .clk(clk),
    .d(ex_ins_pc[43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[43]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b44  (
    .clk(clk),
    .d(ex_ins_pc[44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[44]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b45  (
    .clk(clk),
    .d(ex_ins_pc[45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[45]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b46  (
    .clk(clk),
    .d(ex_ins_pc[46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[46]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b47  (
    .clk(clk),
    .d(ex_ins_pc[47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[47]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b48  (
    .clk(clk),
    .d(ex_ins_pc[48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[48]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b49  (
    .clk(clk),
    .d(ex_ins_pc[49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[49]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b5  (
    .clk(clk),
    .d(ex_ins_pc[5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[5]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b50  (
    .clk(clk),
    .d(ex_ins_pc[50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[50]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b51  (
    .clk(clk),
    .d(ex_ins_pc[51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[51]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b52  (
    .clk(clk),
    .d(ex_ins_pc[52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[52]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b53  (
    .clk(clk),
    .d(ex_ins_pc[53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[53]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b54  (
    .clk(clk),
    .d(ex_ins_pc[54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[54]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b55  (
    .clk(clk),
    .d(ex_ins_pc[55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[55]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b56  (
    .clk(clk),
    .d(ex_ins_pc[56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[56]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b57  (
    .clk(clk),
    .d(ex_ins_pc[57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[57]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b58  (
    .clk(clk),
    .d(ex_ins_pc[58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[58]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b59  (
    .clk(clk),
    .d(ex_ins_pc[59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[59]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b6  (
    .clk(clk),
    .d(ex_ins_pc[6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[6]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b60  (
    .clk(clk),
    .d(ex_ins_pc[60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[60]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b61  (
    .clk(clk),
    .d(ex_ins_pc[61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[61]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b62  (
    .clk(clk),
    .d(ex_ins_pc[62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[62]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b63  (
    .clk(clk),
    .d(ex_ins_pc[63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[63]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b7  (
    .clk(clk),
    .d(ex_ins_pc[7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[7]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b8  (
    .clk(clk),
    .d(ex_ins_pc[8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[8]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg4_b9  (
    .clk(clk),
    .d(ex_ins_pc[9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_ins_pc[9]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b0  (
    .clk(clk),
    .d(\exu/n71 [0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[0]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b1  (
    .clk(clk),
    .d(\exu/n71 [1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[1]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b10  (
    .clk(clk),
    .d(\exu/n71 [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[10]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b11  (
    .clk(clk),
    .d(\exu/n71 [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[11]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b12  (
    .clk(clk),
    .d(\exu/n71 [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[12]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b13  (
    .clk(clk),
    .d(\exu/n71 [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[13]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b14  (
    .clk(clk),
    .d(\exu/n71 [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[14]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b15  (
    .clk(clk),
    .d(\exu/n71 [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[15]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b16  (
    .clk(clk),
    .d(\exu/n71 [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[16]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b17  (
    .clk(clk),
    .d(\exu/n71 [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[17]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b18  (
    .clk(clk),
    .d(\exu/n71 [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[18]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b19  (
    .clk(clk),
    .d(\exu/n71 [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[19]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b2  (
    .clk(clk),
    .d(\exu/n71 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[2]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b20  (
    .clk(clk),
    .d(\exu/n71 [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[20]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b21  (
    .clk(clk),
    .d(\exu/n71 [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[21]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b22  (
    .clk(clk),
    .d(\exu/n71 [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[22]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b23  (
    .clk(clk),
    .d(\exu/n71 [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[23]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b24  (
    .clk(clk),
    .d(\exu/n71 [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[24]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b25  (
    .clk(clk),
    .d(\exu/n71 [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[25]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b26  (
    .clk(clk),
    .d(\exu/n71 [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[26]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b27  (
    .clk(clk),
    .d(\exu/n71 [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[27]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b28  (
    .clk(clk),
    .d(\exu/n71 [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[28]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b29  (
    .clk(clk),
    .d(\exu/n71 [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[29]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b3  (
    .clk(clk),
    .d(\exu/n71 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[3]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b30  (
    .clk(clk),
    .d(\exu/n71 [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[30]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b31  (
    .clk(clk),
    .d(\exu/n71 [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[31]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b32  (
    .clk(clk),
    .d(\exu/n71 [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[32]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b33  (
    .clk(clk),
    .d(\exu/n71 [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[33]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b34  (
    .clk(clk),
    .d(\exu/n71 [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[34]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b35  (
    .clk(clk),
    .d(\exu/n71 [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[35]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b36  (
    .clk(clk),
    .d(\exu/n71 [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[36]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b37  (
    .clk(clk),
    .d(\exu/n71 [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[37]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b38  (
    .clk(clk),
    .d(\exu/n71 [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[38]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b39  (
    .clk(clk),
    .d(\exu/n71 [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[39]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b4  (
    .clk(clk),
    .d(\exu/n71 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[4]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b40  (
    .clk(clk),
    .d(\exu/n71 [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[40]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b41  (
    .clk(clk),
    .d(\exu/n71 [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[41]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b42  (
    .clk(clk),
    .d(\exu/n71 [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[42]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b43  (
    .clk(clk),
    .d(\exu/n71 [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[43]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b44  (
    .clk(clk),
    .d(\exu/n71 [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[44]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b45  (
    .clk(clk),
    .d(\exu/n71 [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[45]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b46  (
    .clk(clk),
    .d(\exu/n71 [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[46]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b47  (
    .clk(clk),
    .d(\exu/n71 [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[47]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b48  (
    .clk(clk),
    .d(\exu/n71 [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[48]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b49  (
    .clk(clk),
    .d(\exu/n71 [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[49]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b5  (
    .clk(clk),
    .d(\exu/n71 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[5]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b50  (
    .clk(clk),
    .d(\exu/n71 [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[50]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b51  (
    .clk(clk),
    .d(\exu/n71 [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[51]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b52  (
    .clk(clk),
    .d(\exu/n71 [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[52]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b53  (
    .clk(clk),
    .d(\exu/n71 [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[53]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b54  (
    .clk(clk),
    .d(\exu/n71 [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[54]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b55  (
    .clk(clk),
    .d(\exu/n71 [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[55]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b56  (
    .clk(clk),
    .d(\exu/n71 [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[56]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b57  (
    .clk(clk),
    .d(\exu/n71 [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[57]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b58  (
    .clk(clk),
    .d(\exu/n71 [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[58]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b59  (
    .clk(clk),
    .d(\exu/n71 [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[59]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b6  (
    .clk(clk),
    .d(\exu/n71 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[6]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b60  (
    .clk(clk),
    .d(\exu/n71 [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[60]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b61  (
    .clk(clk),
    .d(\exu/n71 [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[61]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b62  (
    .clk(clk),
    .d(\exu/n71 [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[62]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b63  (
    .clk(clk),
    .d(\exu/n71 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[63]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b7  (
    .clk(clk),
    .d(\exu/n71 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[7]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b8  (
    .clk(clk),
    .d(\exu/n71 [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[8]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg5_b9  (
    .clk(clk),
    .d(\exu/n71 [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_exc_code[9]));  // ../../RTL/CPU/EX/exu.v(358)
  reg_sr_as_w1 \exu/reg6_b0  (
    .clk(clk),
    .d(ex_csr_index[0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[0]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b1  (
    .clk(clk),
    .d(ex_csr_index[1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[1]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b10  (
    .clk(clk),
    .d(ex_csr_index[10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[10]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b11  (
    .clk(clk),
    .d(ex_csr_index[11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[11]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b2  (
    .clk(clk),
    .d(ex_csr_index[2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[2]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b3  (
    .clk(clk),
    .d(ex_csr_index[3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[3]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b4  (
    .clk(clk),
    .d(ex_csr_index[4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[4]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b5  (
    .clk(clk),
    .d(ex_csr_index[5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[5]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b6  (
    .clk(clk),
    .d(ex_csr_index[6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[6]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b7  (
    .clk(clk),
    .d(ex_csr_index[7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[7]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b8  (
    .clk(clk),
    .d(ex_csr_index[8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[8]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg6_b9  (
    .clk(clk),
    .d(ex_csr_index[9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(csr_index[9]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg7_b0  (
    .clk(clk),
    .d(ex_rd_index[0]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_rd_index[0]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg7_b1  (
    .clk(clk),
    .d(ex_rd_index[1]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_rd_index[1]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg7_b2  (
    .clk(clk),
    .d(ex_rd_index[2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_rd_index[2]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg7_b3  (
    .clk(clk),
    .d(ex_rd_index[3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_rd_index[3]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg7_b4  (
    .clk(clk),
    .d(ex_rd_index[4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(wb_rd_index[4]));  // ../../RTL/CPU/EX/exu.v(383)
  reg_sr_as_w1 \exu/reg8_b0  (
    .clk(clk),
    .d(\exu/n45 [0]),
    .en(~ex_nop),
    .reset(rst),
    .set(1'b0),
    .q(\exu/main_state [0]));  // ../../RTL/CPU/EX/exu.v(268)
  reg_sr_as_w1 \exu/reg8_b1  (
    .clk(clk),
    .d(\exu/n45 [1]),
    .en(~ex_nop),
    .reset(rst),
    .set(1'b0),
    .q(\exu/main_state [1]));  // ../../RTL/CPU/EX/exu.v(268)
  reg_sr_as_w1 \exu/reg8_b2  (
    .clk(clk),
    .d(\exu/n45 [2]),
    .en(~ex_nop),
    .reset(rst),
    .set(1'b0),
    .q(\exu/main_state [2]));  // ../../RTL/CPU/EX/exu.v(268)
  reg_sr_as_w1 \exu/reg8_b3  (
    .clk(clk),
    .d(\exu/n45 [3]),
    .en(~ex_nop),
    .reset(rst),
    .set(1'b0),
    .q(\exu/main_state [3]));  // ../../RTL/CPU/EX/exu.v(268)
  reg_sr_as_w1 \exu/s_ret_reg  (
    .clk(clk),
    .d(ex_s_ret),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_s_ret));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/st_acc_fault_reg  (
    .clk(clk),
    .d(\exu/n90 ),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_st_acc_fault));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/st_addr_mis_reg  (
    .clk(clk),
    .d(\exu/n88 ),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_st_addr_mis));  // ../../RTL/CPU/EX/exu.v(448)
  reg_sr_as_w1 \exu/st_page_fault_reg  (
    .clk(clk),
    .d(\exu/n92 ),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_st_page_fault));  // ../../RTL/CPU/EX/exu.v(448)
  add_pu8_mu8_o8 \exu/sub0  (
    .i0(\exu/shift_count ),
    .i1(8'b00000001),
    .o(\exu/n50 ));  // ../../RTL/CPU/EX/exu.v(288)
  and \exu/u10  (\exu/load_addr_mis , \exu/n0 , \exu/n8 );  // ../../RTL/CPU/EX/exu.v(211)
  or \exu/u100  (\exu/n60 , \exu/c_load_1 , \exu/c_amo_mem01 );  // ../../RTL/CPU/EX/exu.v(324)
  or \exu/u107  (\exu/n86 , rst, ex_nop);  // ../../RTL/CPU/EX/exu.v(388)
  and \exu/u108  (\exu/n87 , \exu/c_amo_mem0 , \exu/load_addr_mis );  // ../../RTL/CPU/EX/exu.v(435)
  or \exu/u109  (\exu/n88 , \exu/n87 , \exu/store_addr_mis );  // ../../RTL/CPU/EX/exu.v(435)
  and \exu/u110  (\exu/n89 , \exu/c_amo_mem0 , load_acc_fault);  // ../../RTL/CPU/EX/exu.v(437)
  or \exu/u111  (\exu/n90 , \exu/n89 , store_acc_fault);  // ../../RTL/CPU/EX/exu.v(437)
  and \exu/u112  (\exu/n91 , \exu/c_amo_mem0 , load_page_fault);  // ../../RTL/CPU/EX/exu.v(439)
  or \exu/u113  (\exu/n92 , \exu/n91 , store_page_fault);  // ../../RTL/CPU/EX/exu.v(439)
  or \exu/u114  (\exu/n93 , ex_ready, ex_more_exception);  // ../../RTL/CPU/EX/exu.v(441)
  or \exu/u115  (\exu/n94 , \exu/n93 , \exu/exception_id );  // ../../RTL/CPU/EX/exu.v(441)
  and \exu/u116  (\exu/n95 , ex_valid, \exu/n94 );  // ../../RTL/CPU/EX/exu.v(441)
  or \exu/u153  (\exu/n132 , load, store);  // ../../RTL/CPU/EX/exu.v(451)
  or \exu/u154  (\exu/n133 , \exu/n132 , amo);  // ../../RTL/CPU/EX/exu.v(451)
  or \exu/u155  (\exu/n134 , \exu/n133 , cache_flush);  // ../../RTL/CPU/EX/exu.v(451)
  or \exu/u156  (\exu/n135 , \exu/n134 , cache_reset);  // ../../RTL/CPU/EX/exu.v(451)
  or \exu/u157  (\exu/n136 , \exu/n135 , shift_l);  // ../../RTL/CPU/EX/exu.v(451)
  or \exu/u158  (\exu/n137 , \exu/n136 , shift_r);  // ../../RTL/CPU/EX/exu.v(451)
  not \exu/u159  (\exu/n138 , \exu/n137 );  // ../../RTL/CPU/EX/exu.v(451)
  and \exu/u160  (\exu/n139 , load, \exu/load_ready );  // ../../RTL/CPU/EX/exu.v(452)
  or \exu/u161  (\exu/n140 , \exu/n138 , \exu/n139 );  // ../../RTL/CPU/EX/exu.v(452)
  and \exu/u162  (\exu/n141 , store, \exu/store_ready );  // ../../RTL/CPU/EX/exu.v(452)
  or \exu/u163  (\exu/n142 , \exu/n140 , \exu/n141 );  // ../../RTL/CPU/EX/exu.v(452)
  and \exu/u164  (\exu/n143 , amo, \exu/amo_ready );  // ../../RTL/CPU/EX/exu.v(452)
  or \exu/u165  (\exu/n144 , \exu/n142 , \exu/n143 );  // ../../RTL/CPU/EX/exu.v(452)
  and \exu/u167  (\exu/n145 , \exu/n21 , \exu/fence_ready );  // ../../RTL/CPU/EX/exu.v(453)
  or \exu/u168  (\exu/n146 , \exu/n144 , \exu/n145 );  // ../../RTL/CPU/EX/exu.v(453)
  and \exu/u170  (\exu/n147 , \exu/n20 , \exu/shift_multi_ready );  // ../../RTL/CPU/EX/exu.v(453)
  or \exu/u171  (ex_ready, \exu/n146 , \exu/n147 );  // ../../RTL/CPU/EX/exu.v(453)
  and \exu/u172  (unpage, mprv, \exu/n148 );  // ../../RTL/CPU/EX/exu.v(506)
  and \exu/u174  (cache_flush_biu, cache_flush, \exu/c_fence );  // ../../RTL/CPU/EX/exu.v(512)
  and \exu/u177  (read, load, \exu/n59 );  // ../../RTL/CPU/EX/exu.v(514)
  or \exu/u178  (\exu/n149 , \exu/c_amo_mem1 , \exu/c_store );  // ../../RTL/CPU/EX/exu.v(515)
  and \exu/u179  (write, store, \exu/n149 );  // ../../RTL/CPU/EX/exu.v(515)
  and \exu/u19  (\exu/store_addr_mis , store, \exu/n8 );  // ../../RTL/CPU/EX/exu.v(212)
  and \exu/u24  (\exu/shift_ready , \exu/c_shift , \exu/n9 );  // ../../RTL/CPU/EX/exu.v(215)
  and \exu/u25  (\exu/n10 , \exu/c_load , uncache_data_rdy);  // ../../RTL/CPU/EX/exu.v(217)
  or \exu/u26  (\exu/load_ready , \exu/n10 , \exu/c_load_1 );  // ../../RTL/CPU/EX/exu.v(217)
  and \exu/u27  (\exu/store_ready , \exu/c_store , cache_ready_ex);  // ../../RTL/CPU/EX/exu.v(218)
  and \exu/u28  (\exu/fence_ready , \exu/c_fence , cache_ready_ex);  // ../../RTL/CPU/EX/exu.v(219)
  and \exu/u29  (\exu/amo_ready , \exu/c_amo_mem1 , cache_ready_ex);  // ../../RTL/CPU/EX/exu.v(220)
  and \exu/u30  (\exu/shift_multi_ready , \exu/c_shift , \exu/shift_ready );  // ../../RTL/CPU/EX/exu.v(221)
  or \exu/u31  (\exu/n11 , ex_ins_acc_fault, ex_ins_addr_mis);  // ../../RTL/CPU/EX/exu.v(223)
  or \exu/u32  (\exu/n12 , \exu/n11 , ex_ins_page_fault);  // ../../RTL/CPU/EX/exu.v(223)
  or \exu/u33  (\exu/exception_id , \exu/n12 , ex_ill_ins);  // ../../RTL/CPU/EX/exu.v(223)
  or \exu/u34  (\exu/n13 , load_acc_fault, load_page_fault);  // ../../RTL/CPU/EX/exu.v(224)
  or \exu/u35  (\exu/n14 , \exu/n13 , store_acc_fault);  // ../../RTL/CPU/EX/exu.v(224)
  or \exu/u36  (\exu/n15 , \exu/n14 , store_page_fault);  // ../../RTL/CPU/EX/exu.v(224)
  or \exu/u37  (\exu/n16 , \exu/n15 , \exu/load_addr_mis );  // ../../RTL/CPU/EX/exu.v(224)
  or \exu/u38  (ex_more_exception, \exu/n16 , \exu/store_addr_mis );  // ../../RTL/CPU/EX/exu.v(224)
  not \exu/u39  (\exu/n17 , \exu/exception_id );  // ../../RTL/CPU/EX/exu.v(235)
  or \exu/u4  (\exu/n0 , amo, load);  // ../../RTL/CPU/EX/exu.v(211)
  and \exu/u40  (\exu/n18 , ex_valid, \exu/n17 );  // ../../RTL/CPU/EX/exu.v(235)
  and \exu/u41  (\exu/n19 , \exu/n18 , \exu/c_stb );  // ../../RTL/CPU/EX/exu.v(235)
  or \exu/u42  (\exu/n20 , shift_l, shift_r);  // ../../RTL/CPU/EX/exu.v(238)
  or \exu/u43  (\exu/n21 , cache_flush, cache_reset);  // ../../RTL/CPU/EX/exu.v(240)
  or \exu/u44  (\exu/n28 , cache_ready_ex, uncache_data_rdy);  // ../../RTL/CPU/EX/exu.v(247)
  not \exu/u47  (\exu/n31 , \exu/shift_ready );  // ../../RTL/CPU/EX/exu.v(250)
  and \exu/u5  (\exu/n2 , ex_size[1], \biu/cache_ctrl_logic/n197 );  // ../../RTL/CPU/EX/exu.v(211)
  not \exu/u58  (\exu/n29 [2], \exu/n28 );  // ../../RTL/CPU/EX/exu.v(247)
  and \exu/u6  (\exu/n4 , ex_size[2], \exu/n3 );  // ../../RTL/CPU/EX/exu.v(211)
  and \exu/u62  (\exu/n48 , \exu/c_stb , ex_valid);  // ../../RTL/CPU/EX/exu.v(284)
  and \exu/u64  (\exu/n49 , \exu/n48 , \exu/n20 );  // ../../RTL/CPU/EX/exu.v(284)
  or \exu/u7  (\exu/n5 , \exu/n2 , \exu/n4 );  // ../../RTL/CPU/EX/exu.v(211)
  and \exu/u8  (\exu/n7 , ex_size[3], \exu/n6 );  // ../../RTL/CPU/EX/exu.v(211)
  or \exu/u9  (\exu/n8 , \exu/n5 , \exu/n7 );  // ../../RTL/CPU/EX/exu.v(211)
  or \exu/u99  (\exu/n59 , \exu/c_load , \exu/c_amo_mem0 );  // ../../RTL/CPU/EX/exu.v(321)
  reg_sr_as_w1 \exu/valid_reg  (
    .clk(clk),
    .d(\exu/n95 ),
    .en(1'b1),
    .reset(\exu/n86 ),
    .set(1'b0),
    .q(wb_valid));  // ../../RTL/CPU/EX/exu.v(448)
  not id_hold_inv (id_hold_neg, id_hold);
  not id_nop_inv (id_nop_neg, id_nop);
  not ins_acc_fault_inv (ins_acc_fault_neg, ins_acc_fault);
  reg_sr_as_w1 \ins_dec/amo_reg  (
    .clk(clk),
    .d(\ins_dec/op_amo ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(amo));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/and_clr_reg  (
    .clk(clk),
    .d(\ins_dec/n71 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(and_clr));  // ../../RTL/CPU/ID/ins_dec.v(674)
  reg_sr_as_w1 \ins_dec/cache_flush_reg  (
    .clk(clk),
    .d(\ins_dec/ins_fence ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(cache_flush));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/cache_reset_reg  (
    .clk(clk),
    .d(\ins_dec/n225 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(cache_reset));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/csr_write_reg  (
    .clk(clk),
    .d(\ins_dec/n239 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_write));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/ebreak_reg  (
    .clk(clk),
    .d(\ins_dec/ins_ebreak ),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ebreak));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/ecall_reg  (
    .clk(clk),
    .d(\ins_dec/ins_ecall ),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ecall));  // ../../RTL/CPU/ID/ins_dec.v(830)
  eq_w7 \ins_dec/eq0  (
    .i0(id_ins[6:0]),
    .i1(7'b0001111),
    .o(id_system));  // ../../RTL/CPU/ID/ins_dec.v(346)
  eq_w7 \ins_dec/eq1  (
    .i0(id_ins[6:0]),
    .i1(7'b0010011),
    .o(\ins_dec/op_imm ));  // ../../RTL/CPU/ID/ins_dec.v(347)
  eq_w7 \ins_dec/eq10  (
    .i0(id_ins[6:0]),
    .i1(7'b0110011),
    .o(\ins_dec/op_reg ));  // ../../RTL/CPU/ID/ins_dec.v(356)
  eq_w7 \ins_dec/eq11  (
    .i0(id_ins[6:0]),
    .i1(7'b0111011),
    .o(\ins_dec/op_32_reg ));  // ../../RTL/CPU/ID/ins_dec.v(357)
  eq_w7 \ins_dec/eq12  (
    .i0(id_ins[6:0]),
    .i1(7'b0101111),
    .o(\ins_dec/op_amo ));  // ../../RTL/CPU/ID/ins_dec.v(358)
  eq_w3 \ins_dec/eq13  (
    .i0(id_ins[14:12]),
    .i1(3'b000),
    .o(\ins_dec/funct3_0 ));  // ../../RTL/CPU/ID/ins_dec.v(363)
  eq_w3 \ins_dec/eq14  (
    .i0(id_ins[14:12]),
    .i1(3'b001),
    .o(\ins_dec/funct3_1 ));  // ../../RTL/CPU/ID/ins_dec.v(364)
  eq_w3 \ins_dec/eq15  (
    .i0(id_ins[14:12]),
    .i1(3'b010),
    .o(\ins_dec/funct3_2 ));  // ../../RTL/CPU/ID/ins_dec.v(365)
  eq_w3 \ins_dec/eq16  (
    .i0(id_ins[14:12]),
    .i1(3'b011),
    .o(\ins_dec/funct3_3 ));  // ../../RTL/CPU/ID/ins_dec.v(366)
  eq_w3 \ins_dec/eq17  (
    .i0(id_ins[14:12]),
    .i1(3'b100),
    .o(\ins_dec/funct3_4 ));  // ../../RTL/CPU/ID/ins_dec.v(367)
  eq_w3 \ins_dec/eq18  (
    .i0(id_ins[14:12]),
    .i1(3'b101),
    .o(\ins_dec/funct3_5 ));  // ../../RTL/CPU/ID/ins_dec.v(368)
  eq_w3 \ins_dec/eq19  (
    .i0(id_ins[14:12]),
    .i1(3'b110),
    .o(\ins_dec/funct3_6 ));  // ../../RTL/CPU/ID/ins_dec.v(369)
  eq_w7 \ins_dec/eq2  (
    .i0(id_ins[6:0]),
    .i1(7'b0011011),
    .o(\ins_dec/op_32_imm ));  // ../../RTL/CPU/ID/ins_dec.v(348)
  eq_w3 \ins_dec/eq20  (
    .i0(id_ins[14:12]),
    .i1(3'b111),
    .o(\ins_dec/funct3_7 ));  // ../../RTL/CPU/ID/ins_dec.v(370)
  eq_w5 \ins_dec/eq21  (
    .i0(id_ins[31:27]),
    .i1(5'b00000),
    .o(\ins_dec/funct5_0 ));  // ../../RTL/CPU/ID/ins_dec.v(372)
  eq_w5 \ins_dec/eq22  (
    .i0(id_ins[31:27]),
    .i1(5'b00001),
    .o(\ins_dec/funct5_1 ));  // ../../RTL/CPU/ID/ins_dec.v(373)
  eq_w5 \ins_dec/eq23  (
    .i0(id_ins[31:27]),
    .i1(5'b00010),
    .o(\ins_dec/funct5_2 ));  // ../../RTL/CPU/ID/ins_dec.v(374)
  eq_w5 \ins_dec/eq24  (
    .i0(id_ins[31:27]),
    .i1(5'b00011),
    .o(\ins_dec/funct5_3 ));  // ../../RTL/CPU/ID/ins_dec.v(375)
  eq_w5 \ins_dec/eq25  (
    .i0(id_ins[31:27]),
    .i1(5'b00100),
    .o(\ins_dec/funct5_4 ));  // ../../RTL/CPU/ID/ins_dec.v(376)
  eq_w5 \ins_dec/eq26  (
    .i0(id_ins[31:27]),
    .i1(5'b01000),
    .o(\ins_dec/funct5_8 ));  // ../../RTL/CPU/ID/ins_dec.v(380)
  eq_w5 \ins_dec/eq27  (
    .i0(id_ins[31:27]),
    .i1(5'b01100),
    .o(\ins_dec/funct5_12 ));  // ../../RTL/CPU/ID/ins_dec.v(384)
  eq_w5 \ins_dec/eq28  (
    .i0(id_ins[31:27]),
    .i1(5'b10000),
    .o(\ins_dec/funct5_16 ));  // ../../RTL/CPU/ID/ins_dec.v(388)
  eq_w5 \ins_dec/eq29  (
    .i0(id_ins[31:27]),
    .i1(5'b10100),
    .o(\ins_dec/funct5_20 ));  // ../../RTL/CPU/ID/ins_dec.v(392)
  eq_w7 \ins_dec/eq3  (
    .i0(id_ins[6:0]),
    .i1(7'b0110111),
    .o(\ins_dec/op_lui ));  // ../../RTL/CPU/ID/ins_dec.v(349)
  eq_w5 \ins_dec/eq30  (
    .i0(id_ins[31:27]),
    .i1(5'b11000),
    .o(\ins_dec/funct5_24 ));  // ../../RTL/CPU/ID/ins_dec.v(396)
  eq_w5 \ins_dec/eq31  (
    .i0(id_ins[31:27]),
    .i1(5'b11100),
    .o(\ins_dec/funct5_28 ));  // ../../RTL/CPU/ID/ins_dec.v(400)
  eq_w6 \ins_dec/eq32  (
    .i0(id_ins[31:26]),
    .i1(6'b000000),
    .o(\ins_dec/funct6_0 ));  // ../../RTL/CPU/ID/ins_dec.v(405)
  eq_w6 \ins_dec/eq33  (
    .i0(id_ins[31:26]),
    .i1(6'b010000),
    .o(\ins_dec/funct6_16 ));  // ../../RTL/CPU/ID/ins_dec.v(406)
  eq_w7 \ins_dec/eq34  (
    .i0(id_ins[31:25]),
    .i1(7'b0000000),
    .o(\ins_dec/funct7_0 ));  // ../../RTL/CPU/ID/ins_dec.v(408)
  eq_w7 \ins_dec/eq35  (
    .i0(id_ins[31:25]),
    .i1(7'b0001000),
    .o(\ins_dec/funct7_8 ));  // ../../RTL/CPU/ID/ins_dec.v(409)
  eq_w7 \ins_dec/eq36  (
    .i0(id_ins[31:25]),
    .i1(7'b0001001),
    .o(\ins_dec/funct7_9 ));  // ../../RTL/CPU/ID/ins_dec.v(410)
  eq_w7 \ins_dec/eq37  (
    .i0(id_ins[31:25]),
    .i1(7'b0011000),
    .o(\ins_dec/funct7_24 ));  // ../../RTL/CPU/ID/ins_dec.v(411)
  eq_w7 \ins_dec/eq38  (
    .i0(id_ins[31:25]),
    .i1(7'b0101111),
    .o(\ins_dec/funct7_32 ));  // ../../RTL/CPU/ID/ins_dec.v(412)
  eq_w12 \ins_dec/eq39  (
    .i0(id_ins[31:20]),
    .i1(12'b000000000000),
    .o(\ins_dec/funct12_0 ));  // ../../RTL/CPU/ID/ins_dec.v(415)
  eq_w7 \ins_dec/eq4  (
    .i0(id_ins[6:0]),
    .i1(7'b0010111),
    .o(\ins_dec/op_auipc ));  // ../../RTL/CPU/ID/ins_dec.v(350)
  eq_w12 \ins_dec/eq40  (
    .i0(id_ins[31:20]),
    .i1(12'b000000000001),
    .o(\ins_dec/funct12_1 ));  // ../../RTL/CPU/ID/ins_dec.v(416)
  eq_w5 \ins_dec/eq41  (
    .i0(id_rs2_index),
    .i1(5'b00010),
    .o(\ins_dec/n44 ));  // ../../RTL/CPU/ID/ins_dec.v(502)
  eq_w2 \ins_dec/eq45  (
    .i0(id_ins[29:28]),
    .i1(2'b00),
    .o(\ins_dec/n80 ));  // ../../RTL/CPU/ID/ins_dec.v(550)
  eq_w7 \ins_dec/eq5  (
    .i0(id_ins[6:0]),
    .i1(7'b1101111),
    .o(\ins_dec/op_jal ));  // ../../RTL/CPU/ID/ins_dec.v(351)
  eq_w7 \ins_dec/eq6  (
    .i0(id_ins[6:0]),
    .i1(7'b1100111),
    .o(\ins_dec/op_jalr ));  // ../../RTL/CPU/ID/ins_dec.v(352)
  eq_w7 \ins_dec/eq7  (
    .i0(id_ins[6:0]),
    .i1(7'b1100011),
    .o(\ins_dec/op_branch ));  // ../../RTL/CPU/ID/ins_dec.v(353)
  eq_w7 \ins_dec/eq8  (
    .i0(id_ins[6:0]),
    .i1(7'b0000011),
    .o(\ins_dec/op_load ));  // ../../RTL/CPU/ID/ins_dec.v(354)
  eq_w7 \ins_dec/eq9  (
    .i0(id_ins[6:0]),
    .i1(7'b0100011),
    .o(\ins_dec/op_store ));  // ../../RTL/CPU/ID/ins_dec.v(355)
  reg_sr_as_w1 \ins_dec/gpr_write_reg  (
    .clk(clk),
    .d(\ins_dec/dec_gpr_write ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_gpr_write));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/id_jmp_reg  (
    .clk(clk),
    .d(\ins_dec/n302 ),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_jmp));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/id_system_reg  (
    .clk(clk),
    .d(id_system),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_system));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/ill_ins_reg  (
    .clk(clk),
    .d(id_ill_ins),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ill_ins));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/ins_acc_fault_reg  (
    .clk(clk),
    .d(id_ins_acc_fault),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_acc_fault));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/ins_addr_mis_reg  (
    .clk(clk),
    .d(id_ins_addr_mis),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_addr_mis));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/ins_page_fault_reg  (
    .clk(clk),
    .d(id_ins_page_fault),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_page_fault));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/int_acc_reg  (
    .clk(clk),
    .d(id_int_acc),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_int_acc));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/jmp_reg  (
    .clk(clk),
    .d(\ins_dec/n59 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(jmp));  // ../../RTL/CPU/ID/ins_dec.v(674)
  reg_sr_as_w1 \ins_dec/load_reg  (
    .clk(clk),
    .d(\ins_dec/op_load ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(load));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/m_ret_reg  (
    .clk(clk),
    .d(\ins_dec/n304 ),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_m_ret));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/mem_csr_data_add_reg  (
    .clk(clk),
    .d(\ins_dec/n146 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_add));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_and_reg  (
    .clk(clk),
    .d(\ins_dec/n148 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_and));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_ds2_reg  (
    .clk(clk),
    .d(\ins_dec/n145 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_ds2));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_max_reg  (
    .clk(clk),
    .d(\ins_dec/n155 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_max));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_min_reg  (
    .clk(clk),
    .d(\ins_dec/n158 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_min));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_or_reg  (
    .clk(clk),
    .d(\ins_dec/n151 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_or));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/mem_csr_data_xor_reg  (
    .clk(clk),
    .d(\ins_dec/n152 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(mem_csr_data_xor));  // ../../RTL/CPU/ID/ins_dec.v(636)
  binary_mux_s1_w1 \ins_dec/mux0_b0  (
    .i0(rs2_data[0]),
    .i1(id_ins[15]),
    .sel(\ins_dec/n57 ),
    .o(\ins_dec/n58 [0]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  binary_mux_s1_w1 \ins_dec/mux0_b1  (
    .i0(rs2_data[1]),
    .i1(id_ins[16]),
    .sel(\ins_dec/n57 ),
    .o(\ins_dec/n58 [1]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  binary_mux_s1_w1 \ins_dec/mux0_b2  (
    .i0(rs2_data[2]),
    .i1(id_ins[17]),
    .sel(\ins_dec/n57 ),
    .o(\ins_dec/n58 [2]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  binary_mux_s1_w1 \ins_dec/mux0_b3  (
    .i0(rs2_data[3]),
    .i1(id_ins[18]),
    .sel(\ins_dec/n57 ),
    .o(\ins_dec/n58 [3]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  binary_mux_s1_w1 \ins_dec/mux0_b4  (
    .i0(rs2_data[4]),
    .i1(id_ins[19]),
    .sel(\ins_dec/n57 ),
    .o(\ins_dec/n58 [4]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  binary_mux_s1_w1 \ins_dec/mux0_b5  (
    .i0(rs2_data[5]),
    .i1(id_ins[20]),
    .sel(\ins_dec/n57 ),
    .o(\ins_dec/n58 [5]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  and \ins_dec/mux13_b0_sel_is_0  (\ins_dec/mux13_b0_sel_is_0_o , \ins_dec/n107_neg , id_hold_neg);
  binary_mux_s1_w1 \ins_dec/mux14_b0  (
    .i0(id_ins_pc[0]),
    .i1(csr_data[0]),
    .sel(id_system),
    .o(\ins_dec/n270 [0]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b1  (
    .i0(id_ins_pc[1]),
    .i1(csr_data[1]),
    .sel(id_system),
    .o(\ins_dec/n270 [1]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b10  (
    .i0(id_ins_pc[10]),
    .i1(csr_data[10]),
    .sel(id_system),
    .o(\ins_dec/n270 [10]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b11  (
    .i0(id_ins_pc[11]),
    .i1(csr_data[11]),
    .sel(id_system),
    .o(\ins_dec/n270 [11]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b12  (
    .i0(id_ins_pc[12]),
    .i1(csr_data[12]),
    .sel(id_system),
    .o(\ins_dec/n270 [12]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b13  (
    .i0(id_ins_pc[13]),
    .i1(csr_data[13]),
    .sel(id_system),
    .o(\ins_dec/n270 [13]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b14  (
    .i0(id_ins_pc[14]),
    .i1(csr_data[14]),
    .sel(id_system),
    .o(\ins_dec/n270 [14]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b15  (
    .i0(id_ins_pc[15]),
    .i1(csr_data[15]),
    .sel(id_system),
    .o(\ins_dec/n270 [15]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b16  (
    .i0(id_ins_pc[16]),
    .i1(csr_data[16]),
    .sel(id_system),
    .o(\ins_dec/n270 [16]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b17  (
    .i0(id_ins_pc[17]),
    .i1(csr_data[17]),
    .sel(id_system),
    .o(\ins_dec/n270 [17]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b18  (
    .i0(id_ins_pc[18]),
    .i1(csr_data[18]),
    .sel(id_system),
    .o(\ins_dec/n270 [18]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b19  (
    .i0(id_ins_pc[19]),
    .i1(csr_data[19]),
    .sel(id_system),
    .o(\ins_dec/n270 [19]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b2  (
    .i0(id_ins_pc[2]),
    .i1(csr_data[2]),
    .sel(id_system),
    .o(\ins_dec/n270 [2]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b20  (
    .i0(id_ins_pc[20]),
    .i1(csr_data[20]),
    .sel(id_system),
    .o(\ins_dec/n270 [20]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b21  (
    .i0(id_ins_pc[21]),
    .i1(csr_data[21]),
    .sel(id_system),
    .o(\ins_dec/n270 [21]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b22  (
    .i0(id_ins_pc[22]),
    .i1(csr_data[22]),
    .sel(id_system),
    .o(\ins_dec/n270 [22]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b23  (
    .i0(id_ins_pc[23]),
    .i1(csr_data[23]),
    .sel(id_system),
    .o(\ins_dec/n270 [23]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b24  (
    .i0(id_ins_pc[24]),
    .i1(csr_data[24]),
    .sel(id_system),
    .o(\ins_dec/n270 [24]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b25  (
    .i0(id_ins_pc[25]),
    .i1(csr_data[25]),
    .sel(id_system),
    .o(\ins_dec/n270 [25]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b26  (
    .i0(id_ins_pc[26]),
    .i1(csr_data[26]),
    .sel(id_system),
    .o(\ins_dec/n270 [26]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b27  (
    .i0(id_ins_pc[27]),
    .i1(csr_data[27]),
    .sel(id_system),
    .o(\ins_dec/n270 [27]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b28  (
    .i0(id_ins_pc[28]),
    .i1(csr_data[28]),
    .sel(id_system),
    .o(\ins_dec/n270 [28]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b29  (
    .i0(id_ins_pc[29]),
    .i1(csr_data[29]),
    .sel(id_system),
    .o(\ins_dec/n270 [29]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b3  (
    .i0(id_ins_pc[3]),
    .i1(csr_data[3]),
    .sel(id_system),
    .o(\ins_dec/n270 [3]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b30  (
    .i0(id_ins_pc[30]),
    .i1(csr_data[30]),
    .sel(id_system),
    .o(\ins_dec/n270 [30]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b31  (
    .i0(id_ins_pc[31]),
    .i1(csr_data[31]),
    .sel(id_system),
    .o(\ins_dec/n270 [31]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b32  (
    .i0(id_ins_pc[32]),
    .i1(csr_data[32]),
    .sel(id_system),
    .o(\ins_dec/n270 [32]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b33  (
    .i0(id_ins_pc[33]),
    .i1(csr_data[33]),
    .sel(id_system),
    .o(\ins_dec/n270 [33]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b34  (
    .i0(id_ins_pc[34]),
    .i1(csr_data[34]),
    .sel(id_system),
    .o(\ins_dec/n270 [34]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b35  (
    .i0(id_ins_pc[35]),
    .i1(csr_data[35]),
    .sel(id_system),
    .o(\ins_dec/n270 [35]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b36  (
    .i0(id_ins_pc[36]),
    .i1(csr_data[36]),
    .sel(id_system),
    .o(\ins_dec/n270 [36]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b37  (
    .i0(id_ins_pc[37]),
    .i1(csr_data[37]),
    .sel(id_system),
    .o(\ins_dec/n270 [37]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b38  (
    .i0(id_ins_pc[38]),
    .i1(csr_data[38]),
    .sel(id_system),
    .o(\ins_dec/n270 [38]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b39  (
    .i0(id_ins_pc[39]),
    .i1(csr_data[39]),
    .sel(id_system),
    .o(\ins_dec/n270 [39]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b4  (
    .i0(id_ins_pc[4]),
    .i1(csr_data[4]),
    .sel(id_system),
    .o(\ins_dec/n270 [4]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b40  (
    .i0(id_ins_pc[40]),
    .i1(csr_data[40]),
    .sel(id_system),
    .o(\ins_dec/n270 [40]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b41  (
    .i0(id_ins_pc[41]),
    .i1(csr_data[41]),
    .sel(id_system),
    .o(\ins_dec/n270 [41]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b42  (
    .i0(id_ins_pc[42]),
    .i1(csr_data[42]),
    .sel(id_system),
    .o(\ins_dec/n270 [42]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b43  (
    .i0(id_ins_pc[43]),
    .i1(csr_data[43]),
    .sel(id_system),
    .o(\ins_dec/n270 [43]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b44  (
    .i0(id_ins_pc[44]),
    .i1(csr_data[44]),
    .sel(id_system),
    .o(\ins_dec/n270 [44]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b45  (
    .i0(id_ins_pc[45]),
    .i1(csr_data[45]),
    .sel(id_system),
    .o(\ins_dec/n270 [45]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b46  (
    .i0(id_ins_pc[46]),
    .i1(csr_data[46]),
    .sel(id_system),
    .o(\ins_dec/n270 [46]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b47  (
    .i0(id_ins_pc[47]),
    .i1(csr_data[47]),
    .sel(id_system),
    .o(\ins_dec/n270 [47]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b48  (
    .i0(id_ins_pc[48]),
    .i1(csr_data[48]),
    .sel(id_system),
    .o(\ins_dec/n270 [48]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b49  (
    .i0(id_ins_pc[49]),
    .i1(csr_data[49]),
    .sel(id_system),
    .o(\ins_dec/n270 [49]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b5  (
    .i0(id_ins_pc[5]),
    .i1(csr_data[5]),
    .sel(id_system),
    .o(\ins_dec/n270 [5]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b50  (
    .i0(id_ins_pc[50]),
    .i1(csr_data[50]),
    .sel(id_system),
    .o(\ins_dec/n270 [50]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b51  (
    .i0(id_ins_pc[51]),
    .i1(csr_data[51]),
    .sel(id_system),
    .o(\ins_dec/n270 [51]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b52  (
    .i0(id_ins_pc[52]),
    .i1(csr_data[52]),
    .sel(id_system),
    .o(\ins_dec/n270 [52]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b53  (
    .i0(id_ins_pc[53]),
    .i1(csr_data[53]),
    .sel(id_system),
    .o(\ins_dec/n270 [53]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b54  (
    .i0(id_ins_pc[54]),
    .i1(csr_data[54]),
    .sel(id_system),
    .o(\ins_dec/n270 [54]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b55  (
    .i0(id_ins_pc[55]),
    .i1(csr_data[55]),
    .sel(id_system),
    .o(\ins_dec/n270 [55]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b56  (
    .i0(id_ins_pc[56]),
    .i1(csr_data[56]),
    .sel(id_system),
    .o(\ins_dec/n270 [56]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b57  (
    .i0(id_ins_pc[57]),
    .i1(csr_data[57]),
    .sel(id_system),
    .o(\ins_dec/n270 [57]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b58  (
    .i0(id_ins_pc[58]),
    .i1(csr_data[58]),
    .sel(id_system),
    .o(\ins_dec/n270 [58]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b59  (
    .i0(id_ins_pc[59]),
    .i1(csr_data[59]),
    .sel(id_system),
    .o(\ins_dec/n270 [59]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b6  (
    .i0(id_ins_pc[6]),
    .i1(csr_data[6]),
    .sel(id_system),
    .o(\ins_dec/n270 [6]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b60  (
    .i0(id_ins_pc[60]),
    .i1(csr_data[60]),
    .sel(id_system),
    .o(\ins_dec/n270 [60]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b61  (
    .i0(id_ins_pc[61]),
    .i1(csr_data[61]),
    .sel(id_system),
    .o(\ins_dec/n270 [61]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b62  (
    .i0(id_ins_pc[62]),
    .i1(csr_data[62]),
    .sel(id_system),
    .o(\ins_dec/n270 [62]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b63  (
    .i0(id_ins_pc[63]),
    .i1(csr_data[63]),
    .sel(id_system),
    .o(\ins_dec/n270 [63]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b7  (
    .i0(id_ins_pc[7]),
    .i1(csr_data[7]),
    .sel(id_system),
    .o(\ins_dec/n270 [7]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b8  (
    .i0(id_ins_pc[8]),
    .i1(csr_data[8]),
    .sel(id_system),
    .o(\ins_dec/n270 [8]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux14_b9  (
    .i0(id_ins_pc[9]),
    .i1(csr_data[9]),
    .sel(id_system),
    .o(\ins_dec/n270 [9]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b0  (
    .i0(\ins_dec/n270 [0]),
    .i1(rs1_data[0]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [0]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b1  (
    .i0(\ins_dec/n270 [1]),
    .i1(rs1_data[1]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [1]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b10  (
    .i0(\ins_dec/n270 [10]),
    .i1(rs1_data[10]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [10]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b11  (
    .i0(\ins_dec/n270 [11]),
    .i1(rs1_data[11]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [11]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b12  (
    .i0(\ins_dec/n270 [12]),
    .i1(rs1_data[12]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [12]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b13  (
    .i0(\ins_dec/n270 [13]),
    .i1(rs1_data[13]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [13]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b14  (
    .i0(\ins_dec/n270 [14]),
    .i1(rs1_data[14]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [14]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b15  (
    .i0(\ins_dec/n270 [15]),
    .i1(rs1_data[15]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [15]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b16  (
    .i0(\ins_dec/n270 [16]),
    .i1(rs1_data[16]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [16]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b17  (
    .i0(\ins_dec/n270 [17]),
    .i1(rs1_data[17]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [17]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b18  (
    .i0(\ins_dec/n270 [18]),
    .i1(rs1_data[18]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [18]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b19  (
    .i0(\ins_dec/n270 [19]),
    .i1(rs1_data[19]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [19]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b2  (
    .i0(\ins_dec/n270 [2]),
    .i1(rs1_data[2]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [2]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b20  (
    .i0(\ins_dec/n270 [20]),
    .i1(rs1_data[20]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [20]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b21  (
    .i0(\ins_dec/n270 [21]),
    .i1(rs1_data[21]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [21]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b22  (
    .i0(\ins_dec/n270 [22]),
    .i1(rs1_data[22]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [22]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b23  (
    .i0(\ins_dec/n270 [23]),
    .i1(rs1_data[23]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [23]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b24  (
    .i0(\ins_dec/n270 [24]),
    .i1(rs1_data[24]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [24]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b25  (
    .i0(\ins_dec/n270 [25]),
    .i1(rs1_data[25]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [25]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b26  (
    .i0(\ins_dec/n270 [26]),
    .i1(rs1_data[26]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [26]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b27  (
    .i0(\ins_dec/n270 [27]),
    .i1(rs1_data[27]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [27]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b28  (
    .i0(\ins_dec/n270 [28]),
    .i1(rs1_data[28]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [28]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b29  (
    .i0(\ins_dec/n270 [29]),
    .i1(rs1_data[29]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [29]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b3  (
    .i0(\ins_dec/n270 [3]),
    .i1(rs1_data[3]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [3]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b30  (
    .i0(\ins_dec/n270 [30]),
    .i1(rs1_data[30]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [30]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b31  (
    .i0(\ins_dec/n270 [31]),
    .i1(rs1_data[31]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [31]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b32  (
    .i0(\ins_dec/n270 [32]),
    .i1(rs1_data[32]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [32]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b33  (
    .i0(\ins_dec/n270 [33]),
    .i1(rs1_data[33]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [33]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b34  (
    .i0(\ins_dec/n270 [34]),
    .i1(rs1_data[34]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [34]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b35  (
    .i0(\ins_dec/n270 [35]),
    .i1(rs1_data[35]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [35]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b36  (
    .i0(\ins_dec/n270 [36]),
    .i1(rs1_data[36]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [36]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b37  (
    .i0(\ins_dec/n270 [37]),
    .i1(rs1_data[37]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [37]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b38  (
    .i0(\ins_dec/n270 [38]),
    .i1(rs1_data[38]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [38]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b39  (
    .i0(\ins_dec/n270 [39]),
    .i1(rs1_data[39]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [39]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b4  (
    .i0(\ins_dec/n270 [4]),
    .i1(rs1_data[4]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [4]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b40  (
    .i0(\ins_dec/n270 [40]),
    .i1(rs1_data[40]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [40]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b41  (
    .i0(\ins_dec/n270 [41]),
    .i1(rs1_data[41]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [41]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b42  (
    .i0(\ins_dec/n270 [42]),
    .i1(rs1_data[42]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [42]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b43  (
    .i0(\ins_dec/n270 [43]),
    .i1(rs1_data[43]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [43]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b44  (
    .i0(\ins_dec/n270 [44]),
    .i1(rs1_data[44]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [44]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b45  (
    .i0(\ins_dec/n270 [45]),
    .i1(rs1_data[45]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [45]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b46  (
    .i0(\ins_dec/n270 [46]),
    .i1(rs1_data[46]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [46]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b47  (
    .i0(\ins_dec/n270 [47]),
    .i1(rs1_data[47]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [47]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b48  (
    .i0(\ins_dec/n270 [48]),
    .i1(rs1_data[48]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [48]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b49  (
    .i0(\ins_dec/n270 [49]),
    .i1(rs1_data[49]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [49]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b5  (
    .i0(\ins_dec/n270 [5]),
    .i1(rs1_data[5]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [5]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b50  (
    .i0(\ins_dec/n270 [50]),
    .i1(rs1_data[50]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [50]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b51  (
    .i0(\ins_dec/n270 [51]),
    .i1(rs1_data[51]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [51]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b52  (
    .i0(\ins_dec/n270 [52]),
    .i1(rs1_data[52]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [52]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b53  (
    .i0(\ins_dec/n270 [53]),
    .i1(rs1_data[53]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [53]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b54  (
    .i0(\ins_dec/n270 [54]),
    .i1(rs1_data[54]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [54]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b55  (
    .i0(\ins_dec/n270 [55]),
    .i1(rs1_data[55]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [55]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b56  (
    .i0(\ins_dec/n270 [56]),
    .i1(rs1_data[56]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [56]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b57  (
    .i0(\ins_dec/n270 [57]),
    .i1(rs1_data[57]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [57]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b58  (
    .i0(\ins_dec/n270 [58]),
    .i1(rs1_data[58]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [58]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b59  (
    .i0(\ins_dec/n270 [59]),
    .i1(rs1_data[59]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [59]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b6  (
    .i0(\ins_dec/n270 [6]),
    .i1(rs1_data[6]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [6]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b60  (
    .i0(\ins_dec/n270 [60]),
    .i1(rs1_data[60]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [60]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b61  (
    .i0(\ins_dec/n270 [61]),
    .i1(rs1_data[61]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [61]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b62  (
    .i0(\ins_dec/n270 [62]),
    .i1(rs1_data[62]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [62]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b63  (
    .i0(\ins_dec/n270 [63]),
    .i1(rs1_data[63]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [63]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b7  (
    .i0(\ins_dec/n270 [7]),
    .i1(rs1_data[7]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [7]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b8  (
    .i0(\ins_dec/n270 [8]),
    .i1(rs1_data[8]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [8]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux15_b9  (
    .i0(\ins_dec/n270 [9]),
    .i1(rs1_data[9]),
    .sel(\ins_dec/n269 ),
    .o(\ins_dec/n271 [9]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b0  (
    .i0(\ins_dec/n271 [0]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [0]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b1  (
    .i0(\ins_dec/n271 [1]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [1]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b10  (
    .i0(\ins_dec/n271 [10]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [10]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b11  (
    .i0(\ins_dec/n271 [11]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [11]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b12  (
    .i0(\ins_dec/n271 [12]),
    .i1(id_ins[12]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [12]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b13  (
    .i0(\ins_dec/n271 [13]),
    .i1(id_ins[13]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [13]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b14  (
    .i0(\ins_dec/n271 [14]),
    .i1(id_ins[14]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [14]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b15  (
    .i0(\ins_dec/n271 [15]),
    .i1(id_ins[15]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [15]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b16  (
    .i0(\ins_dec/n271 [16]),
    .i1(id_ins[16]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [16]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b17  (
    .i0(\ins_dec/n271 [17]),
    .i1(id_ins[17]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [17]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b18  (
    .i0(\ins_dec/n271 [18]),
    .i1(id_ins[18]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [18]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b19  (
    .i0(\ins_dec/n271 [19]),
    .i1(id_ins[19]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [19]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b2  (
    .i0(\ins_dec/n271 [2]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [2]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b20  (
    .i0(\ins_dec/n271 [20]),
    .i1(id_ins[20]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [20]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b21  (
    .i0(\ins_dec/n271 [21]),
    .i1(id_ins[21]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [21]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b22  (
    .i0(\ins_dec/n271 [22]),
    .i1(id_ins[22]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [22]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b23  (
    .i0(\ins_dec/n271 [23]),
    .i1(id_ins[23]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [23]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b24  (
    .i0(\ins_dec/n271 [24]),
    .i1(id_ins[24]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [24]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b25  (
    .i0(\ins_dec/n271 [25]),
    .i1(id_ins[25]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [25]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b26  (
    .i0(\ins_dec/n271 [26]),
    .i1(id_ins[26]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [26]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b27  (
    .i0(\ins_dec/n271 [27]),
    .i1(id_ins[27]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [27]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b28  (
    .i0(\ins_dec/n271 [28]),
    .i1(id_ins[28]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [28]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b29  (
    .i0(\ins_dec/n271 [29]),
    .i1(id_ins[29]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [29]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b3  (
    .i0(\ins_dec/n271 [3]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [3]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b30  (
    .i0(\ins_dec/n271 [30]),
    .i1(id_ins[30]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [30]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b31  (
    .i0(\ins_dec/n271 [31]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [31]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b32  (
    .i0(\ins_dec/n271 [32]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [32]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b33  (
    .i0(\ins_dec/n271 [33]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [33]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b34  (
    .i0(\ins_dec/n271 [34]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [34]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b35  (
    .i0(\ins_dec/n271 [35]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [35]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b36  (
    .i0(\ins_dec/n271 [36]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [36]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b37  (
    .i0(\ins_dec/n271 [37]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [37]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b38  (
    .i0(\ins_dec/n271 [38]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [38]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b39  (
    .i0(\ins_dec/n271 [39]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [39]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b4  (
    .i0(\ins_dec/n271 [4]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [4]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b40  (
    .i0(\ins_dec/n271 [40]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [40]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b41  (
    .i0(\ins_dec/n271 [41]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [41]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b42  (
    .i0(\ins_dec/n271 [42]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [42]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b43  (
    .i0(\ins_dec/n271 [43]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [43]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b44  (
    .i0(\ins_dec/n271 [44]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [44]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b45  (
    .i0(\ins_dec/n271 [45]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [45]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b46  (
    .i0(\ins_dec/n271 [46]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [46]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b47  (
    .i0(\ins_dec/n271 [47]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [47]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b48  (
    .i0(\ins_dec/n271 [48]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [48]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b49  (
    .i0(\ins_dec/n271 [49]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [49]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b5  (
    .i0(\ins_dec/n271 [5]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [5]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b50  (
    .i0(\ins_dec/n271 [50]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [50]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b51  (
    .i0(\ins_dec/n271 [51]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [51]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b52  (
    .i0(\ins_dec/n271 [52]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [52]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b53  (
    .i0(\ins_dec/n271 [53]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [53]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b54  (
    .i0(\ins_dec/n271 [54]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [54]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b55  (
    .i0(\ins_dec/n271 [55]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [55]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b56  (
    .i0(\ins_dec/n271 [56]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [56]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b57  (
    .i0(\ins_dec/n271 [57]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [57]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b58  (
    .i0(\ins_dec/n271 [58]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [58]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b59  (
    .i0(\ins_dec/n271 [59]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [59]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b6  (
    .i0(\ins_dec/n271 [6]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [6]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b60  (
    .i0(\ins_dec/n271 [60]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [60]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b61  (
    .i0(\ins_dec/n271 [61]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [61]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b62  (
    .i0(\ins_dec/n271 [62]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [62]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b63  (
    .i0(\ins_dec/n271 [63]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [63]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b7  (
    .i0(\ins_dec/n271 [7]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [7]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b8  (
    .i0(\ins_dec/n271 [8]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [8]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux16_b9  (
    .i0(\ins_dec/n271 [9]),
    .i1(1'b0),
    .sel(\ins_dec/op_lui ),
    .o(\ins_dec/n272 [9]));  // ../../RTL/CPU/ID/ins_dec.v(762)
  binary_mux_s1_w1 \ins_dec/mux17_b12  (
    .i0(1'b0),
    .i1(id_ins[12]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [12]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b13  (
    .i0(1'b0),
    .i1(id_ins[13]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [13]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b14  (
    .i0(1'b0),
    .i1(id_ins[14]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [14]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b15  (
    .i0(1'b0),
    .i1(id_ins[15]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [15]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b16  (
    .i0(1'b0),
    .i1(id_ins[16]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [16]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b17  (
    .i0(1'b0),
    .i1(id_ins[17]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [17]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b18  (
    .i0(1'b0),
    .i1(id_ins[18]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [18]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b19  (
    .i0(1'b0),
    .i1(id_ins[19]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [19]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b2  (
    .i0(1'b1),
    .i1(1'b0),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [2]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b20  (
    .i0(1'b0),
    .i1(id_ins[20]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [20]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b21  (
    .i0(1'b0),
    .i1(id_ins[21]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [21]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b22  (
    .i0(1'b0),
    .i1(id_ins[22]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [22]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b23  (
    .i0(1'b0),
    .i1(id_ins[23]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [23]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b24  (
    .i0(1'b0),
    .i1(id_ins[24]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [24]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b25  (
    .i0(1'b0),
    .i1(id_ins[25]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [25]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b26  (
    .i0(1'b0),
    .i1(id_ins[26]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [26]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b27  (
    .i0(1'b0),
    .i1(id_ins[27]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [27]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b28  (
    .i0(1'b0),
    .i1(id_ins[28]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [28]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b29  (
    .i0(1'b0),
    .i1(id_ins[29]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [29]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b30  (
    .i0(1'b0),
    .i1(id_ins[30]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [30]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux17_b31  (
    .i0(1'b0),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_auipc ),
    .o(\ins_dec/n280 [31]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b0  (
    .i0(1'b0),
    .i1(rs1_data[0]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [0]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b1  (
    .i0(1'b0),
    .i1(rs1_data[1]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [1]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b12  (
    .i0(\ins_dec/n280 [12]),
    .i1(rs1_data[12]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [12]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b13  (
    .i0(\ins_dec/n280 [13]),
    .i1(rs1_data[13]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [13]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b14  (
    .i0(\ins_dec/n280 [14]),
    .i1(rs1_data[14]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [14]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b15  (
    .i0(\ins_dec/n280 [15]),
    .i1(rs1_data[15]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [15]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b16  (
    .i0(\ins_dec/n280 [16]),
    .i1(rs1_data[16]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [16]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b17  (
    .i0(\ins_dec/n280 [17]),
    .i1(rs1_data[17]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [17]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b18  (
    .i0(\ins_dec/n280 [18]),
    .i1(rs1_data[18]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [18]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b19  (
    .i0(\ins_dec/n280 [19]),
    .i1(rs1_data[19]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [19]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b2  (
    .i0(\ins_dec/n280 [2]),
    .i1(rs1_data[2]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [2]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b20  (
    .i0(\ins_dec/n280 [20]),
    .i1(rs1_data[20]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [20]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b21  (
    .i0(\ins_dec/n280 [21]),
    .i1(rs1_data[21]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [21]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b22  (
    .i0(\ins_dec/n280 [22]),
    .i1(rs1_data[22]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [22]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b23  (
    .i0(\ins_dec/n280 [23]),
    .i1(rs1_data[23]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [23]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b24  (
    .i0(\ins_dec/n280 [24]),
    .i1(rs1_data[24]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [24]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b25  (
    .i0(\ins_dec/n280 [25]),
    .i1(rs1_data[25]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [25]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b26  (
    .i0(\ins_dec/n280 [26]),
    .i1(rs1_data[26]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [26]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b27  (
    .i0(\ins_dec/n280 [27]),
    .i1(rs1_data[27]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [27]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b28  (
    .i0(\ins_dec/n280 [28]),
    .i1(rs1_data[28]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [28]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b29  (
    .i0(\ins_dec/n280 [29]),
    .i1(rs1_data[29]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [29]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b3  (
    .i0(1'b0),
    .i1(rs1_data[3]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [3]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b30  (
    .i0(\ins_dec/n280 [30]),
    .i1(rs1_data[30]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [30]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b31  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[31]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [31]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b32  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[32]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [32]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b33  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[33]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [33]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b34  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[34]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [34]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b35  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[35]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [35]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b36  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[36]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [36]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b37  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[37]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [37]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b38  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[38]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [38]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b39  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[39]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [39]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b4  (
    .i0(1'b0),
    .i1(rs1_data[4]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [4]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b40  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[40]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [40]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b41  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[41]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [41]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b42  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[42]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [42]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b43  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[43]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [43]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b44  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[44]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [44]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b45  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[45]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [45]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b46  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[46]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [46]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b47  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[47]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [47]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b48  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[48]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [48]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b49  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[49]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [49]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b50  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[50]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [50]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b51  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[51]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [51]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b52  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[52]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [52]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b53  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[53]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [53]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b54  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[54]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [54]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b55  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[55]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [55]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b56  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[56]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [56]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b57  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[57]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [57]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b58  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[58]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [58]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b59  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[59]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [59]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b60  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[60]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [60]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b61  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[61]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [61]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b62  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[62]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [62]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux18_b63  (
    .i0(\ins_dec/n280 [31]),
    .i1(rs1_data[63]),
    .sel(\ins_dec/n279 ),
    .o(\ins_dec/n281 [63]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b0  (
    .i0(\ins_dec/n281 [0]),
    .i1(id_ins[7]),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [0]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b1  (
    .i0(\ins_dec/n281 [1]),
    .i1(id_ins[8]),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [1]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  AL_MUX \ins_dec/mux19_b10  (
    .i0(1'b0),
    .i1(rs1_data[10]),
    .sel(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(\ins_dec/n282 [10]));
  and \ins_dec/mux19_b10_sel_is_2  (\ins_dec/mux19_b10_sel_is_2_o , \ins_dec/n277_neg , \ins_dec/n279 );
  AL_MUX \ins_dec/mux19_b11  (
    .i0(1'b0),
    .i1(rs1_data[11]),
    .sel(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(\ins_dec/n282 [11]));
  binary_mux_s1_w1 \ins_dec/mux19_b12  (
    .i0(\ins_dec/n281 [12]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [12]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b13  (
    .i0(\ins_dec/n281 [13]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [13]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b14  (
    .i0(\ins_dec/n281 [14]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [14]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b15  (
    .i0(\ins_dec/n281 [15]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [15]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b16  (
    .i0(\ins_dec/n281 [16]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [16]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b17  (
    .i0(\ins_dec/n281 [17]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [17]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b18  (
    .i0(\ins_dec/n281 [18]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [18]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b19  (
    .i0(\ins_dec/n281 [19]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [19]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b2  (
    .i0(\ins_dec/n281 [2]),
    .i1(id_ins[9]),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [2]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b20  (
    .i0(\ins_dec/n281 [20]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [20]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b21  (
    .i0(\ins_dec/n281 [21]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [21]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b22  (
    .i0(\ins_dec/n281 [22]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [22]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b23  (
    .i0(\ins_dec/n281 [23]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [23]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b24  (
    .i0(\ins_dec/n281 [24]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [24]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b25  (
    .i0(\ins_dec/n281 [25]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [25]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b26  (
    .i0(\ins_dec/n281 [26]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [26]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b27  (
    .i0(\ins_dec/n281 [27]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [27]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b28  (
    .i0(\ins_dec/n281 [28]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [28]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b29  (
    .i0(\ins_dec/n281 [29]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [29]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b3  (
    .i0(\ins_dec/n281 [3]),
    .i1(id_ins[10]),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [3]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b30  (
    .i0(\ins_dec/n281 [30]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [30]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b31  (
    .i0(\ins_dec/n281 [31]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [31]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b32  (
    .i0(\ins_dec/n281 [32]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [32]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b33  (
    .i0(\ins_dec/n281 [33]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [33]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b34  (
    .i0(\ins_dec/n281 [34]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [34]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b35  (
    .i0(\ins_dec/n281 [35]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [35]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b36  (
    .i0(\ins_dec/n281 [36]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [36]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b37  (
    .i0(\ins_dec/n281 [37]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [37]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b38  (
    .i0(\ins_dec/n281 [38]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [38]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b39  (
    .i0(\ins_dec/n281 [39]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [39]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b4  (
    .i0(\ins_dec/n281 [4]),
    .i1(id_ins[11]),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [4]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b40  (
    .i0(\ins_dec/n281 [40]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [40]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b41  (
    .i0(\ins_dec/n281 [41]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [41]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b42  (
    .i0(\ins_dec/n281 [42]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [42]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b43  (
    .i0(\ins_dec/n281 [43]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [43]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b44  (
    .i0(\ins_dec/n281 [44]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [44]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b45  (
    .i0(\ins_dec/n281 [45]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [45]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b46  (
    .i0(\ins_dec/n281 [46]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [46]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b47  (
    .i0(\ins_dec/n281 [47]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [47]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b48  (
    .i0(\ins_dec/n281 [48]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [48]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b49  (
    .i0(\ins_dec/n281 [49]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [49]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  AL_MUX \ins_dec/mux19_b5  (
    .i0(1'b0),
    .i1(rs1_data[5]),
    .sel(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(\ins_dec/n282 [5]));
  binary_mux_s1_w1 \ins_dec/mux19_b50  (
    .i0(\ins_dec/n281 [50]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [50]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b51  (
    .i0(\ins_dec/n281 [51]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [51]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b52  (
    .i0(\ins_dec/n281 [52]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [52]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b53  (
    .i0(\ins_dec/n281 [53]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [53]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b54  (
    .i0(\ins_dec/n281 [54]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [54]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux19_b55  (
    .i0(\ins_dec/n281 [55]),
    .i1(1'b0),
    .sel(\ins_dec/n277 ),
    .o(\ins_dec/n282 [55]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  AL_MUX \ins_dec/mux19_b6  (
    .i0(1'b0),
    .i1(rs1_data[6]),
    .sel(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(\ins_dec/n282 [6]));
  AL_MUX \ins_dec/mux19_b7  (
    .i0(1'b0),
    .i1(rs1_data[7]),
    .sel(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(\ins_dec/n282 [7]));
  AL_MUX \ins_dec/mux19_b8  (
    .i0(1'b0),
    .i1(rs1_data[8]),
    .sel(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(\ins_dec/n282 [8]));
  AL_MUX \ins_dec/mux19_b9  (
    .i0(1'b0),
    .i1(rs1_data[9]),
    .sel(\ins_dec/mux19_b10_sel_is_2_o ),
    .o(\ins_dec/n282 [9]));
  binary_mux_s1_w1 \ins_dec/mux1_b0  (
    .i0(\ins_dec/n58 [0]),
    .i1(id_rs2_index[0]),
    .sel(\ins_dec/n55 ),
    .o(\ins_dec/op_count_decode [0]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  binary_mux_s1_w1 \ins_dec/mux1_b1  (
    .i0(\ins_dec/n58 [1]),
    .i1(id_rs2_index[1]),
    .sel(\ins_dec/n55 ),
    .o(\ins_dec/op_count_decode [1]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  binary_mux_s1_w1 \ins_dec/mux1_b2  (
    .i0(\ins_dec/n58 [2]),
    .i1(id_rs2_index[2]),
    .sel(\ins_dec/n55 ),
    .o(\ins_dec/op_count_decode [2]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  binary_mux_s1_w1 \ins_dec/mux1_b3  (
    .i0(\ins_dec/n58 [3]),
    .i1(id_rs2_index[3]),
    .sel(\ins_dec/n55 ),
    .o(\ins_dec/op_count_decode [3]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  binary_mux_s1_w1 \ins_dec/mux1_b4  (
    .i0(\ins_dec/n58 [4]),
    .i1(id_rs2_index[4]),
    .sel(\ins_dec/n55 ),
    .o(\ins_dec/op_count_decode [4]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  binary_mux_s1_w1 \ins_dec/mux1_b5  (
    .i0(\ins_dec/n58 [5]),
    .i1(1'b0),
    .sel(\ins_dec/n55 ),
    .o(\ins_dec/op_count_decode [5]));  // ../../RTL/CPU/ID/ins_dec.v(524)
  AL_MUX \ins_dec/mux1_b6  (
    .i0(1'b0),
    .i1(rs2_data[6]),
    .sel(\ins_dec/mux1_b6_sel_is_0_o ),
    .o(\ins_dec/op_count_decode [6]));
  and \ins_dec/mux1_b6_sel_is_0  (\ins_dec/mux1_b6_sel_is_0_o , \ins_dec/n55_neg , \ins_dec/n57_neg );
  AL_MUX \ins_dec/mux1_b7  (
    .i0(1'b0),
    .i1(rs2_data[7]),
    .sel(\ins_dec/mux1_b6_sel_is_0_o ),
    .o(\ins_dec/op_count_decode [7]));
  binary_mux_s1_w1 \ins_dec/mux20_b0  (
    .i0(\ins_dec/n282 [0]),
    .i1(id_ins[20]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [0]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b1  (
    .i0(\ins_dec/n282 [1]),
    .i1(id_ins[21]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [1]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b10  (
    .i0(\ins_dec/n282 [10]),
    .i1(id_ins[30]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [10]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b11  (
    .i0(\ins_dec/n282 [11]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [11]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b12  (
    .i0(\ins_dec/n282 [12]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [12]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b13  (
    .i0(\ins_dec/n282 [13]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [13]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b14  (
    .i0(\ins_dec/n282 [14]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [14]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b15  (
    .i0(\ins_dec/n282 [15]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [15]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b16  (
    .i0(\ins_dec/n282 [16]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [16]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b17  (
    .i0(\ins_dec/n282 [17]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [17]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b18  (
    .i0(\ins_dec/n282 [18]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [18]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b19  (
    .i0(\ins_dec/n282 [19]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [19]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b2  (
    .i0(\ins_dec/n282 [2]),
    .i1(id_ins[22]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [2]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b20  (
    .i0(\ins_dec/n282 [20]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [20]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b21  (
    .i0(\ins_dec/n282 [21]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [21]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b22  (
    .i0(\ins_dec/n282 [22]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [22]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b23  (
    .i0(\ins_dec/n282 [23]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [23]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b24  (
    .i0(\ins_dec/n282 [24]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [24]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b25  (
    .i0(\ins_dec/n282 [25]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [25]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b26  (
    .i0(\ins_dec/n282 [26]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [26]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b27  (
    .i0(\ins_dec/n282 [27]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [27]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b28  (
    .i0(\ins_dec/n282 [28]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [28]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b29  (
    .i0(\ins_dec/n282 [29]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [29]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b3  (
    .i0(\ins_dec/n282 [3]),
    .i1(id_ins[23]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [3]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b30  (
    .i0(\ins_dec/n282 [30]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [30]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b31  (
    .i0(\ins_dec/n282 [31]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [31]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b32  (
    .i0(\ins_dec/n282 [32]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [32]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b33  (
    .i0(\ins_dec/n282 [33]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [33]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b34  (
    .i0(\ins_dec/n282 [34]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [34]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b35  (
    .i0(\ins_dec/n282 [35]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [35]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b36  (
    .i0(\ins_dec/n282 [36]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [36]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b37  (
    .i0(\ins_dec/n282 [37]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [37]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b38  (
    .i0(\ins_dec/n282 [38]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [38]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b39  (
    .i0(\ins_dec/n282 [39]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [39]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b4  (
    .i0(\ins_dec/n282 [4]),
    .i1(id_ins[24]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [4]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b40  (
    .i0(\ins_dec/n282 [40]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [40]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b41  (
    .i0(\ins_dec/n282 [41]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [41]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b42  (
    .i0(\ins_dec/n282 [42]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [42]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b43  (
    .i0(\ins_dec/n282 [43]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [43]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b44  (
    .i0(\ins_dec/n282 [44]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [44]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b45  (
    .i0(\ins_dec/n282 [45]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [45]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b46  (
    .i0(\ins_dec/n282 [46]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [46]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b47  (
    .i0(\ins_dec/n282 [47]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [47]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b48  (
    .i0(\ins_dec/n282 [48]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [48]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b49  (
    .i0(\ins_dec/n282 [49]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [49]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b5  (
    .i0(\ins_dec/n282 [5]),
    .i1(id_ins[25]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [5]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b50  (
    .i0(\ins_dec/n282 [50]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [50]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b51  (
    .i0(\ins_dec/n282 [51]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [51]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b52  (
    .i0(\ins_dec/n282 [52]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [52]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b53  (
    .i0(\ins_dec/n282 [53]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [53]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b54  (
    .i0(\ins_dec/n282 [54]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [54]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b55  (
    .i0(\ins_dec/n282 [55]),
    .i1(id_ins[31]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [55]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  AL_MUX \ins_dec/mux20_b56  (
    .i0(1'b0),
    .i1(\ins_dec/n281 [56]),
    .sel(\ins_dec/mux20_b56_sel_is_0_o ),
    .o(\ins_dec/n283 [56]));
  and \ins_dec/mux20_b56_sel_is_0  (\ins_dec/mux20_b56_sel_is_0_o , \ins_dec/n275_neg , \ins_dec/n277_neg );
  AL_MUX \ins_dec/mux20_b57  (
    .i0(1'b0),
    .i1(\ins_dec/n281 [57]),
    .sel(\ins_dec/mux20_b56_sel_is_0_o ),
    .o(\ins_dec/n283 [57]));
  AL_MUX \ins_dec/mux20_b58  (
    .i0(1'b0),
    .i1(\ins_dec/n281 [58]),
    .sel(\ins_dec/mux20_b56_sel_is_0_o ),
    .o(\ins_dec/n283 [58]));
  AL_MUX \ins_dec/mux20_b59  (
    .i0(1'b0),
    .i1(\ins_dec/n281 [59]),
    .sel(\ins_dec/mux20_b56_sel_is_0_o ),
    .o(\ins_dec/n283 [59]));
  binary_mux_s1_w1 \ins_dec/mux20_b6  (
    .i0(\ins_dec/n282 [6]),
    .i1(id_ins[26]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [6]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  AL_MUX \ins_dec/mux20_b60  (
    .i0(1'b0),
    .i1(\ins_dec/n281 [60]),
    .sel(\ins_dec/mux20_b56_sel_is_0_o ),
    .o(\ins_dec/n283 [60]));
  AL_MUX \ins_dec/mux20_b61  (
    .i0(1'b0),
    .i1(\ins_dec/n281 [61]),
    .sel(\ins_dec/mux20_b56_sel_is_0_o ),
    .o(\ins_dec/n283 [61]));
  AL_MUX \ins_dec/mux20_b62  (
    .i0(1'b0),
    .i1(\ins_dec/n281 [62]),
    .sel(\ins_dec/mux20_b56_sel_is_0_o ),
    .o(\ins_dec/n283 [62]));
  AL_MUX \ins_dec/mux20_b63  (
    .i0(1'b0),
    .i1(\ins_dec/n281 [63]),
    .sel(\ins_dec/mux20_b56_sel_is_0_o ),
    .o(\ins_dec/n283 [63]));
  binary_mux_s1_w1 \ins_dec/mux20_b7  (
    .i0(\ins_dec/n282 [7]),
    .i1(id_ins[27]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [7]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b8  (
    .i0(\ins_dec/n282 [8]),
    .i1(id_ins[28]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [8]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux20_b9  (
    .i0(\ins_dec/n282 [9]),
    .i1(id_ins[29]),
    .sel(\ins_dec/n275 ),
    .o(\ins_dec/n283 [9]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b0  (
    .i0(\ins_dec/n283 [0]),
    .i1(rs2_data[0]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [0]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b1  (
    .i0(\ins_dec/n283 [1]),
    .i1(rs2_data[1]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [1]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b10  (
    .i0(\ins_dec/n283 [10]),
    .i1(rs2_data[10]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [10]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b11  (
    .i0(\ins_dec/n283 [11]),
    .i1(rs2_data[11]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [11]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b12  (
    .i0(\ins_dec/n283 [12]),
    .i1(rs2_data[12]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [12]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b13  (
    .i0(\ins_dec/n283 [13]),
    .i1(rs2_data[13]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [13]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b14  (
    .i0(\ins_dec/n283 [14]),
    .i1(rs2_data[14]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [14]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b15  (
    .i0(\ins_dec/n283 [15]),
    .i1(rs2_data[15]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [15]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b16  (
    .i0(\ins_dec/n283 [16]),
    .i1(rs2_data[16]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [16]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b17  (
    .i0(\ins_dec/n283 [17]),
    .i1(rs2_data[17]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [17]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b18  (
    .i0(\ins_dec/n283 [18]),
    .i1(rs2_data[18]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [18]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b19  (
    .i0(\ins_dec/n283 [19]),
    .i1(rs2_data[19]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [19]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b2  (
    .i0(\ins_dec/n283 [2]),
    .i1(rs2_data[2]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [2]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b20  (
    .i0(\ins_dec/n283 [20]),
    .i1(rs2_data[20]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [20]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b21  (
    .i0(\ins_dec/n283 [21]),
    .i1(rs2_data[21]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [21]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b22  (
    .i0(\ins_dec/n283 [22]),
    .i1(rs2_data[22]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [22]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b23  (
    .i0(\ins_dec/n283 [23]),
    .i1(rs2_data[23]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [23]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b24  (
    .i0(\ins_dec/n283 [24]),
    .i1(rs2_data[24]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [24]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b25  (
    .i0(\ins_dec/n283 [25]),
    .i1(rs2_data[25]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [25]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b26  (
    .i0(\ins_dec/n283 [26]),
    .i1(rs2_data[26]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [26]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b27  (
    .i0(\ins_dec/n283 [27]),
    .i1(rs2_data[27]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [27]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b28  (
    .i0(\ins_dec/n283 [28]),
    .i1(rs2_data[28]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [28]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b29  (
    .i0(\ins_dec/n283 [29]),
    .i1(rs2_data[29]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [29]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b3  (
    .i0(\ins_dec/n283 [3]),
    .i1(rs2_data[3]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [3]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b30  (
    .i0(\ins_dec/n283 [30]),
    .i1(rs2_data[30]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [30]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b31  (
    .i0(\ins_dec/n283 [31]),
    .i1(rs2_data[31]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [31]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b32  (
    .i0(\ins_dec/n283 [32]),
    .i1(rs2_data[32]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [32]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b33  (
    .i0(\ins_dec/n283 [33]),
    .i1(rs2_data[33]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [33]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b34  (
    .i0(\ins_dec/n283 [34]),
    .i1(rs2_data[34]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [34]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b35  (
    .i0(\ins_dec/n283 [35]),
    .i1(rs2_data[35]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [35]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b36  (
    .i0(\ins_dec/n283 [36]),
    .i1(rs2_data[36]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [36]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b37  (
    .i0(\ins_dec/n283 [37]),
    .i1(rs2_data[37]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [37]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b38  (
    .i0(\ins_dec/n283 [38]),
    .i1(rs2_data[38]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [38]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b39  (
    .i0(\ins_dec/n283 [39]),
    .i1(rs2_data[39]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [39]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b4  (
    .i0(\ins_dec/n283 [4]),
    .i1(rs2_data[4]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [4]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b40  (
    .i0(\ins_dec/n283 [40]),
    .i1(rs2_data[40]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [40]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b41  (
    .i0(\ins_dec/n283 [41]),
    .i1(rs2_data[41]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [41]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b42  (
    .i0(\ins_dec/n283 [42]),
    .i1(rs2_data[42]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [42]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b43  (
    .i0(\ins_dec/n283 [43]),
    .i1(rs2_data[43]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [43]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b44  (
    .i0(\ins_dec/n283 [44]),
    .i1(rs2_data[44]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [44]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b45  (
    .i0(\ins_dec/n283 [45]),
    .i1(rs2_data[45]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [45]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b46  (
    .i0(\ins_dec/n283 [46]),
    .i1(rs2_data[46]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [46]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b47  (
    .i0(\ins_dec/n283 [47]),
    .i1(rs2_data[47]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [47]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b48  (
    .i0(\ins_dec/n283 [48]),
    .i1(rs2_data[48]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [48]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b49  (
    .i0(\ins_dec/n283 [49]),
    .i1(rs2_data[49]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [49]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b5  (
    .i0(\ins_dec/n283 [5]),
    .i1(rs2_data[5]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [5]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b50  (
    .i0(\ins_dec/n283 [50]),
    .i1(rs2_data[50]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [50]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b51  (
    .i0(\ins_dec/n283 [51]),
    .i1(rs2_data[51]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [51]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b52  (
    .i0(\ins_dec/n283 [52]),
    .i1(rs2_data[52]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [52]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b53  (
    .i0(\ins_dec/n283 [53]),
    .i1(rs2_data[53]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [53]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b54  (
    .i0(\ins_dec/n283 [54]),
    .i1(rs2_data[54]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [54]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b55  (
    .i0(\ins_dec/n283 [55]),
    .i1(rs2_data[55]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [55]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b56  (
    .i0(\ins_dec/n283 [56]),
    .i1(rs2_data[56]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [56]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b57  (
    .i0(\ins_dec/n283 [57]),
    .i1(rs2_data[57]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [57]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b58  (
    .i0(\ins_dec/n283 [58]),
    .i1(rs2_data[58]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [58]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b59  (
    .i0(\ins_dec/n283 [59]),
    .i1(rs2_data[59]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [59]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b6  (
    .i0(\ins_dec/n283 [6]),
    .i1(rs2_data[6]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [6]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b60  (
    .i0(\ins_dec/n283 [60]),
    .i1(rs2_data[60]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [60]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b61  (
    .i0(\ins_dec/n283 [61]),
    .i1(rs2_data[61]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [61]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b62  (
    .i0(\ins_dec/n283 [62]),
    .i1(rs2_data[62]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [62]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b63  (
    .i0(\ins_dec/n283 [63]),
    .i1(rs2_data[63]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [63]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b7  (
    .i0(\ins_dec/n283 [7]),
    .i1(rs2_data[7]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [7]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b8  (
    .i0(\ins_dec/n283 [8]),
    .i1(rs2_data[8]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [8]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux21_b9  (
    .i0(\ins_dec/n283 [9]),
    .i1(rs2_data[9]),
    .sel(\ins_dec/n274 ),
    .o(\ins_dec/n284 [9]));  // ../../RTL/CPU/ID/ins_dec.v(767)
  binary_mux_s1_w1 \ins_dec/mux22_b0  (
    .i0(rs1_data[0]),
    .i1(id_ins_pc[0]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [0]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b1  (
    .i0(rs1_data[1]),
    .i1(id_ins_pc[1]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [1]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b10  (
    .i0(rs1_data[10]),
    .i1(id_ins_pc[10]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [10]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b11  (
    .i0(rs1_data[11]),
    .i1(id_ins_pc[11]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [11]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b12  (
    .i0(rs1_data[12]),
    .i1(id_ins_pc[12]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [12]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b13  (
    .i0(rs1_data[13]),
    .i1(id_ins_pc[13]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [13]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b14  (
    .i0(rs1_data[14]),
    .i1(id_ins_pc[14]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [14]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b15  (
    .i0(rs1_data[15]),
    .i1(id_ins_pc[15]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [15]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b16  (
    .i0(rs1_data[16]),
    .i1(id_ins_pc[16]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [16]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b17  (
    .i0(rs1_data[17]),
    .i1(id_ins_pc[17]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [17]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b18  (
    .i0(rs1_data[18]),
    .i1(id_ins_pc[18]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [18]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b19  (
    .i0(rs1_data[19]),
    .i1(id_ins_pc[19]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [19]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b2  (
    .i0(rs1_data[2]),
    .i1(id_ins_pc[2]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [2]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b20  (
    .i0(rs1_data[20]),
    .i1(id_ins_pc[20]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [20]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b21  (
    .i0(rs1_data[21]),
    .i1(id_ins_pc[21]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [21]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b22  (
    .i0(rs1_data[22]),
    .i1(id_ins_pc[22]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [22]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b23  (
    .i0(rs1_data[23]),
    .i1(id_ins_pc[23]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [23]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b24  (
    .i0(rs1_data[24]),
    .i1(id_ins_pc[24]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [24]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b25  (
    .i0(rs1_data[25]),
    .i1(id_ins_pc[25]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [25]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b26  (
    .i0(rs1_data[26]),
    .i1(id_ins_pc[26]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [26]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b27  (
    .i0(rs1_data[27]),
    .i1(id_ins_pc[27]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [27]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b28  (
    .i0(rs1_data[28]),
    .i1(id_ins_pc[28]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [28]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b29  (
    .i0(rs1_data[29]),
    .i1(id_ins_pc[29]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [29]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b3  (
    .i0(rs1_data[3]),
    .i1(id_ins_pc[3]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [3]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b30  (
    .i0(rs1_data[30]),
    .i1(id_ins_pc[30]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [30]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b31  (
    .i0(rs1_data[31]),
    .i1(id_ins_pc[31]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [31]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b32  (
    .i0(rs1_data[32]),
    .i1(id_ins_pc[32]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [32]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b33  (
    .i0(rs1_data[33]),
    .i1(id_ins_pc[33]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [33]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b34  (
    .i0(rs1_data[34]),
    .i1(id_ins_pc[34]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [34]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b35  (
    .i0(rs1_data[35]),
    .i1(id_ins_pc[35]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [35]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b36  (
    .i0(rs1_data[36]),
    .i1(id_ins_pc[36]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [36]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b37  (
    .i0(rs1_data[37]),
    .i1(id_ins_pc[37]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [37]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b38  (
    .i0(rs1_data[38]),
    .i1(id_ins_pc[38]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [38]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b39  (
    .i0(rs1_data[39]),
    .i1(id_ins_pc[39]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [39]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b4  (
    .i0(rs1_data[4]),
    .i1(id_ins_pc[4]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [4]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b40  (
    .i0(rs1_data[40]),
    .i1(id_ins_pc[40]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [40]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b41  (
    .i0(rs1_data[41]),
    .i1(id_ins_pc[41]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [41]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b42  (
    .i0(rs1_data[42]),
    .i1(id_ins_pc[42]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [42]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b43  (
    .i0(rs1_data[43]),
    .i1(id_ins_pc[43]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [43]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b44  (
    .i0(rs1_data[44]),
    .i1(id_ins_pc[44]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [44]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b45  (
    .i0(rs1_data[45]),
    .i1(id_ins_pc[45]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [45]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b46  (
    .i0(rs1_data[46]),
    .i1(id_ins_pc[46]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [46]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b47  (
    .i0(rs1_data[47]),
    .i1(id_ins_pc[47]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [47]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b48  (
    .i0(rs1_data[48]),
    .i1(id_ins_pc[48]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [48]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b49  (
    .i0(rs1_data[49]),
    .i1(id_ins_pc[49]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [49]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b5  (
    .i0(rs1_data[5]),
    .i1(id_ins_pc[5]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [5]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b50  (
    .i0(rs1_data[50]),
    .i1(id_ins_pc[50]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [50]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b51  (
    .i0(rs1_data[51]),
    .i1(id_ins_pc[51]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [51]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b52  (
    .i0(rs1_data[52]),
    .i1(id_ins_pc[52]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [52]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b53  (
    .i0(rs1_data[53]),
    .i1(id_ins_pc[53]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [53]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b54  (
    .i0(rs1_data[54]),
    .i1(id_ins_pc[54]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [54]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b55  (
    .i0(rs1_data[55]),
    .i1(id_ins_pc[55]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [55]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b56  (
    .i0(rs1_data[56]),
    .i1(id_ins_pc[56]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [56]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b57  (
    .i0(rs1_data[57]),
    .i1(id_ins_pc[57]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [57]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b58  (
    .i0(rs1_data[58]),
    .i1(id_ins_pc[58]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [58]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b59  (
    .i0(rs1_data[59]),
    .i1(id_ins_pc[59]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [59]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b6  (
    .i0(rs1_data[6]),
    .i1(id_ins_pc[6]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [6]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b60  (
    .i0(rs1_data[60]),
    .i1(id_ins_pc[60]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [60]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b61  (
    .i0(rs1_data[61]),
    .i1(id_ins_pc[61]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [61]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b62  (
    .i0(rs1_data[62]),
    .i1(id_ins_pc[62]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [62]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b63  (
    .i0(rs1_data[63]),
    .i1(id_ins_pc[63]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [63]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b7  (
    .i0(rs1_data[7]),
    .i1(id_ins_pc[7]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [7]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b8  (
    .i0(rs1_data[8]),
    .i1(id_ins_pc[8]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [8]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux22_b9  (
    .i0(rs1_data[9]),
    .i1(id_ins_pc[9]),
    .sel(\ins_dec/n285 ),
    .o(\ins_dec/n286 [9]));  // ../../RTL/CPU/ID/ins_dec.v(769)
  binary_mux_s1_w1 \ins_dec/mux23_b0  (
    .i0(1'b0),
    .i1(id_ins[20]),
    .sel(\ins_dec/op_load ),
    .o(\ins_dec/n287 [0]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux23_b1  (
    .i0(1'b0),
    .i1(id_ins[21]),
    .sel(\ins_dec/op_load ),
    .o(\ins_dec/n287 [1]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux23_b2  (
    .i0(1'b0),
    .i1(id_ins[22]),
    .sel(\ins_dec/op_load ),
    .o(\ins_dec/n287 [2]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux23_b3  (
    .i0(1'b0),
    .i1(id_ins[23]),
    .sel(\ins_dec/op_load ),
    .o(\ins_dec/n287 [3]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux23_b4  (
    .i0(1'b0),
    .i1(id_ins[24]),
    .sel(\ins_dec/op_load ),
    .o(\ins_dec/n287 [4]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux24_b0  (
    .i0(\ins_dec/n287 [0]),
    .i1(id_ins[7]),
    .sel(\ins_dec/op_store ),
    .o(\ins_dec/n288 [0]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux24_b1  (
    .i0(\ins_dec/n287 [1]),
    .i1(id_ins[8]),
    .sel(\ins_dec/op_store ),
    .o(\ins_dec/n288 [1]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  AL_MUX \ins_dec/mux24_b10  (
    .i0(id_ins[30]),
    .i1(1'b0),
    .sel(\ins_dec/mux24_b10_sel_is_0_o ),
    .o(\ins_dec/n288 [10]));
  and \ins_dec/mux24_b10_sel_is_0  (\ins_dec/mux24_b10_sel_is_0_o , \ins_dec/op_store_neg , \ins_dec/op_load_neg );
  AL_MUX \ins_dec/mux24_b11  (
    .i0(id_ins[31]),
    .i1(1'b0),
    .sel(\ins_dec/mux24_b10_sel_is_0_o ),
    .o(\ins_dec/n288 [11]));
  binary_mux_s1_w1 \ins_dec/mux24_b2  (
    .i0(\ins_dec/n287 [2]),
    .i1(id_ins[9]),
    .sel(\ins_dec/op_store ),
    .o(\ins_dec/n288 [2]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux24_b3  (
    .i0(\ins_dec/n287 [3]),
    .i1(id_ins[10]),
    .sel(\ins_dec/op_store ),
    .o(\ins_dec/n288 [3]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux24_b4  (
    .i0(\ins_dec/n287 [4]),
    .i1(id_ins[11]),
    .sel(\ins_dec/op_store ),
    .o(\ins_dec/n288 [4]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  AL_MUX \ins_dec/mux24_b5  (
    .i0(id_ins[25]),
    .i1(1'b0),
    .sel(\ins_dec/mux24_b10_sel_is_0_o ),
    .o(\ins_dec/n288 [5]));
  AL_MUX \ins_dec/mux24_b6  (
    .i0(id_ins[26]),
    .i1(1'b0),
    .sel(\ins_dec/mux24_b10_sel_is_0_o ),
    .o(\ins_dec/n288 [6]));
  AL_MUX \ins_dec/mux24_b7  (
    .i0(id_ins[27]),
    .i1(1'b0),
    .sel(\ins_dec/mux24_b10_sel_is_0_o ),
    .o(\ins_dec/n288 [7]));
  AL_MUX \ins_dec/mux24_b8  (
    .i0(id_ins[28]),
    .i1(1'b0),
    .sel(\ins_dec/mux24_b10_sel_is_0_o ),
    .o(\ins_dec/n288 [8]));
  AL_MUX \ins_dec/mux24_b9  (
    .i0(id_ins[29]),
    .i1(1'b0),
    .sel(\ins_dec/mux24_b10_sel_is_0_o ),
    .o(\ins_dec/n288 [9]));
  binary_mux_s1_w1 \ins_dec/mux25_b0  (
    .i0(\ins_dec/n288 [0]),
    .i1(1'b0),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [0]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b1  (
    .i0(\ins_dec/n288 [1]),
    .i1(id_ins[12]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [1]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b10  (
    .i0(\ins_dec/n288 [10]),
    .i1(id_ins[21]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [10]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b11  (
    .i0(\ins_dec/n288 [11]),
    .i1(id_ins[22]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [11]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b12  (
    .i0(\ins_dec/n288 [11]),
    .i1(id_ins[23]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [12]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b13  (
    .i0(\ins_dec/n288 [11]),
    .i1(id_ins[24]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [13]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b14  (
    .i0(\ins_dec/n288 [11]),
    .i1(id_ins[25]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [14]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b15  (
    .i0(\ins_dec/n288 [11]),
    .i1(id_ins[26]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [15]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b16  (
    .i0(\ins_dec/n288 [11]),
    .i1(id_ins[27]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [16]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b17  (
    .i0(\ins_dec/n288 [11]),
    .i1(id_ins[28]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [17]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b18  (
    .i0(\ins_dec/n288 [11]),
    .i1(id_ins[29]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [18]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b19  (
    .i0(\ins_dec/n288 [11]),
    .i1(id_ins[30]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [19]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b2  (
    .i0(\ins_dec/n288 [2]),
    .i1(id_ins[13]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [2]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b3  (
    .i0(\ins_dec/n288 [3]),
    .i1(id_ins[14]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [3]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b4  (
    .i0(\ins_dec/n288 [4]),
    .i1(id_ins[15]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [4]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b5  (
    .i0(\ins_dec/n288 [5]),
    .i1(id_ins[16]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [5]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  and \ins_dec/mux25_b56_sel_is_0  (\ins_dec/mux25_b56_sel_is_0_o , \ins_dec/op_jal_neg , \ins_dec/op_store_neg );
  not \ins_dec/mux25_b56_sel_is_0_o_inv  (\ins_dec/mux25_b56_sel_is_0_o_neg , \ins_dec/mux25_b56_sel_is_0_o );
  binary_mux_s1_w1 \ins_dec/mux25_b6  (
    .i0(\ins_dec/n288 [6]),
    .i1(id_ins[17]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [6]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b7  (
    .i0(\ins_dec/n288 [7]),
    .i1(id_ins[18]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [7]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b8  (
    .i0(\ins_dec/n288 [8]),
    .i1(id_ins[19]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [8]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux25_b9  (
    .i0(\ins_dec/n288 [9]),
    .i1(id_ins[20]),
    .sel(\ins_dec/op_jal ),
    .o(\ins_dec/n289 [9]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux26_b0  (
    .i0(\ins_dec/n289 [0]),
    .i1(id_ins[20]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [0]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux26_b1  (
    .i0(\ins_dec/n289 [1]),
    .i1(id_ins[21]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [1]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux26_b10  (
    .i0(\ins_dec/n289 [10]),
    .i1(id_ins[30]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [10]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux26_b11  (
    .i0(\ins_dec/n289 [11]),
    .i1(id_ins[31]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [11]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux26_b2  (
    .i0(\ins_dec/n289 [2]),
    .i1(id_ins[22]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [2]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  and \ins_dec/mux26_b20_sel_is_0  (\ins_dec/mux26_b20_sel_is_0_o , \ins_dec/op_jalr_neg , \ins_dec/op_jal_neg );
  binary_mux_s1_w1 \ins_dec/mux26_b3  (
    .i0(\ins_dec/n289 [3]),
    .i1(id_ins[23]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [3]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux26_b4  (
    .i0(\ins_dec/n289 [4]),
    .i1(id_ins[24]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [4]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux26_b5  (
    .i0(\ins_dec/n289 [5]),
    .i1(id_ins[25]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [5]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  and \ins_dec/mux26_b56_sel_is_0  (\ins_dec/mux26_b56_sel_is_0_o , \ins_dec/op_jalr_neg , \ins_dec/mux25_b56_sel_is_0_o_neg );
  not \ins_dec/mux26_b56_sel_is_0_o_inv  (\ins_dec/mux26_b56_sel_is_0_o_neg , \ins_dec/mux26_b56_sel_is_0_o );
  binary_mux_s1_w1 \ins_dec/mux26_b6  (
    .i0(\ins_dec/n289 [6]),
    .i1(id_ins[26]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [6]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux26_b7  (
    .i0(\ins_dec/n289 [7]),
    .i1(id_ins[27]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [7]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux26_b8  (
    .i0(\ins_dec/n289 [8]),
    .i1(id_ins[28]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [8]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux26_b9  (
    .i0(\ins_dec/n289 [9]),
    .i1(id_ins[29]),
    .sel(\ins_dec/op_jalr ),
    .o(\ins_dec/n290 [9]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux27_b0  (
    .i0(\ins_dec/n290 [0]),
    .i1(1'b0),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [0]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux27_b1  (
    .i0(\ins_dec/n290 [1]),
    .i1(id_ins[7]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [1]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux27_b10  (
    .i0(\ins_dec/n290 [10]),
    .i1(id_ins[29]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [10]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux27_b11  (
    .i0(\ins_dec/n290 [11]),
    .i1(id_ins[30]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [11]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  AL_MUX \ins_dec/mux27_b12  (
    .i0(id_ins[31]),
    .i1(\ins_dec/n289 [12]),
    .sel(\ins_dec/mux27_b12_sel_is_0_o ),
    .o(\ins_dec/n291 [12]));
  and \ins_dec/mux27_b12_sel_is_0  (\ins_dec/mux27_b12_sel_is_0_o , \ins_dec/op_branch_neg , \ins_dec/op_jalr_neg );
  AL_MUX \ins_dec/mux27_b13  (
    .i0(id_ins[31]),
    .i1(\ins_dec/n289 [13]),
    .sel(\ins_dec/mux27_b12_sel_is_0_o ),
    .o(\ins_dec/n291 [13]));
  AL_MUX \ins_dec/mux27_b14  (
    .i0(id_ins[31]),
    .i1(\ins_dec/n289 [14]),
    .sel(\ins_dec/mux27_b12_sel_is_0_o ),
    .o(\ins_dec/n291 [14]));
  AL_MUX \ins_dec/mux27_b15  (
    .i0(id_ins[31]),
    .i1(\ins_dec/n289 [15]),
    .sel(\ins_dec/mux27_b12_sel_is_0_o ),
    .o(\ins_dec/n291 [15]));
  AL_MUX \ins_dec/mux27_b16  (
    .i0(id_ins[31]),
    .i1(\ins_dec/n289 [16]),
    .sel(\ins_dec/mux27_b12_sel_is_0_o ),
    .o(\ins_dec/n291 [16]));
  AL_MUX \ins_dec/mux27_b17  (
    .i0(id_ins[31]),
    .i1(\ins_dec/n289 [17]),
    .sel(\ins_dec/mux27_b12_sel_is_0_o ),
    .o(\ins_dec/n291 [17]));
  AL_MUX \ins_dec/mux27_b18  (
    .i0(id_ins[31]),
    .i1(\ins_dec/n289 [18]),
    .sel(\ins_dec/mux27_b12_sel_is_0_o ),
    .o(\ins_dec/n291 [18]));
  AL_MUX \ins_dec/mux27_b19  (
    .i0(id_ins[31]),
    .i1(\ins_dec/n289 [19]),
    .sel(\ins_dec/mux27_b12_sel_is_0_o ),
    .o(\ins_dec/n291 [19]));
  binary_mux_s1_w1 \ins_dec/mux27_b2  (
    .i0(\ins_dec/n290 [2]),
    .i1(id_ins[8]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [2]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  AL_MUX \ins_dec/mux27_b20  (
    .i0(id_ins[31]),
    .i1(\ins_dec/n288 [11]),
    .sel(\ins_dec/mux27_b20_sel_is_2_o ),
    .o(\ins_dec/n291 [20]));
  and \ins_dec/mux27_b20_sel_is_2  (\ins_dec/mux27_b20_sel_is_2_o , \ins_dec/op_branch_neg , \ins_dec/mux26_b20_sel_is_0_o );
  binary_mux_s1_w1 \ins_dec/mux27_b3  (
    .i0(\ins_dec/n290 [3]),
    .i1(id_ins[9]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [3]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux27_b4  (
    .i0(\ins_dec/n290 [4]),
    .i1(id_ins[10]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [4]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux27_b5  (
    .i0(\ins_dec/n290 [5]),
    .i1(id_ins[11]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [5]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  AL_MUX \ins_dec/mux27_b56  (
    .i0(id_ins[31]),
    .i1(1'b0),
    .sel(\ins_dec/mux27_b56_sel_is_0_o ),
    .o(\ins_dec/n291 [56]));
  and \ins_dec/mux27_b56_sel_is_0  (\ins_dec/mux27_b56_sel_is_0_o , \ins_dec/op_branch_neg , \ins_dec/mux26_b56_sel_is_0_o_neg );
  binary_mux_s1_w1 \ins_dec/mux27_b6  (
    .i0(\ins_dec/n290 [6]),
    .i1(id_ins[25]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [6]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux27_b7  (
    .i0(\ins_dec/n290 [7]),
    .i1(id_ins[26]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [7]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux27_b8  (
    .i0(\ins_dec/n290 [8]),
    .i1(id_ins[27]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [8]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux27_b9  (
    .i0(\ins_dec/n290 [9]),
    .i1(id_ins[28]),
    .sel(\ins_dec/op_branch ),
    .o(\ins_dec/n291 [9]));  // ../../RTL/CPU/ID/ins_dec.v(774)
  binary_mux_s1_w1 \ins_dec/mux2_b0  (
    .i0(id_ins[15]),
    .i1(1'b0),
    .sel(\ins_dec/n61 ),
    .o(id_rs1_index[0]));  // ../../RTL/CPU/ID/ins_dec.v(529)
  binary_mux_s1_w1 \ins_dec/mux2_b1  (
    .i0(id_ins[16]),
    .i1(1'b0),
    .sel(\ins_dec/n61 ),
    .o(id_rs1_index[1]));  // ../../RTL/CPU/ID/ins_dec.v(529)
  binary_mux_s1_w1 \ins_dec/mux2_b2  (
    .i0(id_ins[17]),
    .i1(1'b0),
    .sel(\ins_dec/n61 ),
    .o(id_rs1_index[2]));  // ../../RTL/CPU/ID/ins_dec.v(529)
  binary_mux_s1_w1 \ins_dec/mux2_b3  (
    .i0(id_ins[18]),
    .i1(1'b0),
    .sel(\ins_dec/n61 ),
    .o(id_rs1_index[3]));  // ../../RTL/CPU/ID/ins_dec.v(529)
  binary_mux_s1_w1 \ins_dec/mux2_b4  (
    .i0(id_ins[19]),
    .i1(1'b0),
    .sel(\ins_dec/n61 ),
    .o(id_rs1_index[4]));  // ../../RTL/CPU/ID/ins_dec.v(529)
  binary_mux_s1_w1 \ins_dec/mux38_b0  (
    .i0(1'b0),
    .i1(id_ins[0]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [0]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b1  (
    .i0(1'b0),
    .i1(id_ins[1]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [1]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b10  (
    .i0(1'b0),
    .i1(id_ins[10]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [10]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b11  (
    .i0(1'b0),
    .i1(id_ins[11]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [11]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b12  (
    .i0(1'b0),
    .i1(id_ins[12]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [12]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b13  (
    .i0(1'b0),
    .i1(id_ins[13]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [13]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b14  (
    .i0(1'b0),
    .i1(id_ins[14]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [14]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b15  (
    .i0(1'b0),
    .i1(id_ins[15]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [15]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b16  (
    .i0(1'b0),
    .i1(id_ins[16]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [16]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b17  (
    .i0(1'b0),
    .i1(id_ins[17]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [17]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b18  (
    .i0(1'b0),
    .i1(id_ins[18]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [18]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b19  (
    .i0(1'b0),
    .i1(id_ins[19]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [19]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b2  (
    .i0(1'b0),
    .i1(id_ins[2]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [2]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b20  (
    .i0(1'b0),
    .i1(id_ins[20]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [20]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b21  (
    .i0(1'b0),
    .i1(id_ins[21]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [21]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b22  (
    .i0(1'b0),
    .i1(id_ins[22]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [22]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b23  (
    .i0(1'b0),
    .i1(id_ins[23]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [23]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b24  (
    .i0(1'b0),
    .i1(id_ins[24]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [24]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b25  (
    .i0(1'b0),
    .i1(id_ins[25]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [25]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b26  (
    .i0(1'b0),
    .i1(id_ins[26]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [26]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b27  (
    .i0(1'b0),
    .i1(id_ins[27]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [27]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b28  (
    .i0(1'b0),
    .i1(id_ins[28]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [28]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b29  (
    .i0(1'b0),
    .i1(id_ins[29]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [29]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b3  (
    .i0(1'b0),
    .i1(id_ins[3]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [3]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b30  (
    .i0(1'b0),
    .i1(id_ins[30]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [30]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b31  (
    .i0(1'b0),
    .i1(id_ins[31]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [31]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b4  (
    .i0(1'b0),
    .i1(id_ins[4]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [4]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b5  (
    .i0(1'b0),
    .i1(id_ins[5]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [5]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b6  (
    .i0(1'b0),
    .i1(id_ins[6]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [6]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b7  (
    .i0(1'b0),
    .i1(id_ins[7]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [7]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b8  (
    .i0(1'b0),
    .i1(id_ins[8]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [8]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux38_b9  (
    .i0(1'b0),
    .i1(id_ins[9]),
    .sel(id_ill_ins),
    .o(\ins_dec/n342 [9]));  // ../../RTL/CPU/ID/ins_dec.v(845)
  binary_mux_s1_w1 \ins_dec/mux3_b0  (
    .i0(1'b0),
    .i1(id_ins[20]),
    .sel(\ins_dec/n65 ),
    .o(id_rs2_index[0]));  // ../../RTL/CPU/ID/ins_dec.v(530)
  binary_mux_s1_w1 \ins_dec/mux3_b1  (
    .i0(1'b0),
    .i1(id_ins[21]),
    .sel(\ins_dec/n65 ),
    .o(id_rs2_index[1]));  // ../../RTL/CPU/ID/ins_dec.v(530)
  binary_mux_s1_w1 \ins_dec/mux3_b2  (
    .i0(1'b0),
    .i1(id_ins[22]),
    .sel(\ins_dec/n65 ),
    .o(id_rs2_index[2]));  // ../../RTL/CPU/ID/ins_dec.v(530)
  binary_mux_s1_w1 \ins_dec/mux3_b3  (
    .i0(1'b0),
    .i1(id_ins[23]),
    .sel(\ins_dec/n65 ),
    .o(id_rs2_index[3]));  // ../../RTL/CPU/ID/ins_dec.v(530)
  binary_mux_s1_w1 \ins_dec/mux3_b4  (
    .i0(1'b0),
    .i1(id_ins[24]),
    .sel(\ins_dec/n65 ),
    .o(id_rs2_index[4]));  // ../../RTL/CPU/ID/ins_dec.v(530)
  not \ins_dec/n107_inv  (\ins_dec/n107_neg , \ins_dec/n107 );
  not \ins_dec/n275_inv  (\ins_dec/n275_neg , \ins_dec/n275 );
  not \ins_dec/n277_inv  (\ins_dec/n277_neg , \ins_dec/n277 );
  not \ins_dec/n55_inv  (\ins_dec/n55_neg , \ins_dec/n55 );
  not \ins_dec/n57_inv  (\ins_dec/n57_neg , \ins_dec/n57 );
  not \ins_dec/op_branch_inv  (\ins_dec/op_branch_neg , \ins_dec/op_branch );
  not \ins_dec/op_jal_inv  (\ins_dec/op_jal_neg , \ins_dec/op_jal );
  not \ins_dec/op_jalr_inv  (\ins_dec/op_jalr_neg , \ins_dec/op_jalr );
  not \ins_dec/op_load_inv  (\ins_dec/op_load_neg , \ins_dec/op_load );
  not \ins_dec/op_store_inv  (\ins_dec/op_store_neg , \ins_dec/op_store );
  reg_sr_as_w1 \ins_dec/rd_data_add_reg  (
    .clk(clk),
    .d(\ins_dec/n132 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_add));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_and_reg  (
    .clk(clk),
    .d(\ins_dec/n134 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_and));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_ds1_reg  (
    .clk(clk),
    .d(\ins_dec/n126 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_ds1));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_or_reg  (
    .clk(clk),
    .d(\ins_dec/n135 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_or));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_slt_reg  (
    .clk(clk),
    .d(\ins_dec/n139 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_slt));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_sub_reg  (
    .clk(clk),
    .d(\ins_dec/n133 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_sub));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/rd_data_xor_reg  (
    .clk(clk),
    .d(\ins_dec/n136 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(rd_data_xor));  // ../../RTL/CPU/ID/ins_dec.v(636)
  reg_sr_as_w1 \ins_dec/reg0_b0  (
    .clk(clk),
    .d(\ins_dec/sbyte ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_size[0]));  // ../../RTL/CPU/ID/ins_dec.v(689)
  reg_sr_as_w1 \ins_dec/reg0_b1  (
    .clk(clk),
    .d(\ins_dec/dbyte ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_size[1]));  // ../../RTL/CPU/ID/ins_dec.v(689)
  reg_ar_ss_w1 \ins_dec/reg0_b2  (
    .clk(clk),
    .d(\ins_dec/qbyte ),
    .en(~id_hold),
    .reset(1'b0),
    .set(\ins_dec/n107 ),
    .q(ex_size[2]));  // ../../RTL/CPU/ID/ins_dec.v(689)
  reg_sr_as_w1 \ins_dec/reg0_b3  (
    .clk(clk),
    .d(\ins_dec/obyte ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_size[3]));  // ../../RTL/CPU/ID/ins_dec.v(689)
  reg_sr_as_w1 \ins_dec/reg10_b0  (
    .clk(clk),
    .d(\ins_dec/n342 [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[0]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b1  (
    .clk(clk),
    .d(\ins_dec/n342 [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[1]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b10  (
    .clk(clk),
    .d(\ins_dec/n342 [10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[10]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b11  (
    .clk(clk),
    .d(\ins_dec/n342 [11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[11]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b12  (
    .clk(clk),
    .d(\ins_dec/n342 [12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[12]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b13  (
    .clk(clk),
    .d(\ins_dec/n342 [13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[13]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b14  (
    .clk(clk),
    .d(\ins_dec/n342 [14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[14]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b15  (
    .clk(clk),
    .d(\ins_dec/n342 [15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[15]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b16  (
    .clk(clk),
    .d(\ins_dec/n342 [16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[16]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b17  (
    .clk(clk),
    .d(\ins_dec/n342 [17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[17]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b18  (
    .clk(clk),
    .d(\ins_dec/n342 [18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[18]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b19  (
    .clk(clk),
    .d(\ins_dec/n342 [19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[19]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b2  (
    .clk(clk),
    .d(\ins_dec/n342 [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[2]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b20  (
    .clk(clk),
    .d(\ins_dec/n342 [20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[20]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b21  (
    .clk(clk),
    .d(\ins_dec/n342 [21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[21]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b22  (
    .clk(clk),
    .d(\ins_dec/n342 [22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[22]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b23  (
    .clk(clk),
    .d(\ins_dec/n342 [23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[23]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b24  (
    .clk(clk),
    .d(\ins_dec/n342 [24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[24]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b25  (
    .clk(clk),
    .d(\ins_dec/n342 [25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[25]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b26  (
    .clk(clk),
    .d(\ins_dec/n342 [26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[26]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b27  (
    .clk(clk),
    .d(\ins_dec/n342 [27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[27]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b28  (
    .clk(clk),
    .d(\ins_dec/n342 [28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[28]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b29  (
    .clk(clk),
    .d(\ins_dec/n342 [29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[29]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b3  (
    .clk(clk),
    .d(\ins_dec/n342 [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[3]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b30  (
    .clk(clk),
    .d(\ins_dec/n342 [30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[30]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b31  (
    .clk(clk),
    .d(\ins_dec/n342 [31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[31]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b4  (
    .clk(clk),
    .d(\ins_dec/n342 [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[4]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b5  (
    .clk(clk),
    .d(\ins_dec/n342 [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[5]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b6  (
    .clk(clk),
    .d(\ins_dec/n342 [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[6]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b7  (
    .clk(clk),
    .d(\ins_dec/n342 [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[7]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b8  (
    .clk(clk),
    .d(\ins_dec/n342 [8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[8]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg10_b9  (
    .clk(clk),
    .d(\ins_dec/n342 [9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_exc_code[9]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b0  (
    .clk(clk),
    .d(id_ins_pc[0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[0]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b1  (
    .clk(clk),
    .d(id_ins_pc[1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[1]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b10  (
    .clk(clk),
    .d(id_ins_pc[10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[10]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b11  (
    .clk(clk),
    .d(id_ins_pc[11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[11]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b12  (
    .clk(clk),
    .d(id_ins_pc[12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[12]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b13  (
    .clk(clk),
    .d(id_ins_pc[13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[13]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b14  (
    .clk(clk),
    .d(id_ins_pc[14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[14]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b15  (
    .clk(clk),
    .d(id_ins_pc[15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[15]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b16  (
    .clk(clk),
    .d(id_ins_pc[16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[16]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b17  (
    .clk(clk),
    .d(id_ins_pc[17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[17]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b18  (
    .clk(clk),
    .d(id_ins_pc[18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[18]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b19  (
    .clk(clk),
    .d(id_ins_pc[19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[19]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b2  (
    .clk(clk),
    .d(id_ins_pc[2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[2]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b20  (
    .clk(clk),
    .d(id_ins_pc[20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[20]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b21  (
    .clk(clk),
    .d(id_ins_pc[21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[21]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b22  (
    .clk(clk),
    .d(id_ins_pc[22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[22]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b23  (
    .clk(clk),
    .d(id_ins_pc[23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[23]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b24  (
    .clk(clk),
    .d(id_ins_pc[24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[24]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b25  (
    .clk(clk),
    .d(id_ins_pc[25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[25]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b26  (
    .clk(clk),
    .d(id_ins_pc[26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[26]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b27  (
    .clk(clk),
    .d(id_ins_pc[27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[27]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b28  (
    .clk(clk),
    .d(id_ins_pc[28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[28]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b29  (
    .clk(clk),
    .d(id_ins_pc[29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[29]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b3  (
    .clk(clk),
    .d(id_ins_pc[3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[3]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b30  (
    .clk(clk),
    .d(id_ins_pc[30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[30]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b31  (
    .clk(clk),
    .d(id_ins_pc[31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[31]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b32  (
    .clk(clk),
    .d(id_ins_pc[32]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[32]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b33  (
    .clk(clk),
    .d(id_ins_pc[33]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[33]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b34  (
    .clk(clk),
    .d(id_ins_pc[34]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[34]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b35  (
    .clk(clk),
    .d(id_ins_pc[35]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[35]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b36  (
    .clk(clk),
    .d(id_ins_pc[36]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[36]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b37  (
    .clk(clk),
    .d(id_ins_pc[37]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[37]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b38  (
    .clk(clk),
    .d(id_ins_pc[38]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[38]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b39  (
    .clk(clk),
    .d(id_ins_pc[39]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[39]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b4  (
    .clk(clk),
    .d(id_ins_pc[4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[4]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b40  (
    .clk(clk),
    .d(id_ins_pc[40]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[40]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b41  (
    .clk(clk),
    .d(id_ins_pc[41]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[41]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b42  (
    .clk(clk),
    .d(id_ins_pc[42]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[42]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b43  (
    .clk(clk),
    .d(id_ins_pc[43]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[43]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b44  (
    .clk(clk),
    .d(id_ins_pc[44]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[44]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b45  (
    .clk(clk),
    .d(id_ins_pc[45]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[45]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b46  (
    .clk(clk),
    .d(id_ins_pc[46]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[46]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b47  (
    .clk(clk),
    .d(id_ins_pc[47]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[47]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b48  (
    .clk(clk),
    .d(id_ins_pc[48]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[48]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b49  (
    .clk(clk),
    .d(id_ins_pc[49]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[49]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b5  (
    .clk(clk),
    .d(id_ins_pc[5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[5]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b50  (
    .clk(clk),
    .d(id_ins_pc[50]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[50]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b51  (
    .clk(clk),
    .d(id_ins_pc[51]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[51]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b52  (
    .clk(clk),
    .d(id_ins_pc[52]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[52]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b53  (
    .clk(clk),
    .d(id_ins_pc[53]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[53]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b54  (
    .clk(clk),
    .d(id_ins_pc[54]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[54]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b55  (
    .clk(clk),
    .d(id_ins_pc[55]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[55]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b56  (
    .clk(clk),
    .d(id_ins_pc[56]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[56]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b57  (
    .clk(clk),
    .d(id_ins_pc[57]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[57]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b58  (
    .clk(clk),
    .d(id_ins_pc[58]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[58]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b59  (
    .clk(clk),
    .d(id_ins_pc[59]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[59]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b6  (
    .clk(clk),
    .d(id_ins_pc[6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[6]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b60  (
    .clk(clk),
    .d(id_ins_pc[60]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[60]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b61  (
    .clk(clk),
    .d(id_ins_pc[61]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[61]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b62  (
    .clk(clk),
    .d(id_ins_pc[62]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[62]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b63  (
    .clk(clk),
    .d(id_ins_pc[63]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[63]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b7  (
    .clk(clk),
    .d(id_ins_pc[7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[7]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b8  (
    .clk(clk),
    .d(id_ins_pc[8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[8]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg11_b9  (
    .clk(clk),
    .d(id_ins_pc[9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_ins_pc[9]));  // ../../RTL/CPU/ID/ins_dec.v(848)
  reg_sr_as_w1 \ins_dec/reg1_b0  (
    .clk(clk),
    .d(id_ins[20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[0]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b1  (
    .clk(clk),
    .d(id_ins[21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[1]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b10  (
    .clk(clk),
    .d(id_ins[30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[10]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b11  (
    .clk(clk),
    .d(id_ins[31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[11]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b2  (
    .clk(clk),
    .d(id_ins[22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[2]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b3  (
    .clk(clk),
    .d(id_ins[23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[3]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b4  (
    .clk(clk),
    .d(id_ins[24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[4]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b5  (
    .clk(clk),
    .d(id_ins[25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[5]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b6  (
    .clk(clk),
    .d(id_ins[26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[6]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b7  (
    .clk(clk),
    .d(id_ins[27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[7]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b8  (
    .clk(clk),
    .d(id_ins[28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[8]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg1_b9  (
    .clk(clk),
    .d(id_ins[29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_csr_index[9]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_ar_as_w1 \ins_dec/reg4_b0  (
    .clk(clk),
    .d(id_ins[7]),
    .en(\ins_dec/mux13_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(ex_rd_index[0]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_ar_as_w1 \ins_dec/reg4_b1  (
    .clk(clk),
    .d(id_ins[8]),
    .en(\ins_dec/mux13_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(ex_rd_index[1]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_ar_as_w1 \ins_dec/reg4_b2  (
    .clk(clk),
    .d(id_ins[9]),
    .en(\ins_dec/mux13_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(ex_rd_index[2]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_ar_as_w1 \ins_dec/reg4_b3  (
    .clk(clk),
    .d(id_ins[10]),
    .en(\ins_dec/mux13_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(ex_rd_index[3]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_ar_as_w1 \ins_dec/reg4_b4  (
    .clk(clk),
    .d(id_ins[11]),
    .en(\ins_dec/mux13_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(ex_rd_index[4]));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/reg5_b0  (
    .clk(clk),
    .d(\ins_dec/n272 [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[0]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b1  (
    .clk(clk),
    .d(\ins_dec/n272 [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[1]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b10  (
    .clk(clk),
    .d(\ins_dec/n272 [10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[10]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b11  (
    .clk(clk),
    .d(\ins_dec/n272 [11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[11]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b12  (
    .clk(clk),
    .d(\ins_dec/n272 [12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[12]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b13  (
    .clk(clk),
    .d(\ins_dec/n272 [13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[13]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b14  (
    .clk(clk),
    .d(\ins_dec/n272 [14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[14]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b15  (
    .clk(clk),
    .d(\ins_dec/n272 [15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[15]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b16  (
    .clk(clk),
    .d(\ins_dec/n272 [16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[16]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b17  (
    .clk(clk),
    .d(\ins_dec/n272 [17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[17]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b18  (
    .clk(clk),
    .d(\ins_dec/n272 [18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[18]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b19  (
    .clk(clk),
    .d(\ins_dec/n272 [19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[19]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b2  (
    .clk(clk),
    .d(\ins_dec/n272 [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[2]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b20  (
    .clk(clk),
    .d(\ins_dec/n272 [20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[20]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b21  (
    .clk(clk),
    .d(\ins_dec/n272 [21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[21]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b22  (
    .clk(clk),
    .d(\ins_dec/n272 [22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[22]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b23  (
    .clk(clk),
    .d(\ins_dec/n272 [23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[23]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b24  (
    .clk(clk),
    .d(\ins_dec/n272 [24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[24]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b25  (
    .clk(clk),
    .d(\ins_dec/n272 [25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[25]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b26  (
    .clk(clk),
    .d(\ins_dec/n272 [26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[26]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b27  (
    .clk(clk),
    .d(\ins_dec/n272 [27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[27]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b28  (
    .clk(clk),
    .d(\ins_dec/n272 [28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[28]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b29  (
    .clk(clk),
    .d(\ins_dec/n272 [29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[29]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b3  (
    .clk(clk),
    .d(\ins_dec/n272 [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[3]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b30  (
    .clk(clk),
    .d(\ins_dec/n272 [30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[30]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b31  (
    .clk(clk),
    .d(\ins_dec/n272 [31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[31]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b32  (
    .clk(clk),
    .d(\ins_dec/n272 [32]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[32]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b33  (
    .clk(clk),
    .d(\ins_dec/n272 [33]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[33]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b34  (
    .clk(clk),
    .d(\ins_dec/n272 [34]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[34]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b35  (
    .clk(clk),
    .d(\ins_dec/n272 [35]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[35]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b36  (
    .clk(clk),
    .d(\ins_dec/n272 [36]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[36]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b37  (
    .clk(clk),
    .d(\ins_dec/n272 [37]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[37]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b38  (
    .clk(clk),
    .d(\ins_dec/n272 [38]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[38]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b39  (
    .clk(clk),
    .d(\ins_dec/n272 [39]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[39]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b4  (
    .clk(clk),
    .d(\ins_dec/n272 [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[4]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b40  (
    .clk(clk),
    .d(\ins_dec/n272 [40]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[40]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b41  (
    .clk(clk),
    .d(\ins_dec/n272 [41]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[41]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b42  (
    .clk(clk),
    .d(\ins_dec/n272 [42]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[42]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b43  (
    .clk(clk),
    .d(\ins_dec/n272 [43]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[43]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b44  (
    .clk(clk),
    .d(\ins_dec/n272 [44]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[44]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b45  (
    .clk(clk),
    .d(\ins_dec/n272 [45]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[45]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b46  (
    .clk(clk),
    .d(\ins_dec/n272 [46]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[46]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b47  (
    .clk(clk),
    .d(\ins_dec/n272 [47]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[47]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b48  (
    .clk(clk),
    .d(\ins_dec/n272 [48]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[48]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b49  (
    .clk(clk),
    .d(\ins_dec/n272 [49]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[49]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b5  (
    .clk(clk),
    .d(\ins_dec/n272 [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[5]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b50  (
    .clk(clk),
    .d(\ins_dec/n272 [50]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[50]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b51  (
    .clk(clk),
    .d(\ins_dec/n272 [51]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[51]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b52  (
    .clk(clk),
    .d(\ins_dec/n272 [52]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[52]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b53  (
    .clk(clk),
    .d(\ins_dec/n272 [53]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[53]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b54  (
    .clk(clk),
    .d(\ins_dec/n272 [54]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[54]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b55  (
    .clk(clk),
    .d(\ins_dec/n272 [55]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[55]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b56  (
    .clk(clk),
    .d(\ins_dec/n272 [56]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[56]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b57  (
    .clk(clk),
    .d(\ins_dec/n272 [57]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[57]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b58  (
    .clk(clk),
    .d(\ins_dec/n272 [58]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[58]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b59  (
    .clk(clk),
    .d(\ins_dec/n272 [59]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[59]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b6  (
    .clk(clk),
    .d(\ins_dec/n272 [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[6]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b60  (
    .clk(clk),
    .d(\ins_dec/n272 [60]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[60]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b61  (
    .clk(clk),
    .d(\ins_dec/n272 [61]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[61]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b62  (
    .clk(clk),
    .d(\ins_dec/n272 [62]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[62]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b63  (
    .clk(clk),
    .d(\ins_dec/n272 [63]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[63]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b7  (
    .clk(clk),
    .d(\ins_dec/n272 [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[7]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b8  (
    .clk(clk),
    .d(\ins_dec/n272 [8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[8]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg5_b9  (
    .clk(clk),
    .d(\ins_dec/n272 [9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds1[9]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b0  (
    .clk(clk),
    .d(\ins_dec/n284 [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[0]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b1  (
    .clk(clk),
    .d(\ins_dec/n284 [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[1]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b10  (
    .clk(clk),
    .d(\ins_dec/n284 [10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[10]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b11  (
    .clk(clk),
    .d(\ins_dec/n284 [11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[11]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b12  (
    .clk(clk),
    .d(\ins_dec/n284 [12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[12]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b13  (
    .clk(clk),
    .d(\ins_dec/n284 [13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[13]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b14  (
    .clk(clk),
    .d(\ins_dec/n284 [14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[14]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b15  (
    .clk(clk),
    .d(\ins_dec/n284 [15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[15]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b16  (
    .clk(clk),
    .d(\ins_dec/n284 [16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[16]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b17  (
    .clk(clk),
    .d(\ins_dec/n284 [17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[17]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b18  (
    .clk(clk),
    .d(\ins_dec/n284 [18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[18]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b19  (
    .clk(clk),
    .d(\ins_dec/n284 [19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[19]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b2  (
    .clk(clk),
    .d(\ins_dec/n284 [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[2]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b20  (
    .clk(clk),
    .d(\ins_dec/n284 [20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[20]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b21  (
    .clk(clk),
    .d(\ins_dec/n284 [21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[21]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b22  (
    .clk(clk),
    .d(\ins_dec/n284 [22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[22]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b23  (
    .clk(clk),
    .d(\ins_dec/n284 [23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[23]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b24  (
    .clk(clk),
    .d(\ins_dec/n284 [24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[24]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b25  (
    .clk(clk),
    .d(\ins_dec/n284 [25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[25]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b26  (
    .clk(clk),
    .d(\ins_dec/n284 [26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[26]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b27  (
    .clk(clk),
    .d(\ins_dec/n284 [27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[27]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b28  (
    .clk(clk),
    .d(\ins_dec/n284 [28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[28]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b29  (
    .clk(clk),
    .d(\ins_dec/n284 [29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[29]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b3  (
    .clk(clk),
    .d(\ins_dec/n284 [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[3]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b30  (
    .clk(clk),
    .d(\ins_dec/n284 [30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[30]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b31  (
    .clk(clk),
    .d(\ins_dec/n284 [31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[31]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b32  (
    .clk(clk),
    .d(\ins_dec/n284 [32]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[32]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b33  (
    .clk(clk),
    .d(\ins_dec/n284 [33]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[33]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b34  (
    .clk(clk),
    .d(\ins_dec/n284 [34]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[34]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b35  (
    .clk(clk),
    .d(\ins_dec/n284 [35]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[35]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b36  (
    .clk(clk),
    .d(\ins_dec/n284 [36]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[36]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b37  (
    .clk(clk),
    .d(\ins_dec/n284 [37]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[37]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b38  (
    .clk(clk),
    .d(\ins_dec/n284 [38]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[38]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b39  (
    .clk(clk),
    .d(\ins_dec/n284 [39]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[39]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b4  (
    .clk(clk),
    .d(\ins_dec/n284 [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[4]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b40  (
    .clk(clk),
    .d(\ins_dec/n284 [40]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[40]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b41  (
    .clk(clk),
    .d(\ins_dec/n284 [41]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[41]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b42  (
    .clk(clk),
    .d(\ins_dec/n284 [42]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[42]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b43  (
    .clk(clk),
    .d(\ins_dec/n284 [43]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[43]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b44  (
    .clk(clk),
    .d(\ins_dec/n284 [44]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[44]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b45  (
    .clk(clk),
    .d(\ins_dec/n284 [45]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[45]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b46  (
    .clk(clk),
    .d(\ins_dec/n284 [46]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[46]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b47  (
    .clk(clk),
    .d(\ins_dec/n284 [47]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[47]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b48  (
    .clk(clk),
    .d(\ins_dec/n284 [48]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[48]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b49  (
    .clk(clk),
    .d(\ins_dec/n284 [49]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[49]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b5  (
    .clk(clk),
    .d(\ins_dec/n284 [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[5]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b50  (
    .clk(clk),
    .d(\ins_dec/n284 [50]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[50]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b51  (
    .clk(clk),
    .d(\ins_dec/n284 [51]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[51]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b52  (
    .clk(clk),
    .d(\ins_dec/n284 [52]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[52]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b53  (
    .clk(clk),
    .d(\ins_dec/n284 [53]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[53]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b54  (
    .clk(clk),
    .d(\ins_dec/n284 [54]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[54]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b55  (
    .clk(clk),
    .d(\ins_dec/n284 [55]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[55]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b56  (
    .clk(clk),
    .d(\ins_dec/n284 [56]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[56]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b57  (
    .clk(clk),
    .d(\ins_dec/n284 [57]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[57]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b58  (
    .clk(clk),
    .d(\ins_dec/n284 [58]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[58]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b59  (
    .clk(clk),
    .d(\ins_dec/n284 [59]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[59]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b6  (
    .clk(clk),
    .d(\ins_dec/n284 [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[6]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b60  (
    .clk(clk),
    .d(\ins_dec/n284 [60]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[60]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b61  (
    .clk(clk),
    .d(\ins_dec/n284 [61]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[61]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b62  (
    .clk(clk),
    .d(\ins_dec/n284 [62]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[62]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b63  (
    .clk(clk),
    .d(\ins_dec/n284 [63]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[63]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b7  (
    .clk(clk),
    .d(\ins_dec/n284 [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[7]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b8  (
    .clk(clk),
    .d(\ins_dec/n284 [8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[8]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg6_b9  (
    .clk(clk),
    .d(\ins_dec/n284 [9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ds2[9]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b0  (
    .clk(clk),
    .d(\ins_dec/n286 [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[0]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b1  (
    .clk(clk),
    .d(\ins_dec/n286 [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[1]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b10  (
    .clk(clk),
    .d(\ins_dec/n286 [10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[10]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b11  (
    .clk(clk),
    .d(\ins_dec/n286 [11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[11]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b12  (
    .clk(clk),
    .d(\ins_dec/n286 [12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[12]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b13  (
    .clk(clk),
    .d(\ins_dec/n286 [13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[13]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b14  (
    .clk(clk),
    .d(\ins_dec/n286 [14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[14]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b15  (
    .clk(clk),
    .d(\ins_dec/n286 [15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[15]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b16  (
    .clk(clk),
    .d(\ins_dec/n286 [16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[16]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b17  (
    .clk(clk),
    .d(\ins_dec/n286 [17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[17]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b18  (
    .clk(clk),
    .d(\ins_dec/n286 [18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[18]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b19  (
    .clk(clk),
    .d(\ins_dec/n286 [19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[19]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b2  (
    .clk(clk),
    .d(\ins_dec/n286 [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[2]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b20  (
    .clk(clk),
    .d(\ins_dec/n286 [20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[20]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b21  (
    .clk(clk),
    .d(\ins_dec/n286 [21]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[21]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b22  (
    .clk(clk),
    .d(\ins_dec/n286 [22]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[22]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b23  (
    .clk(clk),
    .d(\ins_dec/n286 [23]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[23]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b24  (
    .clk(clk),
    .d(\ins_dec/n286 [24]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[24]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b25  (
    .clk(clk),
    .d(\ins_dec/n286 [25]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[25]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b26  (
    .clk(clk),
    .d(\ins_dec/n286 [26]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[26]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b27  (
    .clk(clk),
    .d(\ins_dec/n286 [27]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[27]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b28  (
    .clk(clk),
    .d(\ins_dec/n286 [28]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[28]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b29  (
    .clk(clk),
    .d(\ins_dec/n286 [29]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[29]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b3  (
    .clk(clk),
    .d(\ins_dec/n286 [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[3]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b30  (
    .clk(clk),
    .d(\ins_dec/n286 [30]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[30]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b31  (
    .clk(clk),
    .d(\ins_dec/n286 [31]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[31]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b32  (
    .clk(clk),
    .d(\ins_dec/n286 [32]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[32]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b33  (
    .clk(clk),
    .d(\ins_dec/n286 [33]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[33]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b34  (
    .clk(clk),
    .d(\ins_dec/n286 [34]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[34]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b35  (
    .clk(clk),
    .d(\ins_dec/n286 [35]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[35]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b36  (
    .clk(clk),
    .d(\ins_dec/n286 [36]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[36]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b37  (
    .clk(clk),
    .d(\ins_dec/n286 [37]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[37]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b38  (
    .clk(clk),
    .d(\ins_dec/n286 [38]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[38]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b39  (
    .clk(clk),
    .d(\ins_dec/n286 [39]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[39]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b4  (
    .clk(clk),
    .d(\ins_dec/n286 [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[4]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b40  (
    .clk(clk),
    .d(\ins_dec/n286 [40]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[40]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b41  (
    .clk(clk),
    .d(\ins_dec/n286 [41]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[41]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b42  (
    .clk(clk),
    .d(\ins_dec/n286 [42]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[42]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b43  (
    .clk(clk),
    .d(\ins_dec/n286 [43]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[43]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b44  (
    .clk(clk),
    .d(\ins_dec/n286 [44]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[44]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b45  (
    .clk(clk),
    .d(\ins_dec/n286 [45]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[45]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b46  (
    .clk(clk),
    .d(\ins_dec/n286 [46]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[46]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b47  (
    .clk(clk),
    .d(\ins_dec/n286 [47]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[47]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b48  (
    .clk(clk),
    .d(\ins_dec/n286 [48]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[48]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b49  (
    .clk(clk),
    .d(\ins_dec/n286 [49]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[49]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b5  (
    .clk(clk),
    .d(\ins_dec/n286 [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[5]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b50  (
    .clk(clk),
    .d(\ins_dec/n286 [50]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[50]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b51  (
    .clk(clk),
    .d(\ins_dec/n286 [51]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[51]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b52  (
    .clk(clk),
    .d(\ins_dec/n286 [52]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[52]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b53  (
    .clk(clk),
    .d(\ins_dec/n286 [53]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[53]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b54  (
    .clk(clk),
    .d(\ins_dec/n286 [54]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[54]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b55  (
    .clk(clk),
    .d(\ins_dec/n286 [55]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[55]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b56  (
    .clk(clk),
    .d(\ins_dec/n286 [56]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[56]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b57  (
    .clk(clk),
    .d(\ins_dec/n286 [57]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[57]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b58  (
    .clk(clk),
    .d(\ins_dec/n286 [58]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[58]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b59  (
    .clk(clk),
    .d(\ins_dec/n286 [59]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[59]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b6  (
    .clk(clk),
    .d(\ins_dec/n286 [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[6]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b60  (
    .clk(clk),
    .d(\ins_dec/n286 [60]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[60]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b61  (
    .clk(clk),
    .d(\ins_dec/n286 [61]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[61]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b62  (
    .clk(clk),
    .d(\ins_dec/n286 [62]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[62]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b63  (
    .clk(clk),
    .d(\ins_dec/n286 [63]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[63]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b7  (
    .clk(clk),
    .d(\ins_dec/n286 [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[7]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b8  (
    .clk(clk),
    .d(\ins_dec/n286 [8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[8]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg7_b9  (
    .clk(clk),
    .d(\ins_dec/n286 [9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as1[9]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b0  (
    .clk(clk),
    .d(\ins_dec/n291 [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[0]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b1  (
    .clk(clk),
    .d(\ins_dec/n291 [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[1]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b10  (
    .clk(clk),
    .d(\ins_dec/n291 [10]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[10]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b11  (
    .clk(clk),
    .d(\ins_dec/n291 [11]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[11]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b12  (
    .clk(clk),
    .d(\ins_dec/n291 [12]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[12]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b13  (
    .clk(clk),
    .d(\ins_dec/n291 [13]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[13]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b14  (
    .clk(clk),
    .d(\ins_dec/n291 [14]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[14]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b15  (
    .clk(clk),
    .d(\ins_dec/n291 [15]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[15]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b16  (
    .clk(clk),
    .d(\ins_dec/n291 [16]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[16]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b17  (
    .clk(clk),
    .d(\ins_dec/n291 [17]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[17]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b18  (
    .clk(clk),
    .d(\ins_dec/n291 [18]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[18]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b19  (
    .clk(clk),
    .d(\ins_dec/n291 [19]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[19]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b2  (
    .clk(clk),
    .d(\ins_dec/n291 [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[2]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b20  (
    .clk(clk),
    .d(\ins_dec/n291 [20]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[20]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b3  (
    .clk(clk),
    .d(\ins_dec/n291 [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[3]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b4  (
    .clk(clk),
    .d(\ins_dec/n291 [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[4]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b5  (
    .clk(clk),
    .d(\ins_dec/n291 [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[5]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b56  (
    .clk(clk),
    .d(\ins_dec/n291 [56]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[56]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b6  (
    .clk(clk),
    .d(\ins_dec/n291 [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[6]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b7  (
    .clk(clk),
    .d(\ins_dec/n291 [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[7]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b8  (
    .clk(clk),
    .d(\ins_dec/n291 [8]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[8]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg8_b9  (
    .clk(clk),
    .d(\ins_dec/n291 [9]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(as2[9]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b0  (
    .clk(clk),
    .d(\ins_dec/op_count_decode [0]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[0]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b1  (
    .clk(clk),
    .d(\ins_dec/op_count_decode [1]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[1]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b2  (
    .clk(clk),
    .d(\ins_dec/op_count_decode [2]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[2]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b3  (
    .clk(clk),
    .d(\ins_dec/op_count_decode [3]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[3]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b4  (
    .clk(clk),
    .d(\ins_dec/op_count_decode [4]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[4]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b5  (
    .clk(clk),
    .d(\ins_dec/op_count_decode [5]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[5]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b6  (
    .clk(clk),
    .d(\ins_dec/op_count_decode [6]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[6]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/reg9_b7  (
    .clk(clk),
    .d(\ins_dec/op_count_decode [7]),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(op_count[7]));  // ../../RTL/CPU/ID/ins_dec.v(777)
  reg_sr_as_w1 \ins_dec/s_ret_reg  (
    .clk(clk),
    .d(\ins_dec/n305 ),
    .en(\ins_dec/u461_sel_is_0_o ),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(ex_s_ret));  // ../../RTL/CPU/ID/ins_dec.v(830)
  reg_sr_as_w1 \ins_dec/shift_l_reg  (
    .clk(clk),
    .d(\ins_dec/n235 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(shift_l));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/shift_r_reg  (
    .clk(clk),
    .d(\ins_dec/n232 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(shift_r));  // ../../RTL/CPU/ID/ins_dec.v(739)
  reg_sr_as_w1 \ins_dec/store_reg  (
    .clk(clk),
    .d(\ins_dec/op_store ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(store));  // ../../RTL/CPU/ID/ins_dec.v(739)
  or \ins_dec/u10  (\ins_dec/n6 , \ins_dec/n5 , \ins_dec/ins_amoandd );  // ../../RTL/CPU/ID/ins_dec.v(341)
  and \ins_dec/u100  (\ins_dec/n34 , \ins_dec/op_reg , \ins_dec/funct3_7 );  // ../../RTL/CPU/ID/ins_dec.v(454)
  and \ins_dec/u101  (\ins_dec/ins_and , \ins_dec/n34 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(454)
  or \ins_dec/u102  (\ins_dec/n35 , \ins_dec/funct3_0 , \ins_dec/funct3_1 );  // ../../RTL/CPU/ID/ins_dec.v(455)
  and \ins_dec/u103  (\ins_dec/ins_fence , id_system, \ins_dec/n35 );  // ../../RTL/CPU/ID/ins_dec.v(455)
  and \ins_dec/u104  (\ins_dec/n36 , id_system, \ins_dec/funct3_0 );  // ../../RTL/CPU/ID/ins_dec.v(456)
  and \ins_dec/u105  (\ins_dec/ins_ecall , \ins_dec/n36 , \ins_dec/funct12_0 );  // ../../RTL/CPU/ID/ins_dec.v(456)
  and \ins_dec/u107  (\ins_dec/ins_ebreak , \ins_dec/n36 , \ins_dec/funct12_1 );  // ../../RTL/CPU/ID/ins_dec.v(457)
  and \ins_dec/u108  (\ins_dec/ins_csrrw , id_system, \ins_dec/funct3_1 );  // ../../RTL/CPU/ID/ins_dec.v(458)
  and \ins_dec/u109  (\ins_dec/ins_csrrs , id_system, \ins_dec/funct3_2 );  // ../../RTL/CPU/ID/ins_dec.v(459)
  or \ins_dec/u11  (\ins_dec/n7 , \ins_dec/n6 , \ins_dec/ins_amoorw );  // ../../RTL/CPU/ID/ins_dec.v(341)
  and \ins_dec/u110  (\ins_dec/ins_csrrc , id_system, \ins_dec/funct3_3 );  // ../../RTL/CPU/ID/ins_dec.v(460)
  and \ins_dec/u111  (\ins_dec/ins_csrrwi , id_system, \ins_dec/funct3_5 );  // ../../RTL/CPU/ID/ins_dec.v(461)
  and \ins_dec/u112  (\ins_dec/ins_csrrsi , id_system, \ins_dec/funct3_6 );  // ../../RTL/CPU/ID/ins_dec.v(462)
  and \ins_dec/u113  (\ins_dec/ins_csrrci , id_system, \ins_dec/funct3_7 );  // ../../RTL/CPU/ID/ins_dec.v(463)
  and \ins_dec/u114  (\ins_dec/ins_lwu , \ins_dec/op_load , \ins_dec/funct3_6 );  // ../../RTL/CPU/ID/ins_dec.v(465)
  and \ins_dec/u115  (\ins_dec/ins_ld , \ins_dec/op_load , \ins_dec/funct3_3 );  // ../../RTL/CPU/ID/ins_dec.v(466)
  and \ins_dec/u117  (\ins_dec/ins_addiw , \ins_dec/op_32_imm , \ins_dec/funct3_0 );  // ../../RTL/CPU/ID/ins_dec.v(468)
  and \ins_dec/u118  (\ins_dec/n37 , \ins_dec/op_32_imm , \ins_dec/funct3_1 );  // ../../RTL/CPU/ID/ins_dec.v(469)
  and \ins_dec/u119  (\ins_dec/ins_slliw , \ins_dec/n37 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(469)
  or \ins_dec/u12  (\ins_dec/n8 , \ins_dec/n7 , \ins_dec/ins_amoord );  // ../../RTL/CPU/ID/ins_dec.v(341)
  and \ins_dec/u120  (\ins_dec/n38 , \ins_dec/op_32_imm , \ins_dec/funct3_5 );  // ../../RTL/CPU/ID/ins_dec.v(470)
  and \ins_dec/u121  (\ins_dec/ins_srliw , \ins_dec/n38 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(470)
  and \ins_dec/u123  (\ins_dec/ins_sraiw , \ins_dec/n38 , \ins_dec/funct7_32 );  // ../../RTL/CPU/ID/ins_dec.v(471)
  and \ins_dec/u124  (\ins_dec/n39 , \ins_dec/op_32_reg , \ins_dec/funct3_0 );  // ../../RTL/CPU/ID/ins_dec.v(472)
  and \ins_dec/u125  (\ins_dec/ins_addw , \ins_dec/n39 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(472)
  and \ins_dec/u127  (\ins_dec/ins_subw , \ins_dec/n39 , \ins_dec/funct7_32 );  // ../../RTL/CPU/ID/ins_dec.v(473)
  and \ins_dec/u128  (\ins_dec/n40 , \ins_dec/op_32_reg , \ins_dec/funct3_1 );  // ../../RTL/CPU/ID/ins_dec.v(474)
  and \ins_dec/u129  (\ins_dec/ins_sllw , \ins_dec/n40 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(474)
  or \ins_dec/u13  (\ins_dec/n9 , \ins_dec/n8 , \ins_dec/ins_amominw );  // ../../RTL/CPU/ID/ins_dec.v(341)
  and \ins_dec/u130  (\ins_dec/n41 , \ins_dec/op_32_reg , \ins_dec/funct3_5 );  // ../../RTL/CPU/ID/ins_dec.v(475)
  and \ins_dec/u131  (\ins_dec/ins_srlw , \ins_dec/n41 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(475)
  and \ins_dec/u133  (\ins_dec/ins_sraw , \ins_dec/n41 , \ins_dec/funct7_32 );  // ../../RTL/CPU/ID/ins_dec.v(476)
  and \ins_dec/u134  (\ins_dec/n42 , \ins_dec/op_amo , \ins_dec/funct3_2 );  // ../../RTL/CPU/ID/ins_dec.v(478)
  and \ins_dec/u135  (\ins_dec/ins_lrw , \ins_dec/n42 , \ins_dec/funct5_2 );  // ../../RTL/CPU/ID/ins_dec.v(478)
  and \ins_dec/u137  (\ins_dec/ins_scw , \ins_dec/n42 , \ins_dec/funct5_3 );  // ../../RTL/CPU/ID/ins_dec.v(479)
  and \ins_dec/u139  (\ins_dec/ins_amoswapw , \ins_dec/n42 , \ins_dec/funct5_1 );  // ../../RTL/CPU/ID/ins_dec.v(480)
  or \ins_dec/u14  (\ins_dec/n10 , \ins_dec/n9 , \ins_dec/ins_amomind );  // ../../RTL/CPU/ID/ins_dec.v(341)
  and \ins_dec/u141  (\ins_dec/ins_amoaddw , \ins_dec/n42 , \ins_dec/funct5_0 );  // ../../RTL/CPU/ID/ins_dec.v(481)
  and \ins_dec/u143  (\ins_dec/ins_amoxorw , \ins_dec/n42 , \ins_dec/funct5_4 );  // ../../RTL/CPU/ID/ins_dec.v(482)
  and \ins_dec/u145  (\ins_dec/ins_amoandw , \ins_dec/n42 , \ins_dec/funct5_12 );  // ../../RTL/CPU/ID/ins_dec.v(483)
  and \ins_dec/u147  (\ins_dec/ins_amoorw , \ins_dec/n42 , \ins_dec/funct5_8 );  // ../../RTL/CPU/ID/ins_dec.v(484)
  and \ins_dec/u149  (\ins_dec/ins_amominw , \ins_dec/n42 , \ins_dec/funct5_16 );  // ../../RTL/CPU/ID/ins_dec.v(485)
  or \ins_dec/u15  (\ins_dec/n11 , \ins_dec/n10 , \ins_dec/ins_amomaxw );  // ../../RTL/CPU/ID/ins_dec.v(342)
  and \ins_dec/u151  (\ins_dec/ins_amomaxw , \ins_dec/n42 , \ins_dec/funct5_20 );  // ../../RTL/CPU/ID/ins_dec.v(486)
  and \ins_dec/u153  (\ins_dec/ins_amominuw , \ins_dec/n42 , \ins_dec/funct5_24 );  // ../../RTL/CPU/ID/ins_dec.v(487)
  and \ins_dec/u155  (\ins_dec/ins_amomaxuw , \ins_dec/n42 , \ins_dec/funct5_28 );  // ../../RTL/CPU/ID/ins_dec.v(488)
  and \ins_dec/u156  (\ins_dec/n43 , \ins_dec/op_amo , \ins_dec/funct3_3 );  // ../../RTL/CPU/ID/ins_dec.v(490)
  and \ins_dec/u157  (\ins_dec/ins_lrd , \ins_dec/n43 , \ins_dec/funct5_2 );  // ../../RTL/CPU/ID/ins_dec.v(490)
  and \ins_dec/u159  (\ins_dec/ins_scd , \ins_dec/n43 , \ins_dec/funct5_3 );  // ../../RTL/CPU/ID/ins_dec.v(491)
  or \ins_dec/u16  (\ins_dec/n12 , \ins_dec/n11 , \ins_dec/ins_amomaxd );  // ../../RTL/CPU/ID/ins_dec.v(342)
  and \ins_dec/u161  (\ins_dec/ins_amoswapd , \ins_dec/n43 , \ins_dec/funct5_1 );  // ../../RTL/CPU/ID/ins_dec.v(492)
  and \ins_dec/u163  (\ins_dec/ins_amoaddd , \ins_dec/n43 , \ins_dec/funct5_0 );  // ../../RTL/CPU/ID/ins_dec.v(493)
  and \ins_dec/u165  (\ins_dec/ins_amoxord , \ins_dec/n43 , \ins_dec/funct5_4 );  // ../../RTL/CPU/ID/ins_dec.v(494)
  and \ins_dec/u167  (\ins_dec/ins_amoandd , \ins_dec/n43 , \ins_dec/funct5_12 );  // ../../RTL/CPU/ID/ins_dec.v(495)
  and \ins_dec/u169  (\ins_dec/ins_amoord , \ins_dec/n43 , \ins_dec/funct5_8 );  // ../../RTL/CPU/ID/ins_dec.v(496)
  or \ins_dec/u17  (\ins_dec/n13 , \ins_dec/ins_amomaxd , \ins_dec/ins_amomaxud );  // ../../RTL/CPU/ID/ins_dec.v(342)
  and \ins_dec/u171  (\ins_dec/ins_amomind , \ins_dec/n43 , \ins_dec/funct5_16 );  // ../../RTL/CPU/ID/ins_dec.v(497)
  and \ins_dec/u173  (\ins_dec/ins_amomaxd , \ins_dec/n43 , \ins_dec/funct5_20 );  // ../../RTL/CPU/ID/ins_dec.v(498)
  and \ins_dec/u175  (\ins_dec/ins_amominud , \ins_dec/n43 , \ins_dec/funct5_24 );  // ../../RTL/CPU/ID/ins_dec.v(499)
  and \ins_dec/u177  (\ins_dec/ins_amomaxud , \ins_dec/n43 , \ins_dec/funct5_28 );  // ../../RTL/CPU/ID/ins_dec.v(500)
  and \ins_dec/u178  (\ins_dec/n45 , id_system, \ins_dec/n44 );  // ../../RTL/CPU/ID/ins_dec.v(502)
  and \ins_dec/u179  (\ins_dec/ins_mret , \ins_dec/n45 , \ins_dec/funct7_24 );  // ../../RTL/CPU/ID/ins_dec.v(502)
  or \ins_dec/u18  (\ins_dec/n14 , \ins_dec/n13 , \ins_dec/ins_amomind );  // ../../RTL/CPU/ID/ins_dec.v(342)
  and \ins_dec/u182  (\ins_dec/ins_sret , \ins_dec/n45 , \ins_dec/funct7_8 );  // ../../RTL/CPU/ID/ins_dec.v(503)
  and \ins_dec/u183  (\ins_dec/ins_sfencevma , id_system, \ins_dec/funct7_9 );  // ../../RTL/CPU/ID/ins_dec.v(504)
  and \ins_dec/u184  (\ins_dec/ins_wfi , id_system, \ins_dec/funct7_8 );  // ../../RTL/CPU/ID/ins_dec.v(505)
  or \ins_dec/u19  (\ins_dec/n15 , \ins_dec/n14 , \ins_dec/ins_amominud );  // ../../RTL/CPU/ID/ins_dec.v(342)
  or \ins_dec/u190  (\ins_dec/n46 , \ins_dec/ins_lb , \ins_dec/ins_lbu );  // ../../RTL/CPU/ID/ins_dec.v(517)
  or \ins_dec/u191  (\ins_dec/sbyte , \ins_dec/n46 , \ins_dec/ins_sb );  // ../../RTL/CPU/ID/ins_dec.v(517)
  or \ins_dec/u192  (\ins_dec/n47 , \ins_dec/ins_lh , \ins_dec/ins_lhu );  // ../../RTL/CPU/ID/ins_dec.v(518)
  or \ins_dec/u193  (\ins_dec/dbyte , \ins_dec/n47 , \ins_dec/ins_sh );  // ../../RTL/CPU/ID/ins_dec.v(518)
  or \ins_dec/u194  (\ins_dec/n48 , \ins_dec/ins_lw , \ins_dec/ins_lwu );  // ../../RTL/CPU/ID/ins_dec.v(519)
  or \ins_dec/u195  (\ins_dec/n49 , \ins_dec/n48 , \ins_dec/ins_sw );  // ../../RTL/CPU/ID/ins_dec.v(519)
  or \ins_dec/u196  (\ins_dec/n50 , \ins_dec/n49 , \ins_dec/op_32_imm );  // ../../RTL/CPU/ID/ins_dec.v(519)
  or \ins_dec/u197  (\ins_dec/n51 , \ins_dec/n50 , \ins_dec/op_32_reg );  // ../../RTL/CPU/ID/ins_dec.v(519)
  or \ins_dec/u199  (\ins_dec/qbyte , \ins_dec/n51 , \ins_dec/n42 );  // ../../RTL/CPU/ID/ins_dec.v(519)
  or \ins_dec/u20  (\ins_dec/n16 , \ins_dec/n15 , \ins_dec/ins_lb );  // ../../RTL/CPU/ID/ins_dec.v(343)
  or \ins_dec/u200  (\ins_dec/n52 , \ins_dec/sbyte , \ins_dec/dbyte );  // ../../RTL/CPU/ID/ins_dec.v(520)
  or \ins_dec/u201  (\ins_dec/n53 , \ins_dec/n52 , \ins_dec/qbyte );  // ../../RTL/CPU/ID/ins_dec.v(520)
  not \ins_dec/u202  (\ins_dec/obyte , \ins_dec/n53 );  // ../../RTL/CPU/ID/ins_dec.v(520)
  or \ins_dec/u203  (\ins_dec/n54 , \ins_dec/ins_slliw , \ins_dec/ins_srliw );  // ../../RTL/CPU/ID/ins_dec.v(522)
  or \ins_dec/u204  (\ins_dec/n55 , \ins_dec/n54 , \ins_dec/ins_sraiw );  // ../../RTL/CPU/ID/ins_dec.v(522)
  or \ins_dec/u205  (\ins_dec/n56 , \ins_dec/ins_slli , \ins_dec/ins_srli );  // ../../RTL/CPU/ID/ins_dec.v(523)
  or \ins_dec/u206  (\ins_dec/n57 , \ins_dec/n56 , \ins_dec/ins_srai );  // ../../RTL/CPU/ID/ins_dec.v(523)
  or \ins_dec/u207  (\ins_dec/n59 , \ins_dec/op_jal , \ins_dec/op_jalr );  // ../../RTL/CPU/ID/ins_dec.v(529)
  or \ins_dec/u208  (\ins_dec/n60 , \ins_dec/n59 , \ins_dec/op_lui );  // ../../RTL/CPU/ID/ins_dec.v(529)
  or \ins_dec/u209  (\ins_dec/n61 , \ins_dec/n60 , \ins_dec/op_auipc );  // ../../RTL/CPU/ID/ins_dec.v(529)
  or \ins_dec/u21  (\ins_dec/n17 , \ins_dec/n16 , \ins_dec/ins_lbu );  // ../../RTL/CPU/ID/ins_dec.v(343)
  or \ins_dec/u210  (\ins_dec/n62 , \ins_dec/op_reg , \ins_dec/op_32_reg );  // ../../RTL/CPU/ID/ins_dec.v(530)
  or \ins_dec/u211  (\ins_dec/n63 , \ins_dec/n62 , \ins_dec/op_branch );  // ../../RTL/CPU/ID/ins_dec.v(530)
  or \ins_dec/u212  (\ins_dec/n64 , \ins_dec/n63 , \ins_dec/op_store );  // ../../RTL/CPU/ID/ins_dec.v(530)
  or \ins_dec/u213  (\ins_dec/n65 , \ins_dec/n64 , \ins_dec/op_amo );  // ../../RTL/CPU/ID/ins_dec.v(530)
  or \ins_dec/u217  (\ins_dec/n66 , \ins_dec/op_branch , \ins_dec/op_jalr );  // ../../RTL/CPU/ID/ins_dec.v(538)
  or \ins_dec/u218  (id_branch, \ins_dec/n66 , \ins_dec/op_jal );  // ../../RTL/CPU/ID/ins_dec.v(538)
  or \ins_dec/u219  (\ins_dec/n67 , \ins_dec/op_branch , \ins_dec/op_store );  // ../../RTL/CPU/ID/ins_dec.v(545)
  or \ins_dec/u22  (\ins_dec/n18 , \ins_dec/n17 , \ins_dec/ins_lh );  // ../../RTL/CPU/ID/ins_dec.v(343)
  or \ins_dec/u220  (\ins_dec/n68 , \ins_dec/n67 , \ins_dec/ins_fence );  // ../../RTL/CPU/ID/ins_dec.v(545)
  or \ins_dec/u221  (\ins_dec/n69 , \ins_dec/n68 , \ins_dec/ins_mret );  // ../../RTL/CPU/ID/ins_dec.v(545)
  or \ins_dec/u222  (\ins_dec/n70 , \ins_dec/n69 , \ins_dec/ins_sret );  // ../../RTL/CPU/ID/ins_dec.v(545)
  not \ins_dec/u223  (\ins_dec/dec_gpr_write , \ins_dec/n70 );  // ../../RTL/CPU/ID/ins_dec.v(545)
  or \ins_dec/u224  (\ins_dec/n71 , \ins_dec/ins_csrrc , \ins_dec/ins_csrrci );  // ../../RTL/CPU/ID/ins_dec.v(550)
  or \ins_dec/u225  (\ins_dec/n72 , \ins_dec/n71 , \ins_dec/ins_csrrs );  // ../../RTL/CPU/ID/ins_dec.v(550)
  or \ins_dec/u226  (\ins_dec/n73 , \ins_dec/n72 , \ins_dec/ins_csrrsi );  // ../../RTL/CPU/ID/ins_dec.v(550)
  or \ins_dec/u227  (\ins_dec/n74 , \ins_dec/n73 , \ins_dec/ins_csrrw );  // ../../RTL/CPU/ID/ins_dec.v(550)
  or \ins_dec/u228  (\ins_dec/n75 , \ins_dec/n74 , \ins_dec/ins_csrrwi );  // ../../RTL/CPU/ID/ins_dec.v(550)
  or \ins_dec/u229  (\ins_dec/n78 , \biu/cache_ctrl_logic/n52 , \biu/cache_ctrl_logic/n50 );  // ../../RTL/CPU/ID/ins_dec.v(550)
  or \ins_dec/u23  (\ins_dec/n19 , \ins_dec/n18 , \ins_dec/ins_lhu );  // ../../RTL/CPU/ID/ins_dec.v(343)
  and \ins_dec/u230  (\ins_dec/n81 , \biu/cache_ctrl_logic/n48 , \ins_dec/n80 );  // ../../RTL/CPU/ID/ins_dec.v(550)
  or \ins_dec/u231  (\ins_dec/n82 , \ins_dec/n78 , \ins_dec/n81 );  // ../../RTL/CPU/ID/ins_dec.v(550)
  AL_MUX \ins_dec/u232  (
    .i0(1'b0),
    .i1(\ins_dec/n82 ),
    .sel(\ins_dec/n75 ),
    .o(\ins_dec/dec_csr_acc_fault ));  // ../../RTL/CPU/ID/ins_dec.v(550)
  and \ins_dec/u233  (\ins_dec/n83 , tsr, \ins_dec/ins_sret );  // ../../RTL/CPU/ID/ins_dec.v(552)
  or \ins_dec/u24  (\ins_dec/n20 , \ins_dec/n19 , \ins_dec/ins_lw );  // ../../RTL/CPU/ID/ins_dec.v(343)
  and \ins_dec/u240  (\ins_dec/n84 , \ins_dec/n75 , \biu/cache_ctrl_logic/n50 );  // ../../RTL/CPU/ID/ins_dec.v(552)
  and \ins_dec/u241  (\ins_dec/n86 , \ins_dec/n84 , \cu_ru/read_satp_sel );  // ../../RTL/CPU/ID/ins_dec.v(552)
  or \ins_dec/u242  (\ins_dec/n87 , \ins_dec/ins_sfencevma , \ins_dec/n86 );  // ../../RTL/CPU/ID/ins_dec.v(552)
  and \ins_dec/u243  (\ins_dec/n88 , tvm, \ins_dec/n87 );  // ../../RTL/CPU/ID/ins_dec.v(552)
  or \ins_dec/u244  (\ins_dec/n89 , \ins_dec/n83 , \ins_dec/n88 );  // ../../RTL/CPU/ID/ins_dec.v(552)
  and \ins_dec/u245  (\ins_dec/n90 , tw, \ins_dec/ins_wfi );  // ../../RTL/CPU/ID/ins_dec.v(553)
  or \ins_dec/u246  (\ins_dec/n91 , \ins_dec/n89 , \ins_dec/n90 );  // ../../RTL/CPU/ID/ins_dec.v(553)
  and \ins_dec/u248  (\ins_dec/n92 , \biu/cache_ctrl_logic/n50 , \ins_dec/ins_mret );  // ../../RTL/CPU/ID/ins_dec.v(554)
  or \ins_dec/u249  (\ins_dec/dec_ins_unpermit , \ins_dec/n91 , \ins_dec/n92 );  // ../../RTL/CPU/ID/ins_dec.v(554)
  or \ins_dec/u25  (\ins_dec/n21 , \ins_dec/n20 , \ins_dec/ins_lwu );  // ../../RTL/CPU/ID/ins_dec.v(343)
  or \ins_dec/u250  (\ins_dec/n93 , id_system, \ins_dec/op_imm );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u251  (\ins_dec/n94 , \ins_dec/n93 , \ins_dec/op_32_imm );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u252  (\ins_dec/n95 , \ins_dec/n94 , \ins_dec/op_lui );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u253  (\ins_dec/n96 , \ins_dec/n95 , \ins_dec/op_auipc );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u254  (\ins_dec/n97 , \ins_dec/n96 , \ins_dec/op_jal );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u255  (\ins_dec/n98 , \ins_dec/n97 , \ins_dec/op_jalr );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u256  (\ins_dec/n99 , \ins_dec/n98 , \ins_dec/op_branch );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u257  (\ins_dec/n100 , \ins_dec/n99 , \ins_dec/op_store );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u258  (\ins_dec/n101 , \ins_dec/n100 , \ins_dec/op_load );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u259  (\ins_dec/n102 , \ins_dec/n101 , \ins_dec/op_reg );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u26  (\ins_dec/n22 , \ins_dec/n21 , \ins_dec/ins_ld );  // ../../RTL/CPU/ID/ins_dec.v(343)
  or \ins_dec/u260  (\ins_dec/n103 , \ins_dec/n102 , \ins_dec/op_32_reg );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u261  (\ins_dec/n104 , \ins_dec/n103 , \ins_dec/op_amo );  // ../../RTL/CPU/ID/ins_dec.v(556)
  not \ins_dec/u262  (\ins_dec/dec_ins_dec_fault , \ins_dec/n104 );  // ../../RTL/CPU/ID/ins_dec.v(556)
  or \ins_dec/u263  (\ins_dec/n105 , \ins_dec/dec_ins_unpermit , \ins_dec/dec_csr_acc_fault );  // ../../RTL/CPU/ID/ins_dec.v(557)
  or \ins_dec/u264  (id_ill_ins, \ins_dec/n105 , \ins_dec/dec_ins_dec_fault );  // ../../RTL/CPU/ID/ins_dec.v(557)
  not \ins_dec/u265  (\ins_dec/n106 , id_valid);  // ../../RTL/CPU/ID/ins_dec.v(561)
  or \ins_dec/u266  (\ins_dec/n107 , rst, \ins_dec/n106 );  // ../../RTL/CPU/ID/ins_dec.v(561)
  or \ins_dec/u267  (\ins_dec/n108 , \ins_dec/op_lui , \ins_dec/ins_slli );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u268  (\ins_dec/n109 , \ins_dec/n108 , \ins_dec/ins_slliw );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u269  (\ins_dec/n110 , \ins_dec/n109 , \ins_dec/ins_srli );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u27  (\ins_dec/n23 , \ins_dec/n22 , \ins_dec/ins_lrw );  // ../../RTL/CPU/ID/ins_dec.v(343)
  or \ins_dec/u270  (\ins_dec/n111 , \ins_dec/n110 , \ins_dec/ins_srliw );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u271  (\ins_dec/n112 , \ins_dec/n111 , \ins_dec/ins_srai );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u272  (\ins_dec/n113 , \ins_dec/n112 , \ins_dec/ins_sraiw );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u273  (\ins_dec/n114 , \ins_dec/n113 , \ins_dec/ins_sll );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u274  (\ins_dec/n115 , \ins_dec/n114 , \ins_dec/ins_sllw );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u275  (\ins_dec/n116 , \ins_dec/n115 , \ins_dec/ins_srl );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u276  (\ins_dec/n117 , \ins_dec/n116 , \ins_dec/ins_srlw );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u277  (\ins_dec/n118 , \ins_dec/n117 , \ins_dec/ins_sra );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u278  (\ins_dec/n119 , \ins_dec/n118 , \ins_dec/ins_sraw );  // ../../RTL/CPU/ID/ins_dec.v(613)
  or \ins_dec/u279  (\ins_dec/n120 , \ins_dec/n119 , \ins_dec/ins_csrrc );  // ../../RTL/CPU/ID/ins_dec.v(614)
  or \ins_dec/u28  (\ins_dec/n24 , \ins_dec/n23 , \ins_dec/ins_lrd );  // ../../RTL/CPU/ID/ins_dec.v(343)
  or \ins_dec/u280  (\ins_dec/n121 , \ins_dec/n120 , \ins_dec/ins_csrrci );  // ../../RTL/CPU/ID/ins_dec.v(614)
  or \ins_dec/u281  (\ins_dec/n122 , \ins_dec/n121 , \ins_dec/ins_csrrs );  // ../../RTL/CPU/ID/ins_dec.v(614)
  or \ins_dec/u282  (\ins_dec/n123 , \ins_dec/n122 , \ins_dec/ins_csrrsi );  // ../../RTL/CPU/ID/ins_dec.v(614)
  or \ins_dec/u283  (\ins_dec/n124 , \ins_dec/n123 , \ins_dec/ins_csrrw );  // ../../RTL/CPU/ID/ins_dec.v(614)
  or \ins_dec/u284  (\ins_dec/n125 , \ins_dec/n124 , \ins_dec/ins_csrrwi );  // ../../RTL/CPU/ID/ins_dec.v(614)
  or \ins_dec/u285  (\ins_dec/n126 , \ins_dec/n125 , \ins_dec/ds1_mem_iden );  // ../../RTL/CPU/ID/ins_dec.v(614)
  or \ins_dec/u286  (\ins_dec/n127 , \ins_dec/op_auipc , \ins_dec/op_jal );  // ../../RTL/CPU/ID/ins_dec.v(617)
  or \ins_dec/u287  (\ins_dec/n128 , \ins_dec/n127 , \ins_dec/op_jalr );  // ../../RTL/CPU/ID/ins_dec.v(617)
  or \ins_dec/u288  (\ins_dec/n129 , \ins_dec/n128 , \ins_dec/ins_addi );  // ../../RTL/CPU/ID/ins_dec.v(617)
  or \ins_dec/u289  (\ins_dec/n130 , \ins_dec/n129 , \ins_dec/ins_addiw );  // ../../RTL/CPU/ID/ins_dec.v(617)
  or \ins_dec/u29  (\ins_dec/ds1_mem_iden , \ins_dec/n12 , \ins_dec/n24 );  // ../../RTL/CPU/ID/ins_dec.v(343)
  or \ins_dec/u290  (\ins_dec/n131 , \ins_dec/n130 , \ins_dec/ins_add );  // ../../RTL/CPU/ID/ins_dec.v(617)
  or \ins_dec/u291  (\ins_dec/n132 , \ins_dec/n131 , \ins_dec/ins_addw );  // ../../RTL/CPU/ID/ins_dec.v(617)
  or \ins_dec/u292  (\ins_dec/n133 , \ins_dec/ins_sub , \ins_dec/ins_subw );  // ../../RTL/CPU/ID/ins_dec.v(618)
  or \ins_dec/u293  (\ins_dec/n134 , \ins_dec/ins_andi , \ins_dec/ins_and );  // ../../RTL/CPU/ID/ins_dec.v(619)
  or \ins_dec/u294  (\ins_dec/n135 , \ins_dec/ins_ori , \ins_dec/ins_or );  // ../../RTL/CPU/ID/ins_dec.v(620)
  or \ins_dec/u295  (\ins_dec/n136 , \ins_dec/ins_xori , \ins_dec/ins_xor );  // ../../RTL/CPU/ID/ins_dec.v(621)
  or \ins_dec/u296  (\ins_dec/n137 , \ins_dec/ins_slti , \ins_dec/ins_sltiu );  // ../../RTL/CPU/ID/ins_dec.v(622)
  or \ins_dec/u297  (\ins_dec/n138 , \ins_dec/n137 , \ins_dec/ins_slt );  // ../../RTL/CPU/ID/ins_dec.v(622)
  or \ins_dec/u298  (\ins_dec/n139 , \ins_dec/n138 , \ins_dec/ins_sltu );  // ../../RTL/CPU/ID/ins_dec.v(622)
  or \ins_dec/u300  (\ins_dec/n141 , \ins_dec/ins_csrrw , \ins_dec/ins_csrrwi );  // ../../RTL/CPU/ID/ins_dec.v(628)
  or \ins_dec/u301  (\ins_dec/n142 , \ins_dec/n141 , \ins_dec/ins_scw );  // ../../RTL/CPU/ID/ins_dec.v(628)
  or \ins_dec/u302  (\ins_dec/n143 , \ins_dec/n142 , \ins_dec/ins_scd );  // ../../RTL/CPU/ID/ins_dec.v(628)
  or \ins_dec/u303  (\ins_dec/n144 , \ins_dec/n143 , \ins_dec/ins_amoswapd );  // ../../RTL/CPU/ID/ins_dec.v(628)
  or \ins_dec/u304  (\ins_dec/n145 , \ins_dec/n144 , \ins_dec/ins_amoswapw );  // ../../RTL/CPU/ID/ins_dec.v(628)
  or \ins_dec/u305  (\ins_dec/n146 , \ins_dec/ins_amoaddd , \ins_dec/ins_addw );  // ../../RTL/CPU/ID/ins_dec.v(629)
  or \ins_dec/u307  (\ins_dec/n147 , \ins_dec/n71 , \ins_dec/ins_amoandd );  // ../../RTL/CPU/ID/ins_dec.v(630)
  or \ins_dec/u308  (\ins_dec/n148 , \ins_dec/n147 , \ins_dec/ins_amoandw );  // ../../RTL/CPU/ID/ins_dec.v(630)
  or \ins_dec/u309  (\ins_dec/n149 , \ins_dec/ins_csrrs , \ins_dec/ins_csrrsi );  // ../../RTL/CPU/ID/ins_dec.v(631)
  or \ins_dec/u310  (\ins_dec/n150 , \ins_dec/n149 , \ins_dec/ins_amoord );  // ../../RTL/CPU/ID/ins_dec.v(631)
  or \ins_dec/u311  (\ins_dec/n151 , \ins_dec/n150 , \ins_dec/ins_amoorw );  // ../../RTL/CPU/ID/ins_dec.v(631)
  or \ins_dec/u312  (\ins_dec/n152 , \ins_dec/ins_amoxord , \ins_dec/ins_amoxorw );  // ../../RTL/CPU/ID/ins_dec.v(632)
  or \ins_dec/u313  (\ins_dec/n153 , \ins_dec/ins_amomaxw , \ins_dec/ins_amomaxuw );  // ../../RTL/CPU/ID/ins_dec.v(633)
  or \ins_dec/u314  (\ins_dec/n154 , \ins_dec/n153 , \ins_dec/ins_amomaxd );  // ../../RTL/CPU/ID/ins_dec.v(633)
  or \ins_dec/u315  (\ins_dec/n155 , \ins_dec/n154 , \ins_dec/ins_amomaxud );  // ../../RTL/CPU/ID/ins_dec.v(633)
  or \ins_dec/u316  (\ins_dec/n156 , \ins_dec/ins_amominw , \ins_dec/ins_amominuw );  // ../../RTL/CPU/ID/ins_dec.v(634)
  or \ins_dec/u317  (\ins_dec/n157 , \ins_dec/n156 , \ins_dec/ins_amomind );  // ../../RTL/CPU/ID/ins_dec.v(634)
  or \ins_dec/u318  (\ins_dec/n158 , \ins_dec/n157 , \ins_dec/ins_amominud );  // ../../RTL/CPU/ID/ins_dec.v(634)
  or \ins_dec/u357  (\ins_dec/n195 , \ins_dec/ins_bltu , \ins_dec/ins_bgeu );  // ../../RTL/CPU/ID/ins_dec.v(668)
  or \ins_dec/u358  (\ins_dec/n196 , \ins_dec/n195 , \ins_dec/ins_lbu );  // ../../RTL/CPU/ID/ins_dec.v(668)
  or \ins_dec/u359  (\ins_dec/n197 , \ins_dec/n196 , \ins_dec/ins_lhu );  // ../../RTL/CPU/ID/ins_dec.v(668)
  or \ins_dec/u360  (\ins_dec/n198 , \ins_dec/n197 , \ins_dec/ins_lwu );  // ../../RTL/CPU/ID/ins_dec.v(668)
  or \ins_dec/u361  (\ins_dec/n199 , \ins_dec/n198 , \ins_dec/ins_srai );  // ../../RTL/CPU/ID/ins_dec.v(668)
  or \ins_dec/u362  (\ins_dec/n200 , \ins_dec/n199 , \ins_dec/ins_sraiw );  // ../../RTL/CPU/ID/ins_dec.v(668)
  or \ins_dec/u363  (\ins_dec/n201 , \ins_dec/n200 , \ins_dec/ins_sraw );  // ../../RTL/CPU/ID/ins_dec.v(669)
  or \ins_dec/u364  (\ins_dec/n202 , \ins_dec/n201 , \ins_dec/ins_sra );  // ../../RTL/CPU/ID/ins_dec.v(669)
  or \ins_dec/u365  (\ins_dec/n203 , \ins_dec/n202 , \ins_dec/ins_amomaxuw );  // ../../RTL/CPU/ID/ins_dec.v(669)
  or \ins_dec/u366  (\ins_dec/n204 , \ins_dec/n203 , \ins_dec/ins_amomaxud );  // ../../RTL/CPU/ID/ins_dec.v(669)
  or \ins_dec/u367  (\ins_dec/n205 , \ins_dec/n204 , \ins_dec/ins_amominud );  // ../../RTL/CPU/ID/ins_dec.v(669)
  or \ins_dec/u368  (\ins_dec/n206 , \ins_dec/n205 , \ins_dec/ins_amominuw );  // ../../RTL/CPU/ID/ins_dec.v(669)
  or \ins_dec/u390  (\ins_dec/n225 , \ins_dec/ins_sfencevma , \ins_dec/ins_fence );  // ../../RTL/CPU/ID/ins_dec.v(729)
  or \ins_dec/u391  (\ins_dec/n226 , \ins_dec/ins_srli , \ins_dec/ins_srliw );  // ../../RTL/CPU/ID/ins_dec.v(730)
  or \ins_dec/u392  (\ins_dec/n227 , \ins_dec/n226 , \ins_dec/ins_srai );  // ../../RTL/CPU/ID/ins_dec.v(730)
  or \ins_dec/u393  (\ins_dec/n228 , \ins_dec/n227 , \ins_dec/ins_sraiw );  // ../../RTL/CPU/ID/ins_dec.v(730)
  or \ins_dec/u394  (\ins_dec/n229 , \ins_dec/n228 , \ins_dec/ins_srl );  // ../../RTL/CPU/ID/ins_dec.v(730)
  or \ins_dec/u395  (\ins_dec/n230 , \ins_dec/n229 , \ins_dec/ins_srlw );  // ../../RTL/CPU/ID/ins_dec.v(730)
  or \ins_dec/u396  (\ins_dec/n231 , \ins_dec/n230 , \ins_dec/ins_sra );  // ../../RTL/CPU/ID/ins_dec.v(730)
  or \ins_dec/u397  (\ins_dec/n232 , \ins_dec/n231 , \ins_dec/ins_sraw );  // ../../RTL/CPU/ID/ins_dec.v(730)
  or \ins_dec/u398  (\ins_dec/n233 , \ins_dec/ins_slli , \ins_dec/ins_slliw );  // ../../RTL/CPU/ID/ins_dec.v(731)
  or \ins_dec/u399  (\ins_dec/n234 , \ins_dec/n233 , \ins_dec/ins_sll );  // ../../RTL/CPU/ID/ins_dec.v(731)
  or \ins_dec/u4  (\ins_dec/n0 , \ins_dec/ins_amoswapd , \ins_dec/ins_amoswapw );  // ../../RTL/CPU/ID/ins_dec.v(340)
  or \ins_dec/u400  (\ins_dec/n235 , \ins_dec/n234 , \ins_dec/ins_sllw );  // ../../RTL/CPU/ID/ins_dec.v(731)
  or \ins_dec/u402  (\ins_dec/n236 , \ins_dec/n141 , \ins_dec/ins_csrrci );  // ../../RTL/CPU/ID/ins_dec.v(732)
  or \ins_dec/u403  (\ins_dec/n237 , \ins_dec/n236 , \ins_dec/ins_csrrc );  // ../../RTL/CPU/ID/ins_dec.v(732)
  or \ins_dec/u404  (\ins_dec/n238 , \ins_dec/n237 , \ins_dec/ins_csrrs );  // ../../RTL/CPU/ID/ins_dec.v(732)
  or \ins_dec/u405  (\ins_dec/n239 , \ins_dec/n238 , \ins_dec/ins_csrrsi );  // ../../RTL/CPU/ID/ins_dec.v(732)
  or \ins_dec/u426  (\ins_dec/n266 , \ins_dec/op_branch , \ins_dec/op_reg );  // ../../RTL/CPU/ID/ins_dec.v(760)
  or \ins_dec/u427  (\ins_dec/n267 , \ins_dec/n266 , \ins_dec/op_32_reg );  // ../../RTL/CPU/ID/ins_dec.v(760)
  or \ins_dec/u428  (\ins_dec/n268 , \ins_dec/n267 , \ins_dec/op_imm );  // ../../RTL/CPU/ID/ins_dec.v(760)
  or \ins_dec/u429  (\ins_dec/n269 , \ins_dec/n268 , \ins_dec/op_32_imm );  // ../../RTL/CPU/ID/ins_dec.v(760)
  or \ins_dec/u432  (\ins_dec/n273 , \ins_dec/n267 , \ins_dec/op_store );  // ../../RTL/CPU/ID/ins_dec.v(763)
  or \ins_dec/u433  (\ins_dec/n274 , \ins_dec/n273 , \ins_dec/op_amo );  // ../../RTL/CPU/ID/ins_dec.v(763)
  or \ins_dec/u434  (\ins_dec/n275 , \ins_dec/op_32_imm , \ins_dec/op_imm );  // ../../RTL/CPU/ID/ins_dec.v(764)
  or \ins_dec/u435  (\ins_dec/n276 , \ins_dec/ins_csrrwi , \ins_dec/ins_csrrci );  // ../../RTL/CPU/ID/ins_dec.v(765)
  or \ins_dec/u436  (\ins_dec/n277 , \ins_dec/n276 , \ins_dec/ins_csrrsi );  // ../../RTL/CPU/ID/ins_dec.v(765)
  or \ins_dec/u437  (\ins_dec/n278 , \ins_dec/ins_csrrw , \ins_dec/ins_csrrc );  // ../../RTL/CPU/ID/ins_dec.v(766)
  or \ins_dec/u438  (\ins_dec/n279 , \ins_dec/n278 , \ins_dec/ins_csrrs );  // ../../RTL/CPU/ID/ins_dec.v(766)
  or \ins_dec/u439  (\ins_dec/n285 , \ins_dec/op_branch , \ins_dec/op_jal );  // ../../RTL/CPU/ID/ins_dec.v(769)
  or \ins_dec/u443  (\ins_dec/n302 , \ins_dec/n285 , \ins_dec/op_jalr );  // ../../RTL/CPU/ID/ins_dec.v(817)
  not \ins_dec/u444  (\ins_dec/n303 , id_ill_ins);  // ../../RTL/CPU/ID/ins_dec.v(824)
  and \ins_dec/u445  (\ins_dec/n304 , \ins_dec/n303 , \ins_dec/ins_mret );  // ../../RTL/CPU/ID/ins_dec.v(824)
  and \ins_dec/u447  (\ins_dec/n305 , \ins_dec/n303 , \ins_dec/ins_sret );  // ../../RTL/CPU/ID/ins_dec.v(825)
  and \ins_dec/u461_sel_is_0  (\ins_dec/u461_sel_is_0_o , id_nop_neg, id_hold_neg);
  and \ins_dec/u478_sel_is_0  (\ins_dec/u478_sel_is_0_o , \ins_dec/n107_neg , id_nop_neg);
  or \ins_dec/u5  (\ins_dec/n1 , \ins_dec/n0 , \ins_dec/ins_amoaddw );  // ../../RTL/CPU/ID/ins_dec.v(340)
  or \ins_dec/u6  (\ins_dec/n2 , \ins_dec/n1 , \ins_dec/ins_amoaddd );  // ../../RTL/CPU/ID/ins_dec.v(340)
  and \ins_dec/u60  (\ins_dec/ins_bltu , \ins_dec/op_branch , \ins_dec/funct3_6 );  // ../../RTL/CPU/ID/ins_dec.v(426)
  and \ins_dec/u61  (\ins_dec/ins_bgeu , \ins_dec/op_branch , \ins_dec/funct3_7 );  // ../../RTL/CPU/ID/ins_dec.v(427)
  and \ins_dec/u62  (\ins_dec/ins_lb , \ins_dec/op_load , \ins_dec/funct3_0 );  // ../../RTL/CPU/ID/ins_dec.v(428)
  and \ins_dec/u63  (\ins_dec/ins_lh , \ins_dec/op_load , \ins_dec/funct3_1 );  // ../../RTL/CPU/ID/ins_dec.v(429)
  and \ins_dec/u64  (\ins_dec/ins_lw , \ins_dec/op_load , \ins_dec/funct3_2 );  // ../../RTL/CPU/ID/ins_dec.v(430)
  and \ins_dec/u65  (\ins_dec/ins_lbu , \ins_dec/op_load , \ins_dec/funct3_4 );  // ../../RTL/CPU/ID/ins_dec.v(431)
  and \ins_dec/u66  (\ins_dec/ins_lhu , \ins_dec/op_load , \ins_dec/funct3_5 );  // ../../RTL/CPU/ID/ins_dec.v(432)
  and \ins_dec/u67  (\ins_dec/ins_sb , \ins_dec/op_store , \ins_dec/funct3_0 );  // ../../RTL/CPU/ID/ins_dec.v(433)
  and \ins_dec/u68  (\ins_dec/ins_sh , \ins_dec/op_store , \ins_dec/funct3_1 );  // ../../RTL/CPU/ID/ins_dec.v(434)
  and \ins_dec/u69  (\ins_dec/ins_sw , \ins_dec/op_store , \ins_dec/funct3_2 );  // ../../RTL/CPU/ID/ins_dec.v(435)
  or \ins_dec/u7  (\ins_dec/n3 , \ins_dec/n2 , \ins_dec/ins_amoxorw );  // ../../RTL/CPU/ID/ins_dec.v(340)
  and \ins_dec/u70  (\ins_dec/ins_addi , \ins_dec/op_imm , \ins_dec/funct3_0 );  // ../../RTL/CPU/ID/ins_dec.v(436)
  and \ins_dec/u71  (\ins_dec/ins_slti , \ins_dec/op_imm , \ins_dec/funct3_2 );  // ../../RTL/CPU/ID/ins_dec.v(437)
  and \ins_dec/u72  (\ins_dec/ins_sltiu , \ins_dec/op_imm , \ins_dec/funct3_3 );  // ../../RTL/CPU/ID/ins_dec.v(438)
  and \ins_dec/u73  (\ins_dec/ins_xori , \ins_dec/op_imm , \ins_dec/funct3_4 );  // ../../RTL/CPU/ID/ins_dec.v(439)
  and \ins_dec/u74  (\ins_dec/ins_ori , \ins_dec/op_imm , \ins_dec/funct3_6 );  // ../../RTL/CPU/ID/ins_dec.v(440)
  and \ins_dec/u75  (\ins_dec/ins_andi , \ins_dec/op_imm , \ins_dec/funct3_7 );  // ../../RTL/CPU/ID/ins_dec.v(441)
  and \ins_dec/u76  (\ins_dec/n25 , \ins_dec/op_imm , \ins_dec/funct3_1 );  // ../../RTL/CPU/ID/ins_dec.v(442)
  and \ins_dec/u77  (\ins_dec/ins_slli , \ins_dec/n25 , \ins_dec/funct6_0 );  // ../../RTL/CPU/ID/ins_dec.v(442)
  and \ins_dec/u78  (\ins_dec/n26 , \ins_dec/op_imm , \ins_dec/funct3_5 );  // ../../RTL/CPU/ID/ins_dec.v(443)
  and \ins_dec/u79  (\ins_dec/ins_srli , \ins_dec/n26 , \ins_dec/funct6_0 );  // ../../RTL/CPU/ID/ins_dec.v(443)
  or \ins_dec/u8  (\ins_dec/n4 , \ins_dec/n3 , \ins_dec/ins_amoxord );  // ../../RTL/CPU/ID/ins_dec.v(340)
  and \ins_dec/u81  (\ins_dec/ins_srai , \ins_dec/n26 , \ins_dec/funct6_16 );  // ../../RTL/CPU/ID/ins_dec.v(444)
  and \ins_dec/u82  (\ins_dec/n27 , \ins_dec/op_reg , \ins_dec/funct3_0 );  // ../../RTL/CPU/ID/ins_dec.v(445)
  and \ins_dec/u83  (\ins_dec/ins_add , \ins_dec/n27 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(445)
  and \ins_dec/u85  (\ins_dec/ins_sub , \ins_dec/n27 , \ins_dec/funct7_32 );  // ../../RTL/CPU/ID/ins_dec.v(446)
  and \ins_dec/u86  (\ins_dec/n28 , \ins_dec/op_reg , \ins_dec/funct3_1 );  // ../../RTL/CPU/ID/ins_dec.v(447)
  and \ins_dec/u87  (\ins_dec/ins_sll , \ins_dec/n28 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(447)
  and \ins_dec/u88  (\ins_dec/n29 , \ins_dec/op_reg , \ins_dec/funct3_2 );  // ../../RTL/CPU/ID/ins_dec.v(448)
  and \ins_dec/u89  (\ins_dec/ins_slt , \ins_dec/n29 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(448)
  or \ins_dec/u9  (\ins_dec/n5 , \ins_dec/n4 , \ins_dec/ins_amoandw );  // ../../RTL/CPU/ID/ins_dec.v(341)
  and \ins_dec/u90  (\ins_dec/n30 , \ins_dec/op_reg , \ins_dec/funct3_3 );  // ../../RTL/CPU/ID/ins_dec.v(449)
  and \ins_dec/u91  (\ins_dec/ins_sltu , \ins_dec/n30 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(449)
  and \ins_dec/u92  (\ins_dec/n31 , \ins_dec/op_reg , \ins_dec/funct3_4 );  // ../../RTL/CPU/ID/ins_dec.v(450)
  and \ins_dec/u93  (\ins_dec/ins_xor , \ins_dec/n31 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(450)
  and \ins_dec/u94  (\ins_dec/n32 , \ins_dec/op_reg , \ins_dec/funct3_5 );  // ../../RTL/CPU/ID/ins_dec.v(451)
  and \ins_dec/u95  (\ins_dec/ins_srl , \ins_dec/n32 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(451)
  and \ins_dec/u97  (\ins_dec/ins_sra , \ins_dec/n32 , \ins_dec/funct7_32 );  // ../../RTL/CPU/ID/ins_dec.v(452)
  and \ins_dec/u98  (\ins_dec/n33 , \ins_dec/op_reg , \ins_dec/funct3_6 );  // ../../RTL/CPU/ID/ins_dec.v(453)
  and \ins_dec/u99  (\ins_dec/ins_or , \ins_dec/n33 , \ins_dec/funct7_0 );  // ../../RTL/CPU/ID/ins_dec.v(453)
  reg_sr_as_w1 \ins_dec/unsign_reg  (
    .clk(clk),
    .d(\ins_dec/n206 ),
    .en(~id_hold),
    .reset(\ins_dec/n107 ),
    .set(1'b0),
    .q(unsign));  // ../../RTL/CPU/ID/ins_dec.v(674)
  reg_sr_as_w1 \ins_dec/valid_reg  (
    .clk(clk),
    .d(id_valid),
    .en(~id_hold),
    .reset(~\ins_dec/u478_sel_is_0_o ),
    .set(1'b0),
    .q(ex_valid));  // ../../RTL/CPU/ID/ins_dec.v(830)
  add_pu62_pu62_o62 \ins_fetch/add0  (
    .i0(addr_if[63:2]),
    .i1(62'b00000000000000000000000000000000000000000000000000000000000001),
    .o(\ins_fetch/n1 ));  // ../../RTL/CPU/IF/ins_fetch.v(81)
  not \ins_fetch/hold_inv  (\ins_fetch/hold_neg , \ins_fetch/hold );
  reg_sr_as_w1 \ins_fetch/hold_reg  (
    .clk(clk),
    .d(if_hold),
    .en(~\ins_fetch/u72_sel_is_1_o ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/hold ));  // ../../RTL/CPU/IF/ins_fetch.v(115)
  reg_sr_as_w1 \ins_fetch/ins_acc_fault_reg  (
    .clk(clk),
    .d(ins_acc_fault),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_acc_fault));  // ../../RTL/CPU/IF/ins_fetch.v(137)
  reg_sr_as_w1 \ins_fetch/ins_addr_mis_reg  (
    .clk(clk),
    .d(\ins_fetch/addr_mis ),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_addr_mis));  // ../../RTL/CPU/IF/ins_fetch.v(137)
  reg_sr_as_w1 \ins_fetch/ins_page_fault_reg  (
    .clk(clk),
    .d(ins_page_fault),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_page_fault));  // ../../RTL/CPU/IF/ins_fetch.v(137)
  reg_sr_as_w1 \ins_fetch/int_acc_reg  (
    .clk(clk),
    .d(int_req),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_int_acc));  // ../../RTL/CPU/IF/ins_fetch.v(137)
  binary_mux_s1_w1 \ins_fetch/mux0_b0  (
    .i0(ins_read[0]),
    .i1(ins_read[32]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [0]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b1  (
    .i0(ins_read[1]),
    .i1(ins_read[33]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [1]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b10  (
    .i0(ins_read[10]),
    .i1(ins_read[42]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [10]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b11  (
    .i0(ins_read[11]),
    .i1(ins_read[43]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [11]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b12  (
    .i0(ins_read[12]),
    .i1(ins_read[44]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [12]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b13  (
    .i0(ins_read[13]),
    .i1(ins_read[45]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [13]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b14  (
    .i0(ins_read[14]),
    .i1(ins_read[46]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [14]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b15  (
    .i0(ins_read[15]),
    .i1(ins_read[47]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [15]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b16  (
    .i0(ins_read[16]),
    .i1(ins_read[48]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [16]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b17  (
    .i0(ins_read[17]),
    .i1(ins_read[49]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [17]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b18  (
    .i0(ins_read[18]),
    .i1(ins_read[50]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [18]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b19  (
    .i0(ins_read[19]),
    .i1(ins_read[51]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [19]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b2  (
    .i0(ins_read[2]),
    .i1(ins_read[34]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [2]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b20  (
    .i0(ins_read[20]),
    .i1(ins_read[52]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [20]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b21  (
    .i0(ins_read[21]),
    .i1(ins_read[53]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [21]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b22  (
    .i0(ins_read[22]),
    .i1(ins_read[54]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [22]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b23  (
    .i0(ins_read[23]),
    .i1(ins_read[55]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [23]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b24  (
    .i0(ins_read[24]),
    .i1(ins_read[56]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [24]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b25  (
    .i0(ins_read[25]),
    .i1(ins_read[57]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [25]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b26  (
    .i0(ins_read[26]),
    .i1(ins_read[58]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [26]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b27  (
    .i0(ins_read[27]),
    .i1(ins_read[59]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [27]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b28  (
    .i0(ins_read[28]),
    .i1(ins_read[60]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [28]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b29  (
    .i0(ins_read[29]),
    .i1(ins_read[61]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [29]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b3  (
    .i0(ins_read[3]),
    .i1(ins_read[35]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [3]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b30  (
    .i0(ins_read[30]),
    .i1(ins_read[62]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [30]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b31  (
    .i0(ins_read[31]),
    .i1(ins_read[63]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [31]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b4  (
    .i0(ins_read[4]),
    .i1(ins_read[36]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [4]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b5  (
    .i0(ins_read[5]),
    .i1(ins_read[37]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [5]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b6  (
    .i0(ins_read[6]),
    .i1(ins_read[38]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [6]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b7  (
    .i0(ins_read[7]),
    .i1(ins_read[39]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [7]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b8  (
    .i0(ins_read[8]),
    .i1(ins_read[40]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [8]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux0_b9  (
    .i0(ins_read[9]),
    .i1(ins_read[41]),
    .sel(id_ins_pc[2]),
    .o(\ins_fetch/ins_shift [9]));  // ../../RTL/CPU/IF/ins_fetch.v(64)
  binary_mux_s1_w1 \ins_fetch/mux2_b10  (
    .i0(\ins_fetch/n3 [8]),
    .i1(flush_pc[10]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [10]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b11  (
    .i0(\ins_fetch/n3 [9]),
    .i1(flush_pc[11]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [11]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b12  (
    .i0(\ins_fetch/n3 [10]),
    .i1(flush_pc[12]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [12]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b13  (
    .i0(\ins_fetch/n3 [11]),
    .i1(flush_pc[13]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [13]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b14  (
    .i0(\ins_fetch/n3 [12]),
    .i1(flush_pc[14]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [14]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b15  (
    .i0(\ins_fetch/n3 [13]),
    .i1(flush_pc[15]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [15]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b16  (
    .i0(\ins_fetch/n3 [14]),
    .i1(flush_pc[16]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [16]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b17  (
    .i0(\ins_fetch/n3 [15]),
    .i1(flush_pc[17]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [17]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b18  (
    .i0(\ins_fetch/n3 [16]),
    .i1(flush_pc[18]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [18]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b19  (
    .i0(\ins_fetch/n3 [17]),
    .i1(flush_pc[19]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [19]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b2  (
    .i0(\ins_fetch/n3 [0]),
    .i1(flush_pc[2]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [2]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b20  (
    .i0(\ins_fetch/n3 [18]),
    .i1(flush_pc[20]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [20]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b21  (
    .i0(\ins_fetch/n3 [19]),
    .i1(flush_pc[21]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [21]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b22  (
    .i0(\ins_fetch/n3 [20]),
    .i1(flush_pc[22]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [22]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b23  (
    .i0(\ins_fetch/n3 [21]),
    .i1(flush_pc[23]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [23]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b24  (
    .i0(\ins_fetch/n3 [22]),
    .i1(flush_pc[24]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [24]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b25  (
    .i0(\ins_fetch/n3 [23]),
    .i1(flush_pc[25]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [25]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b26  (
    .i0(\ins_fetch/n3 [24]),
    .i1(flush_pc[26]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [26]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b27  (
    .i0(\ins_fetch/n3 [25]),
    .i1(flush_pc[27]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [27]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b28  (
    .i0(\ins_fetch/n3 [26]),
    .i1(flush_pc[28]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [28]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b29  (
    .i0(\ins_fetch/n3 [27]),
    .i1(flush_pc[29]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [29]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b3  (
    .i0(\ins_fetch/n3 [1]),
    .i1(flush_pc[3]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [3]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b30  (
    .i0(\ins_fetch/n3 [28]),
    .i1(flush_pc[30]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [30]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b31  (
    .i0(\ins_fetch/n3 [29]),
    .i1(flush_pc[31]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [31]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b32  (
    .i0(\ins_fetch/n3 [30]),
    .i1(flush_pc[32]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [32]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b33  (
    .i0(\ins_fetch/n3 [31]),
    .i1(flush_pc[33]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [33]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b34  (
    .i0(\ins_fetch/n3 [32]),
    .i1(flush_pc[34]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [34]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b35  (
    .i0(\ins_fetch/n3 [33]),
    .i1(flush_pc[35]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [35]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b36  (
    .i0(\ins_fetch/n3 [34]),
    .i1(flush_pc[36]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [36]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b37  (
    .i0(\ins_fetch/n3 [35]),
    .i1(flush_pc[37]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [37]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b38  (
    .i0(\ins_fetch/n3 [36]),
    .i1(flush_pc[38]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [38]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b39  (
    .i0(\ins_fetch/n3 [37]),
    .i1(flush_pc[39]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [39]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b4  (
    .i0(\ins_fetch/n3 [2]),
    .i1(flush_pc[4]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [4]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b40  (
    .i0(\ins_fetch/n3 [38]),
    .i1(flush_pc[40]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [40]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b41  (
    .i0(\ins_fetch/n3 [39]),
    .i1(flush_pc[41]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [41]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b42  (
    .i0(\ins_fetch/n3 [40]),
    .i1(flush_pc[42]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [42]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b43  (
    .i0(\ins_fetch/n3 [41]),
    .i1(flush_pc[43]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [43]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b44  (
    .i0(\ins_fetch/n3 [42]),
    .i1(flush_pc[44]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [44]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b45  (
    .i0(\ins_fetch/n3 [43]),
    .i1(flush_pc[45]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [45]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b46  (
    .i0(\ins_fetch/n3 [44]),
    .i1(flush_pc[46]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [46]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b47  (
    .i0(\ins_fetch/n3 [45]),
    .i1(flush_pc[47]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [47]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b48  (
    .i0(\ins_fetch/n3 [46]),
    .i1(flush_pc[48]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [48]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b49  (
    .i0(\ins_fetch/n3 [47]),
    .i1(flush_pc[49]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [49]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b5  (
    .i0(\ins_fetch/n3 [3]),
    .i1(flush_pc[5]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [5]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b50  (
    .i0(\ins_fetch/n3 [48]),
    .i1(flush_pc[50]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [50]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b51  (
    .i0(\ins_fetch/n3 [49]),
    .i1(flush_pc[51]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [51]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b52  (
    .i0(\ins_fetch/n3 [50]),
    .i1(flush_pc[52]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [52]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b53  (
    .i0(\ins_fetch/n3 [51]),
    .i1(flush_pc[53]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [53]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b54  (
    .i0(\ins_fetch/n3 [52]),
    .i1(flush_pc[54]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [54]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b55  (
    .i0(\ins_fetch/n3 [53]),
    .i1(flush_pc[55]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [55]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b56  (
    .i0(\ins_fetch/n3 [54]),
    .i1(flush_pc[56]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [56]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b57  (
    .i0(\ins_fetch/n3 [55]),
    .i1(flush_pc[57]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [57]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b58  (
    .i0(\ins_fetch/n3 [56]),
    .i1(flush_pc[58]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [58]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b59  (
    .i0(\ins_fetch/n3 [57]),
    .i1(flush_pc[59]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [59]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b6  (
    .i0(\ins_fetch/n3 [4]),
    .i1(flush_pc[6]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [6]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b60  (
    .i0(\ins_fetch/n3 [58]),
    .i1(flush_pc[60]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [60]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b61  (
    .i0(\ins_fetch/n3 [59]),
    .i1(flush_pc[61]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [61]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b62  (
    .i0(\ins_fetch/n3 [60]),
    .i1(flush_pc[62]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [62]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b63  (
    .i0(\ins_fetch/n3 [61]),
    .i1(flush_pc[63]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [63]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b7  (
    .i0(\ins_fetch/n3 [5]),
    .i1(flush_pc[7]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [7]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b8  (
    .i0(\ins_fetch/n3 [6]),
    .i1(flush_pc[8]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [8]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  binary_mux_s1_w1 \ins_fetch/mux2_b9  (
    .i0(\ins_fetch/n3 [7]),
    .i1(flush_pc[9]),
    .sel(pip_flush),
    .o(\ins_fetch/n4 [9]));  // ../../RTL/CPU/IF/ins_fetch.v(82)
  AL_MUX \ins_fetch/mux8_b0  (
    .i0(addr_if[2]),
    .i1(\ins_fetch/n1 [0]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [0]));
  and \ins_fetch/mux8_b0_sel_is_2  (\ins_fetch/mux8_b0_sel_is_2_o , \ins_fetch/n0_neg , cache_ready_if);
  AL_MUX \ins_fetch/mux8_b1  (
    .i0(addr_if[3]),
    .i1(\ins_fetch/n1 [1]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [1]));
  AL_MUX \ins_fetch/mux8_b10  (
    .i0(addr_if[12]),
    .i1(\ins_fetch/n1 [10]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [10]));
  AL_MUX \ins_fetch/mux8_b11  (
    .i0(addr_if[13]),
    .i1(\ins_fetch/n1 [11]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [11]));
  AL_MUX \ins_fetch/mux8_b12  (
    .i0(addr_if[14]),
    .i1(\ins_fetch/n1 [12]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [12]));
  AL_MUX \ins_fetch/mux8_b13  (
    .i0(addr_if[15]),
    .i1(\ins_fetch/n1 [13]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [13]));
  AL_MUX \ins_fetch/mux8_b14  (
    .i0(addr_if[16]),
    .i1(\ins_fetch/n1 [14]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [14]));
  AL_MUX \ins_fetch/mux8_b15  (
    .i0(addr_if[17]),
    .i1(\ins_fetch/n1 [15]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [15]));
  AL_MUX \ins_fetch/mux8_b16  (
    .i0(addr_if[18]),
    .i1(\ins_fetch/n1 [16]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [16]));
  AL_MUX \ins_fetch/mux8_b17  (
    .i0(addr_if[19]),
    .i1(\ins_fetch/n1 [17]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [17]));
  AL_MUX \ins_fetch/mux8_b18  (
    .i0(addr_if[20]),
    .i1(\ins_fetch/n1 [18]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [18]));
  AL_MUX \ins_fetch/mux8_b19  (
    .i0(addr_if[21]),
    .i1(\ins_fetch/n1 [19]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [19]));
  AL_MUX \ins_fetch/mux8_b2  (
    .i0(addr_if[4]),
    .i1(\ins_fetch/n1 [2]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [2]));
  AL_MUX \ins_fetch/mux8_b20  (
    .i0(addr_if[22]),
    .i1(\ins_fetch/n1 [20]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [20]));
  AL_MUX \ins_fetch/mux8_b21  (
    .i0(addr_if[23]),
    .i1(\ins_fetch/n1 [21]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [21]));
  AL_MUX \ins_fetch/mux8_b22  (
    .i0(addr_if[24]),
    .i1(\ins_fetch/n1 [22]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [22]));
  AL_MUX \ins_fetch/mux8_b23  (
    .i0(addr_if[25]),
    .i1(\ins_fetch/n1 [23]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [23]));
  AL_MUX \ins_fetch/mux8_b24  (
    .i0(addr_if[26]),
    .i1(\ins_fetch/n1 [24]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [24]));
  AL_MUX \ins_fetch/mux8_b25  (
    .i0(addr_if[27]),
    .i1(\ins_fetch/n1 [25]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [25]));
  AL_MUX \ins_fetch/mux8_b26  (
    .i0(addr_if[28]),
    .i1(\ins_fetch/n1 [26]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [26]));
  AL_MUX \ins_fetch/mux8_b27  (
    .i0(addr_if[29]),
    .i1(\ins_fetch/n1 [27]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [27]));
  AL_MUX \ins_fetch/mux8_b28  (
    .i0(addr_if[30]),
    .i1(\ins_fetch/n1 [28]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [28]));
  AL_MUX \ins_fetch/mux8_b29  (
    .i0(addr_if[31]),
    .i1(\ins_fetch/n1 [29]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [29]));
  AL_MUX \ins_fetch/mux8_b3  (
    .i0(addr_if[5]),
    .i1(\ins_fetch/n1 [3]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [3]));
  AL_MUX \ins_fetch/mux8_b30  (
    .i0(addr_if[32]),
    .i1(\ins_fetch/n1 [30]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [30]));
  AL_MUX \ins_fetch/mux8_b31  (
    .i0(addr_if[33]),
    .i1(\ins_fetch/n1 [31]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [31]));
  AL_MUX \ins_fetch/mux8_b32  (
    .i0(addr_if[34]),
    .i1(\ins_fetch/n1 [32]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [32]));
  AL_MUX \ins_fetch/mux8_b33  (
    .i0(addr_if[35]),
    .i1(\ins_fetch/n1 [33]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [33]));
  AL_MUX \ins_fetch/mux8_b34  (
    .i0(addr_if[36]),
    .i1(\ins_fetch/n1 [34]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [34]));
  AL_MUX \ins_fetch/mux8_b35  (
    .i0(addr_if[37]),
    .i1(\ins_fetch/n1 [35]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [35]));
  AL_MUX \ins_fetch/mux8_b36  (
    .i0(addr_if[38]),
    .i1(\ins_fetch/n1 [36]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [36]));
  AL_MUX \ins_fetch/mux8_b37  (
    .i0(addr_if[39]),
    .i1(\ins_fetch/n1 [37]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [37]));
  AL_MUX \ins_fetch/mux8_b38  (
    .i0(addr_if[40]),
    .i1(\ins_fetch/n1 [38]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [38]));
  AL_MUX \ins_fetch/mux8_b39  (
    .i0(addr_if[41]),
    .i1(\ins_fetch/n1 [39]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [39]));
  AL_MUX \ins_fetch/mux8_b4  (
    .i0(addr_if[6]),
    .i1(\ins_fetch/n1 [4]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [4]));
  AL_MUX \ins_fetch/mux8_b40  (
    .i0(addr_if[42]),
    .i1(\ins_fetch/n1 [40]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [40]));
  AL_MUX \ins_fetch/mux8_b41  (
    .i0(addr_if[43]),
    .i1(\ins_fetch/n1 [41]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [41]));
  AL_MUX \ins_fetch/mux8_b42  (
    .i0(addr_if[44]),
    .i1(\ins_fetch/n1 [42]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [42]));
  AL_MUX \ins_fetch/mux8_b43  (
    .i0(addr_if[45]),
    .i1(\ins_fetch/n1 [43]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [43]));
  AL_MUX \ins_fetch/mux8_b44  (
    .i0(addr_if[46]),
    .i1(\ins_fetch/n1 [44]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [44]));
  AL_MUX \ins_fetch/mux8_b45  (
    .i0(addr_if[47]),
    .i1(\ins_fetch/n1 [45]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [45]));
  AL_MUX \ins_fetch/mux8_b46  (
    .i0(addr_if[48]),
    .i1(\ins_fetch/n1 [46]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [46]));
  AL_MUX \ins_fetch/mux8_b47  (
    .i0(addr_if[49]),
    .i1(\ins_fetch/n1 [47]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [47]));
  AL_MUX \ins_fetch/mux8_b48  (
    .i0(addr_if[50]),
    .i1(\ins_fetch/n1 [48]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [48]));
  AL_MUX \ins_fetch/mux8_b49  (
    .i0(addr_if[51]),
    .i1(\ins_fetch/n1 [49]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [49]));
  AL_MUX \ins_fetch/mux8_b5  (
    .i0(addr_if[7]),
    .i1(\ins_fetch/n1 [5]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [5]));
  AL_MUX \ins_fetch/mux8_b50  (
    .i0(addr_if[52]),
    .i1(\ins_fetch/n1 [50]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [50]));
  AL_MUX \ins_fetch/mux8_b51  (
    .i0(addr_if[53]),
    .i1(\ins_fetch/n1 [51]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [51]));
  AL_MUX \ins_fetch/mux8_b52  (
    .i0(addr_if[54]),
    .i1(\ins_fetch/n1 [52]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [52]));
  AL_MUX \ins_fetch/mux8_b53  (
    .i0(addr_if[55]),
    .i1(\ins_fetch/n1 [53]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [53]));
  AL_MUX \ins_fetch/mux8_b54  (
    .i0(addr_if[56]),
    .i1(\ins_fetch/n1 [54]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [54]));
  AL_MUX \ins_fetch/mux8_b55  (
    .i0(addr_if[57]),
    .i1(\ins_fetch/n1 [55]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [55]));
  AL_MUX \ins_fetch/mux8_b56  (
    .i0(addr_if[58]),
    .i1(\ins_fetch/n1 [56]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [56]));
  AL_MUX \ins_fetch/mux8_b57  (
    .i0(addr_if[59]),
    .i1(\ins_fetch/n1 [57]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [57]));
  AL_MUX \ins_fetch/mux8_b58  (
    .i0(addr_if[60]),
    .i1(\ins_fetch/n1 [58]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [58]));
  AL_MUX \ins_fetch/mux8_b59  (
    .i0(addr_if[61]),
    .i1(\ins_fetch/n1 [59]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [59]));
  AL_MUX \ins_fetch/mux8_b6  (
    .i0(addr_if[8]),
    .i1(\ins_fetch/n1 [6]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [6]));
  AL_MUX \ins_fetch/mux8_b60  (
    .i0(addr_if[62]),
    .i1(\ins_fetch/n1 [60]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [60]));
  AL_MUX \ins_fetch/mux8_b61  (
    .i0(addr_if[63]),
    .i1(\ins_fetch/n1 [61]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [61]));
  AL_MUX \ins_fetch/mux8_b7  (
    .i0(addr_if[9]),
    .i1(\ins_fetch/n1 [7]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [7]));
  AL_MUX \ins_fetch/mux8_b8  (
    .i0(addr_if[10]),
    .i1(\ins_fetch/n1 [8]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [8]));
  AL_MUX \ins_fetch/mux8_b9  (
    .i0(addr_if[11]),
    .i1(\ins_fetch/n1 [9]),
    .sel(\ins_fetch/mux8_b0_sel_is_2_o ),
    .o(\ins_fetch/n3 [9]));
  binary_mux_s1_w1 \ins_fetch/mux9_b0  (
    .i0(\ins_fetch/ins_shift [0]),
    .i1(\ins_fetch/ins_hold [0]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[0]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b1  (
    .i0(\ins_fetch/ins_shift [1]),
    .i1(\ins_fetch/ins_hold [1]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[1]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b10  (
    .i0(\ins_fetch/ins_shift [10]),
    .i1(\ins_fetch/ins_hold [10]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[10]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b11  (
    .i0(\ins_fetch/ins_shift [11]),
    .i1(\ins_fetch/ins_hold [11]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[11]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b12  (
    .i0(\ins_fetch/ins_shift [12]),
    .i1(\ins_fetch/ins_hold [12]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[12]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b13  (
    .i0(\ins_fetch/ins_shift [13]),
    .i1(\ins_fetch/ins_hold [13]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[13]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b14  (
    .i0(\ins_fetch/ins_shift [14]),
    .i1(\ins_fetch/ins_hold [14]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[14]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b15  (
    .i0(\ins_fetch/ins_shift [15]),
    .i1(\ins_fetch/ins_hold [15]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[15]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b16  (
    .i0(\ins_fetch/ins_shift [16]),
    .i1(\ins_fetch/ins_hold [16]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[16]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b17  (
    .i0(\ins_fetch/ins_shift [17]),
    .i1(\ins_fetch/ins_hold [17]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[17]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b18  (
    .i0(\ins_fetch/ins_shift [18]),
    .i1(\ins_fetch/ins_hold [18]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[18]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b19  (
    .i0(\ins_fetch/ins_shift [19]),
    .i1(\ins_fetch/ins_hold [19]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[19]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b2  (
    .i0(\ins_fetch/ins_shift [2]),
    .i1(\ins_fetch/ins_hold [2]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[2]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b20  (
    .i0(\ins_fetch/ins_shift [20]),
    .i1(\ins_fetch/ins_hold [20]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[20]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b21  (
    .i0(\ins_fetch/ins_shift [21]),
    .i1(\ins_fetch/ins_hold [21]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[21]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b22  (
    .i0(\ins_fetch/ins_shift [22]),
    .i1(\ins_fetch/ins_hold [22]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[22]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b23  (
    .i0(\ins_fetch/ins_shift [23]),
    .i1(\ins_fetch/ins_hold [23]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[23]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b24  (
    .i0(\ins_fetch/ins_shift [24]),
    .i1(\ins_fetch/ins_hold [24]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[24]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b25  (
    .i0(\ins_fetch/ins_shift [25]),
    .i1(\ins_fetch/ins_hold [25]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[25]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b26  (
    .i0(\ins_fetch/ins_shift [26]),
    .i1(\ins_fetch/ins_hold [26]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[26]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b27  (
    .i0(\ins_fetch/ins_shift [27]),
    .i1(\ins_fetch/ins_hold [27]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[27]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b28  (
    .i0(\ins_fetch/ins_shift [28]),
    .i1(\ins_fetch/ins_hold [28]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[28]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b29  (
    .i0(\ins_fetch/ins_shift [29]),
    .i1(\ins_fetch/ins_hold [29]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[29]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b3  (
    .i0(\ins_fetch/ins_shift [3]),
    .i1(\ins_fetch/ins_hold [3]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[3]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b30  (
    .i0(\ins_fetch/ins_shift [30]),
    .i1(\ins_fetch/ins_hold [30]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[30]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b31  (
    .i0(\ins_fetch/ins_shift [31]),
    .i1(\ins_fetch/ins_hold [31]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[31]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b4  (
    .i0(\ins_fetch/ins_shift [4]),
    .i1(\ins_fetch/ins_hold [4]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[4]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b5  (
    .i0(\ins_fetch/ins_shift [5]),
    .i1(\ins_fetch/ins_hold [5]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[5]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b6  (
    .i0(\ins_fetch/ins_shift [6]),
    .i1(\ins_fetch/ins_hold [6]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[6]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b7  (
    .i0(\ins_fetch/ins_shift [7]),
    .i1(\ins_fetch/ins_hold [7]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[7]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b8  (
    .i0(\ins_fetch/ins_shift [8]),
    .i1(\ins_fetch/ins_hold [8]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[8]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  binary_mux_s1_w1 \ins_fetch/mux9_b9  (
    .i0(\ins_fetch/ins_shift [9]),
    .i1(\ins_fetch/ins_hold [9]),
    .sel(\ins_fetch/hold ),
    .o(id_ins[9]));  // ../../RTL/CPU/IF/ins_fetch.v(156)
  not \ins_fetch/n0_inv  (\ins_fetch/n0_neg , \ins_fetch/n0 );
  ne_w2 \ins_fetch/neq0  (
    .i0(addr_if[1:0]),
    .i1(2'b00),
    .o(\ins_fetch/addr_mis ));  // ../../RTL/CPU/IF/ins_fetch.v(62)
  reg_sr_as_w1 \ins_fetch/reg0_b0  (
    .clk(clk),
    .d(addr_if[0]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[0]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b1  (
    .clk(clk),
    .d(addr_if[1]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[1]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b10  (
    .clk(clk),
    .d(addr_if[10]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[10]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b11  (
    .clk(clk),
    .d(addr_if[11]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[11]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b12  (
    .clk(clk),
    .d(addr_if[12]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[12]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b13  (
    .clk(clk),
    .d(addr_if[13]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[13]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b14  (
    .clk(clk),
    .d(addr_if[14]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[14]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b15  (
    .clk(clk),
    .d(addr_if[15]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[15]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b16  (
    .clk(clk),
    .d(addr_if[16]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[16]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b17  (
    .clk(clk),
    .d(addr_if[17]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[17]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b18  (
    .clk(clk),
    .d(addr_if[18]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[18]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b19  (
    .clk(clk),
    .d(addr_if[19]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[19]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b2  (
    .clk(clk),
    .d(addr_if[2]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[2]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b20  (
    .clk(clk),
    .d(addr_if[20]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[20]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b21  (
    .clk(clk),
    .d(addr_if[21]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[21]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b22  (
    .clk(clk),
    .d(addr_if[22]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[22]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b23  (
    .clk(clk),
    .d(addr_if[23]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[23]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b24  (
    .clk(clk),
    .d(addr_if[24]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[24]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b25  (
    .clk(clk),
    .d(addr_if[25]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[25]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b26  (
    .clk(clk),
    .d(addr_if[26]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[26]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b27  (
    .clk(clk),
    .d(addr_if[27]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[27]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b28  (
    .clk(clk),
    .d(addr_if[28]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[28]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b29  (
    .clk(clk),
    .d(addr_if[29]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[29]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b3  (
    .clk(clk),
    .d(addr_if[3]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[3]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b30  (
    .clk(clk),
    .d(addr_if[30]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[30]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b31  (
    .clk(clk),
    .d(addr_if[31]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[31]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b32  (
    .clk(clk),
    .d(addr_if[32]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[32]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b33  (
    .clk(clk),
    .d(addr_if[33]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[33]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b34  (
    .clk(clk),
    .d(addr_if[34]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[34]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b35  (
    .clk(clk),
    .d(addr_if[35]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[35]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b36  (
    .clk(clk),
    .d(addr_if[36]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[36]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b37  (
    .clk(clk),
    .d(addr_if[37]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[37]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b38  (
    .clk(clk),
    .d(addr_if[38]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[38]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b39  (
    .clk(clk),
    .d(addr_if[39]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[39]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b4  (
    .clk(clk),
    .d(addr_if[4]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[4]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b40  (
    .clk(clk),
    .d(addr_if[40]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[40]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b41  (
    .clk(clk),
    .d(addr_if[41]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[41]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b42  (
    .clk(clk),
    .d(addr_if[42]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[42]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b43  (
    .clk(clk),
    .d(addr_if[43]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[43]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b44  (
    .clk(clk),
    .d(addr_if[44]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[44]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b45  (
    .clk(clk),
    .d(addr_if[45]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[45]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b46  (
    .clk(clk),
    .d(addr_if[46]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[46]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b47  (
    .clk(clk),
    .d(addr_if[47]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[47]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b48  (
    .clk(clk),
    .d(addr_if[48]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[48]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b49  (
    .clk(clk),
    .d(addr_if[49]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[49]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b5  (
    .clk(clk),
    .d(addr_if[5]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[5]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b50  (
    .clk(clk),
    .d(addr_if[50]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[50]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b51  (
    .clk(clk),
    .d(addr_if[51]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[51]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b52  (
    .clk(clk),
    .d(addr_if[52]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[52]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b53  (
    .clk(clk),
    .d(addr_if[53]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[53]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b54  (
    .clk(clk),
    .d(addr_if[54]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[54]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b55  (
    .clk(clk),
    .d(addr_if[55]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[55]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b56  (
    .clk(clk),
    .d(addr_if[56]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[56]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b57  (
    .clk(clk),
    .d(addr_if[57]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[57]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b58  (
    .clk(clk),
    .d(addr_if[58]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[58]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b59  (
    .clk(clk),
    .d(addr_if[59]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[59]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b6  (
    .clk(clk),
    .d(addr_if[6]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[6]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b60  (
    .clk(clk),
    .d(addr_if[60]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[60]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b61  (
    .clk(clk),
    .d(addr_if[61]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[61]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b62  (
    .clk(clk),
    .d(addr_if[62]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[62]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b63  (
    .clk(clk),
    .d(addr_if[63]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[63]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b7  (
    .clk(clk),
    .d(addr_if[7]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[7]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b8  (
    .clk(clk),
    .d(addr_if[8]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[8]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg0_b9  (
    .clk(clk),
    .d(addr_if[9]),
    .en(~if_hold),
    .reset(rst),
    .set(1'b0),
    .q(id_ins_pc[9]));  // ../../RTL/CPU/IF/ins_fetch.v(95)
  reg_sr_as_w1 \ins_fetch/reg1_b0  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [0]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [0]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b1  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [1]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [1]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b10  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [10]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [10]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b11  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [11]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [11]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b12  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [12]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [12]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b13  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [13]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [13]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b14  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [14]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [14]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b15  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [15]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [15]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b16  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [16]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [16]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b17  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [17]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [17]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b18  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [18]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [18]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b19  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [19]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [19]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b2  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [2]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [2]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b20  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [20]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [20]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b21  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [21]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [21]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b22  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [22]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [22]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b23  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [23]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [23]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b24  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [24]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [24]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b25  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [25]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [25]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b26  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [26]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [26]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b27  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [27]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [27]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b28  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [28]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [28]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b29  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [29]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [29]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b3  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [3]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [3]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b30  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [30]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [30]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b31  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [31]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [31]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b4  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [4]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [4]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b5  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [5]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [5]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b6  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [6]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [6]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b7  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [7]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [7]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b8  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [8]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [8]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg1_b9  (
    .clk(clk),
    .d(\ins_fetch/ins_shift [9]),
    .en(\ins_fetch/n9 ),
    .reset(rst),
    .set(1'b0),
    .q(\ins_fetch/ins_hold [9]));  // ../../RTL/CPU/IF/ins_fetch.v(104)
  reg_sr_as_w1 \ins_fetch/reg2_b0  (
    .clk(clk),
    .d(flush_pc[0]),
    .en(pip_flush),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[0]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b1  (
    .clk(clk),
    .d(flush_pc[1]),
    .en(pip_flush),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[1]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b10  (
    .clk(clk),
    .d(\ins_fetch/n4 [10]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[10]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b11  (
    .clk(clk),
    .d(\ins_fetch/n4 [11]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[11]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b12  (
    .clk(clk),
    .d(\ins_fetch/n4 [12]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[12]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b13  (
    .clk(clk),
    .d(\ins_fetch/n4 [13]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[13]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b14  (
    .clk(clk),
    .d(\ins_fetch/n4 [14]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[14]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b15  (
    .clk(clk),
    .d(\ins_fetch/n4 [15]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[15]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b16  (
    .clk(clk),
    .d(\ins_fetch/n4 [16]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[16]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b17  (
    .clk(clk),
    .d(\ins_fetch/n4 [17]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[17]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b18  (
    .clk(clk),
    .d(\ins_fetch/n4 [18]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[18]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b19  (
    .clk(clk),
    .d(\ins_fetch/n4 [19]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[19]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b2  (
    .clk(clk),
    .d(\ins_fetch/n4 [2]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[2]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b20  (
    .clk(clk),
    .d(\ins_fetch/n4 [20]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[20]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b21  (
    .clk(clk),
    .d(\ins_fetch/n4 [21]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[21]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b22  (
    .clk(clk),
    .d(\ins_fetch/n4 [22]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[22]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b23  (
    .clk(clk),
    .d(\ins_fetch/n4 [23]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[23]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b24  (
    .clk(clk),
    .d(\ins_fetch/n4 [24]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[24]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b25  (
    .clk(clk),
    .d(\ins_fetch/n4 [25]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[25]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b26  (
    .clk(clk),
    .d(\ins_fetch/n4 [26]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[26]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b27  (
    .clk(clk),
    .d(\ins_fetch/n4 [27]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[27]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b28  (
    .clk(clk),
    .d(\ins_fetch/n4 [28]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[28]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b29  (
    .clk(clk),
    .d(\ins_fetch/n4 [29]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[29]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b3  (
    .clk(clk),
    .d(\ins_fetch/n4 [3]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[3]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b30  (
    .clk(clk),
    .d(\ins_fetch/n4 [30]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[30]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b31  (
    .clk(clk),
    .d(\ins_fetch/n4 [31]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[31]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b32  (
    .clk(clk),
    .d(\ins_fetch/n4 [32]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[32]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b33  (
    .clk(clk),
    .d(\ins_fetch/n4 [33]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[33]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b34  (
    .clk(clk),
    .d(\ins_fetch/n4 [34]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[34]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b35  (
    .clk(clk),
    .d(\ins_fetch/n4 [35]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[35]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b36  (
    .clk(clk),
    .d(\ins_fetch/n4 [36]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[36]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b37  (
    .clk(clk),
    .d(\ins_fetch/n4 [37]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[37]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b38  (
    .clk(clk),
    .d(\ins_fetch/n4 [38]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[38]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b39  (
    .clk(clk),
    .d(\ins_fetch/n4 [39]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[39]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b4  (
    .clk(clk),
    .d(\ins_fetch/n4 [4]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[4]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b40  (
    .clk(clk),
    .d(\ins_fetch/n4 [40]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[40]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b41  (
    .clk(clk),
    .d(\ins_fetch/n4 [41]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[41]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b42  (
    .clk(clk),
    .d(\ins_fetch/n4 [42]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[42]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b43  (
    .clk(clk),
    .d(\ins_fetch/n4 [43]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[43]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b44  (
    .clk(clk),
    .d(\ins_fetch/n4 [44]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[44]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b45  (
    .clk(clk),
    .d(\ins_fetch/n4 [45]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[45]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b46  (
    .clk(clk),
    .d(\ins_fetch/n4 [46]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[46]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b47  (
    .clk(clk),
    .d(\ins_fetch/n4 [47]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[47]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b48  (
    .clk(clk),
    .d(\ins_fetch/n4 [48]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[48]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b49  (
    .clk(clk),
    .d(\ins_fetch/n4 [49]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[49]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b5  (
    .clk(clk),
    .d(\ins_fetch/n4 [5]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[5]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b50  (
    .clk(clk),
    .d(\ins_fetch/n4 [50]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[50]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b51  (
    .clk(clk),
    .d(\ins_fetch/n4 [51]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[51]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b52  (
    .clk(clk),
    .d(\ins_fetch/n4 [52]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[52]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b53  (
    .clk(clk),
    .d(\ins_fetch/n4 [53]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[53]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b54  (
    .clk(clk),
    .d(\ins_fetch/n4 [54]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[54]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b55  (
    .clk(clk),
    .d(\ins_fetch/n4 [55]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[55]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b56  (
    .clk(clk),
    .d(\ins_fetch/n4 [56]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[56]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b57  (
    .clk(clk),
    .d(\ins_fetch/n4 [57]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[57]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b58  (
    .clk(clk),
    .d(\ins_fetch/n4 [58]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[58]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b59  (
    .clk(clk),
    .d(\ins_fetch/n4 [59]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[59]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b6  (
    .clk(clk),
    .d(\ins_fetch/n4 [6]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[6]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b60  (
    .clk(clk),
    .d(\ins_fetch/n4 [60]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[60]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b61  (
    .clk(clk),
    .d(\ins_fetch/n4 [61]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[61]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b62  (
    .clk(clk),
    .d(\ins_fetch/n4 [62]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[62]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b63  (
    .clk(clk),
    .d(\ins_fetch/n4 [63]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[63]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b7  (
    .clk(clk),
    .d(\ins_fetch/n4 [7]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[7]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b8  (
    .clk(clk),
    .d(\ins_fetch/n4 [8]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[8]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  reg_sr_as_w1 \ins_fetch/reg2_b9  (
    .clk(clk),
    .d(\ins_fetch/n4 [9]),
    .en(1'b1),
    .reset(rst),
    .set(1'b0),
    .q(addr_if[9]));  // ../../RTL/CPU/IF/ins_fetch.v(83)
  or \ins_fetch/u4  (\ins_fetch/n0 , if_nop, if_hold);  // ../../RTL/CPU/IF/ins_fetch.v(77)
  and \ins_fetch/u67  (\ins_fetch/n9 , if_hold, \ins_fetch/hold_neg );  // ../../RTL/CPU/IF/ins_fetch.v(101)
  and \ins_fetch/u72_sel_is_1  (\ins_fetch/u72_sel_is_1_o , \ins_fetch/hold , \ins_fetch/hold_neg );
  or \ins_fetch/u82  (\ins_fetch/n23 , rst, id_ins_acc_fault);  // ../../RTL/CPU/IF/ins_fetch.v(142)
  or \ins_fetch/u83  (\ins_fetch/n24 , \ins_fetch/n23 , id_ins_page_fault);  // ../../RTL/CPU/IF/ins_fetch.v(142)
  or \ins_fetch/u84  (\ins_fetch/n25 , \ins_fetch/n24 , id_ins_addr_mis);  // ../../RTL/CPU/IF/ins_fetch.v(142)
  not \ins_fetch/u85  (\ins_fetch/n26 , if_nop);  // ../../RTL/CPU/IF/ins_fetch.v(145)
  and \ins_fetch/u86  (\ins_fetch/n27 , cache_ready_if, \ins_fetch/n26 );  // ../../RTL/CPU/IF/ins_fetch.v(145)
  not \ins_fetch/u92  (\ins_fetch/n31 , if_hold);  // ../../RTL/CPU/IF/ins_fetch.v(159)
  and \ins_fetch/u93  (rd_ins, \ins_fetch/n26 , \ins_fetch/n31 );  // ../../RTL/CPU/IF/ins_fetch.v(159)
  reg_sr_ss_w1 \ins_fetch/valid_reg  (
    .clk(clk),
    .d(1'b0),
    .en(~if_hold),
    .reset(\ins_fetch/n25 ),
    .set(\ins_fetch/n27 ),
    .q(id_valid));  // ../../RTL/CPU/IF/ins_fetch.v(154)
  not load_acc_fault_inv (load_acc_fault_neg, load_acc_fault);
  not load_inv (load_neg, load);
  eq_w5 \pip_ctrl/eq0  (
    .i0(id_rs1_index),
    .i1(ex_rd_index),
    .o(\pip_ctrl/n36 ));  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(96)
  eq_w5 \pip_ctrl/eq1  (
    .i0(id_rs2_index),
    .i1(ex_rd_index),
    .o(\pip_ctrl/n42 ));  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(97)
  eq_w5 \pip_ctrl/eq2  (
    .i0(id_rs1_index),
    .i1(wb_rd_index),
    .o(\pip_ctrl/n46 ));  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(100)
  eq_w5 \pip_ctrl/eq3  (
    .i0(id_rs2_index),
    .i1(wb_rd_index),
    .o(\pip_ctrl/n50 ));  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(101)
  ne_w5 \pip_ctrl/neq0  (
    .i0(id_rs1_index),
    .i1(5'b00000),
    .o(\pip_ctrl/n33 ));  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(96)
  ne_w5 \pip_ctrl/neq1  (
    .i0(id_rs2_index),
    .i1(5'b00000),
    .o(\pip_ctrl/n39 ));  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(97)
  or \pip_ctrl/u1  (\pip_ctrl/n0 , id_ill_ins, id_system);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(86)
  or \pip_ctrl/u10  (\pip_ctrl/n8 , \pip_ctrl/n7 , ex_ins_acc_fault);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(88)
  or \pip_ctrl/u11  (\pip_ctrl/n9 , \pip_ctrl/n8 , ex_ins_addr_mis);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(88)
  or \pip_ctrl/u12  (\pip_ctrl/n10 , \pip_ctrl/n9 , ex_ins_page_fault);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(88)
  or \pip_ctrl/u13  (\pip_ctrl/n11 , \pip_ctrl/n10 , ex_int_acc);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(89)
  or \pip_ctrl/u14  (\pip_ctrl/n12 , \pip_ctrl/n11 , ex_ill_ins);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(89)
  or \pip_ctrl/u15  (\pip_ctrl/n13 , \pip_ctrl/n12 , ex_m_ret);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(89)
  or \pip_ctrl/u16  (\pip_ctrl/n14 , \pip_ctrl/n13 , ex_s_ret);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(89)
  or \pip_ctrl/u17  (\pip_ctrl/n15 , \pip_ctrl/n14 , ex_ecall);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(89)
  or \pip_ctrl/u18  (\pip_ctrl/n16 , \pip_ctrl/n15 , ex_ebreak);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(89)
  and \pip_ctrl/u19  (\pip_ctrl/ex_exception , ex_valid, \pip_ctrl/n16 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(89)
  or \pip_ctrl/u2  (\pip_ctrl/n1 , \pip_ctrl/n0 , id_branch);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(86)
  or \pip_ctrl/u20  (\pip_ctrl/n17 , wb_system, wb_jmp);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(90)
  or \pip_ctrl/u21  (\pip_ctrl/n18 , \pip_ctrl/n17 , wb_ins_acc_fault);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(90)
  or \pip_ctrl/u22  (\pip_ctrl/n19 , \pip_ctrl/n18 , wb_ins_addr_mis);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(90)
  or \pip_ctrl/u23  (\pip_ctrl/n20 , \pip_ctrl/n19 , wb_ins_page_fault);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(90)
  or \pip_ctrl/u24  (\pip_ctrl/n21 , \pip_ctrl/n20 , wb_ld_addr_mis);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(90)
  or \pip_ctrl/u25  (\pip_ctrl/n22 , \pip_ctrl/n21 , wb_st_addr_mis);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(91)
  or \pip_ctrl/u26  (\pip_ctrl/n23 , \pip_ctrl/n22 , wb_ld_acc_fault);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(91)
  or \pip_ctrl/u27  (\pip_ctrl/n24 , \pip_ctrl/n23 , wb_st_acc_fault);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(91)
  or \pip_ctrl/u28  (\pip_ctrl/n25 , \pip_ctrl/n24 , wb_ld_page_fault);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(91)
  or \pip_ctrl/u29  (\pip_ctrl/n26 , \pip_ctrl/n25 , wb_st_page_fault);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(91)
  or \pip_ctrl/u3  (\pip_ctrl/n2 , \pip_ctrl/n1 , id_ins_acc_fault);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(86)
  or \pip_ctrl/u30  (\pip_ctrl/n27 , \pip_ctrl/n26 , wb_int_acc);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(91)
  or \pip_ctrl/u31  (\pip_ctrl/n28 , \pip_ctrl/n27 , wb_ill_ins);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(91)
  or \pip_ctrl/u32  (\pip_ctrl/n29 , \pip_ctrl/n28 , wb_m_ret);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(92)
  or \pip_ctrl/u33  (\pip_ctrl/n30 , \pip_ctrl/n29 , wb_s_ret);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(92)
  or \pip_ctrl/u34  (\pip_ctrl/n31 , \pip_ctrl/n30 , wb_ecall);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(92)
  or \pip_ctrl/u35  (\pip_ctrl/n32 , \pip_ctrl/n31 , wb_ebreak);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(92)
  and \pip_ctrl/u36  (ex_nop, wb_valid, \pip_ctrl/n32 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(92)
  and \pip_ctrl/u37  (\pip_ctrl/n34 , id_valid, \pip_ctrl/n33 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(96)
  and \pip_ctrl/u38  (\pip_ctrl/n35 , \pip_ctrl/n34 , ex_valid);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(96)
  and \pip_ctrl/u39  (\pip_ctrl/n37 , \pip_ctrl/n35 , \pip_ctrl/n36 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(96)
  or \pip_ctrl/u4  (\pip_ctrl/n3 , \pip_ctrl/n2 , id_ins_addr_mis);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(86)
  and \pip_ctrl/u40  (\pip_ctrl/n38 , \pip_ctrl/n37 , ex_gpr_write);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(96)
  and \pip_ctrl/u41  (\pip_ctrl/n40 , id_valid, \pip_ctrl/n39 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(97)
  and \pip_ctrl/u42  (\pip_ctrl/n41 , \pip_ctrl/n40 , ex_valid);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(97)
  and \pip_ctrl/u43  (\pip_ctrl/n43 , \pip_ctrl/n41 , \pip_ctrl/n42 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(97)
  and \pip_ctrl/u44  (\pip_ctrl/n44 , \pip_ctrl/n43 , ex_gpr_write);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(97)
  or \pip_ctrl/u45  (\pip_ctrl/id_ex_war , \pip_ctrl/n38 , \pip_ctrl/n44 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(97)
  and \pip_ctrl/u46  (\pip_ctrl/n45 , \pip_ctrl/n34 , wb_valid);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(100)
  and \pip_ctrl/u47  (\pip_ctrl/n47 , \pip_ctrl/n45 , \pip_ctrl/n46 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(100)
  and \pip_ctrl/u48  (\pip_ctrl/n48 , \pip_ctrl/n47 , wb_gpr_write);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(100)
  and \pip_ctrl/u49  (\pip_ctrl/n49 , \pip_ctrl/n40 , wb_valid);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(101)
  or \pip_ctrl/u5  (\pip_ctrl/n4 , \pip_ctrl/n3 , id_ins_page_fault);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(86)
  and \pip_ctrl/u50  (\pip_ctrl/n51 , \pip_ctrl/n49 , \pip_ctrl/n50 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(101)
  and \pip_ctrl/u51  (\pip_ctrl/n52 , \pip_ctrl/n51 , wb_gpr_write);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(101)
  or \pip_ctrl/u52  (\pip_ctrl/id_wb_war , \pip_ctrl/n48 , \pip_ctrl/n52 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(101)
  or \pip_ctrl/u53  (\pip_ctrl/n53 , \pip_ctrl/id_exception , \pip_ctrl/ex_exception );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(105)
  or \pip_ctrl/u54  (if_nop, \pip_ctrl/n53 , ex_nop);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(105)
  or \pip_ctrl/u56  (\pip_ctrl/n55 , \pip_ctrl/id_ex_war , \pip_ctrl/id_wb_war );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(109)
  not \pip_ctrl/u57  (\pip_ctrl/n56 , ex_ready);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(109)
  or \pip_ctrl/u58  (\pip_ctrl/n57 , \pip_ctrl/n55 , \pip_ctrl/n56 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(109)
  and \pip_ctrl/u59  (if_hold, \ins_fetch/n26 , \pip_ctrl/n57 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(109)
  or \pip_ctrl/u6  (\pip_ctrl/n5 , \pip_ctrl/n4 , id_int_acc);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(86)
  or \pip_ctrl/u60  (\pip_ctrl/n58 , \pip_ctrl/ex_exception , ex_nop);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(112)
  or \pip_ctrl/u61  (\pip_ctrl/n59 , \pip_ctrl/n58 , \pip_ctrl/id_ex_war );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(112)
  or \pip_ctrl/u62  (id_nop, \pip_ctrl/n59 , \pip_ctrl/id_wb_war );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(112)
  and \pip_ctrl/u64  (id_hold, id_nop_neg, \pip_ctrl/n56 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(114)
  and \pip_ctrl/u7  (\pip_ctrl/id_exception , id_valid, \pip_ctrl/n5 );  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(86)
  or \pip_ctrl/u8  (\pip_ctrl/n6 , ex_more_exception, ex_system);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(88)
  or \pip_ctrl/u9  (\pip_ctrl/n7 , \pip_ctrl/n6 , ex_jmp);  // ../../RTL/CPU/PIP_CTRL/pip_ctrl.v(88)
  not \priv[1]_inv  (\priv[1]_neg , priv[1]);
  not \priv[3]_inv  (\priv[3]_neg , priv[3]);
  not rst_inv (rst_neg, rst);
  not store_acc_fault_inv (store_acc_fault_neg, store_acc_fault);
  not store_inv (store_neg, store);

endmodule 

module add_pu9_pu9_o9
  (
  i0,
  i1,
  o
  );

  input [8:0] i0;
  input [8:0] i1;
  output [8:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;

  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));

endmodule 

module add_pu61_pu61_o61
  (
  i0,
  i1,
  o
  );

  input [60:0] i0;
  input [60:0] i1;
  output [60:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a32;
  wire net_a33;
  wire net_a34;
  wire net_a35;
  wire net_a36;
  wire net_a37;
  wire net_a38;
  wire net_a39;
  wire net_a4;
  wire net_a40;
  wire net_a41;
  wire net_a42;
  wire net_a43;
  wire net_a44;
  wire net_a45;
  wire net_a46;
  wire net_a47;
  wire net_a48;
  wire net_a49;
  wire net_a5;
  wire net_a50;
  wire net_a51;
  wire net_a52;
  wire net_a53;
  wire net_a54;
  wire net_a55;
  wire net_a56;
  wire net_a57;
  wire net_a58;
  wire net_a59;
  wire net_a6;
  wire net_a60;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b32;
  wire net_b33;
  wire net_b34;
  wire net_b35;
  wire net_b36;
  wire net_b37;
  wire net_b38;
  wire net_b39;
  wire net_b4;
  wire net_b40;
  wire net_b41;
  wire net_b42;
  wire net_b43;
  wire net_b44;
  wire net_b45;
  wire net_b46;
  wire net_b47;
  wire net_b48;
  wire net_b49;
  wire net_b5;
  wire net_b50;
  wire net_b51;
  wire net_b52;
  wire net_b53;
  wire net_b54;
  wire net_b55;
  wire net_b56;
  wire net_b57;
  wire net_b58;
  wire net_b59;
  wire net_b6;
  wire net_b60;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout32;
  wire net_cout33;
  wire net_cout34;
  wire net_cout35;
  wire net_cout36;
  wire net_cout37;
  wire net_cout38;
  wire net_cout39;
  wire net_cout4;
  wire net_cout40;
  wire net_cout41;
  wire net_cout42;
  wire net_cout43;
  wire net_cout44;
  wire net_cout45;
  wire net_cout46;
  wire net_cout47;
  wire net_cout48;
  wire net_cout49;
  wire net_cout5;
  wire net_cout50;
  wire net_cout51;
  wire net_cout52;
  wire net_cout53;
  wire net_cout54;
  wire net_cout55;
  wire net_cout56;
  wire net_cout57;
  wire net_cout58;
  wire net_cout59;
  wire net_cout6;
  wire net_cout60;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum32;
  wire net_sum33;
  wire net_sum34;
  wire net_sum35;
  wire net_sum36;
  wire net_sum37;
  wire net_sum38;
  wire net_sum39;
  wire net_sum4;
  wire net_sum40;
  wire net_sum41;
  wire net_sum42;
  wire net_sum43;
  wire net_sum44;
  wire net_sum45;
  wire net_sum46;
  wire net_sum47;
  wire net_sum48;
  wire net_sum49;
  wire net_sum5;
  wire net_sum50;
  wire net_sum51;
  wire net_sum52;
  wire net_sum53;
  wire net_sum54;
  wire net_sum55;
  wire net_sum56;
  wire net_sum57;
  wire net_sum58;
  wire net_sum59;
  wire net_sum6;
  wire net_sum60;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a60 = i0[60];
  assign net_a59 = i0[59];
  assign net_a58 = i0[58];
  assign net_a57 = i0[57];
  assign net_a56 = i0[56];
  assign net_a55 = i0[55];
  assign net_a54 = i0[54];
  assign net_a53 = i0[53];
  assign net_a52 = i0[52];
  assign net_a51 = i0[51];
  assign net_a50 = i0[50];
  assign net_a49 = i0[49];
  assign net_a48 = i0[48];
  assign net_a47 = i0[47];
  assign net_a46 = i0[46];
  assign net_a45 = i0[45];
  assign net_a44 = i0[44];
  assign net_a43 = i0[43];
  assign net_a42 = i0[42];
  assign net_a41 = i0[41];
  assign net_a40 = i0[40];
  assign net_a39 = i0[39];
  assign net_a38 = i0[38];
  assign net_a37 = i0[37];
  assign net_a36 = i0[36];
  assign net_a35 = i0[35];
  assign net_a34 = i0[34];
  assign net_a33 = i0[33];
  assign net_a32 = i0[32];
  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b60 = i1[60];
  assign net_b59 = i1[59];
  assign net_b58 = i1[58];
  assign net_b57 = i1[57];
  assign net_b56 = i1[56];
  assign net_b55 = i1[55];
  assign net_b54 = i1[54];
  assign net_b53 = i1[53];
  assign net_b52 = i1[52];
  assign net_b51 = i1[51];
  assign net_b50 = i1[50];
  assign net_b49 = i1[49];
  assign net_b48 = i1[48];
  assign net_b47 = i1[47];
  assign net_b46 = i1[46];
  assign net_b45 = i1[45];
  assign net_b44 = i1[44];
  assign net_b43 = i1[43];
  assign net_b42 = i1[42];
  assign net_b41 = i1[41];
  assign net_b40 = i1[40];
  assign net_b39 = i1[39];
  assign net_b38 = i1[38];
  assign net_b37 = i1[37];
  assign net_b36 = i1[36];
  assign net_b35 = i1[35];
  assign net_b34 = i1[34];
  assign net_b33 = i1[33];
  assign net_b32 = i1[32];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[60] = net_sum60;
  assign o[59] = net_sum59;
  assign o[58] = net_sum58;
  assign o[57] = net_sum57;
  assign o[56] = net_sum56;
  assign o[55] = net_sum55;
  assign o[54] = net_sum54;
  assign o[53] = net_sum53;
  assign o[52] = net_sum52;
  assign o[51] = net_sum51;
  assign o[50] = net_sum50;
  assign o[49] = net_sum49;
  assign o[48] = net_sum48;
  assign o[47] = net_sum47;
  assign o[46] = net_sum46;
  assign o[45] = net_sum45;
  assign o[44] = net_sum44;
  assign o[43] = net_sum43;
  assign o[42] = net_sum42;
  assign o[41] = net_sum41;
  assign o[40] = net_sum40;
  assign o[39] = net_sum39;
  assign o[38] = net_sum38;
  assign o[37] = net_sum37;
  assign o[36] = net_sum36;
  assign o[35] = net_sum35;
  assign o[34] = net_sum34;
  assign o[33] = net_sum33;
  assign o[32] = net_sum32;
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_32 (
    .a(net_a32),
    .b(net_b32),
    .c(net_cout31),
    .cout(net_cout32),
    .sum(net_sum32));
  AL_FADD comp_33 (
    .a(net_a33),
    .b(net_b33),
    .c(net_cout32),
    .cout(net_cout33),
    .sum(net_sum33));
  AL_FADD comp_34 (
    .a(net_a34),
    .b(net_b34),
    .c(net_cout33),
    .cout(net_cout34),
    .sum(net_sum34));
  AL_FADD comp_35 (
    .a(net_a35),
    .b(net_b35),
    .c(net_cout34),
    .cout(net_cout35),
    .sum(net_sum35));
  AL_FADD comp_36 (
    .a(net_a36),
    .b(net_b36),
    .c(net_cout35),
    .cout(net_cout36),
    .sum(net_sum36));
  AL_FADD comp_37 (
    .a(net_a37),
    .b(net_b37),
    .c(net_cout36),
    .cout(net_cout37),
    .sum(net_sum37));
  AL_FADD comp_38 (
    .a(net_a38),
    .b(net_b38),
    .c(net_cout37),
    .cout(net_cout38),
    .sum(net_sum38));
  AL_FADD comp_39 (
    .a(net_a39),
    .b(net_b39),
    .c(net_cout38),
    .cout(net_cout39),
    .sum(net_sum39));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_40 (
    .a(net_a40),
    .b(net_b40),
    .c(net_cout39),
    .cout(net_cout40),
    .sum(net_sum40));
  AL_FADD comp_41 (
    .a(net_a41),
    .b(net_b41),
    .c(net_cout40),
    .cout(net_cout41),
    .sum(net_sum41));
  AL_FADD comp_42 (
    .a(net_a42),
    .b(net_b42),
    .c(net_cout41),
    .cout(net_cout42),
    .sum(net_sum42));
  AL_FADD comp_43 (
    .a(net_a43),
    .b(net_b43),
    .c(net_cout42),
    .cout(net_cout43),
    .sum(net_sum43));
  AL_FADD comp_44 (
    .a(net_a44),
    .b(net_b44),
    .c(net_cout43),
    .cout(net_cout44),
    .sum(net_sum44));
  AL_FADD comp_45 (
    .a(net_a45),
    .b(net_b45),
    .c(net_cout44),
    .cout(net_cout45),
    .sum(net_sum45));
  AL_FADD comp_46 (
    .a(net_a46),
    .b(net_b46),
    .c(net_cout45),
    .cout(net_cout46),
    .sum(net_sum46));
  AL_FADD comp_47 (
    .a(net_a47),
    .b(net_b47),
    .c(net_cout46),
    .cout(net_cout47),
    .sum(net_sum47));
  AL_FADD comp_48 (
    .a(net_a48),
    .b(net_b48),
    .c(net_cout47),
    .cout(net_cout48),
    .sum(net_sum48));
  AL_FADD comp_49 (
    .a(net_a49),
    .b(net_b49),
    .c(net_cout48),
    .cout(net_cout49),
    .sum(net_sum49));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_50 (
    .a(net_a50),
    .b(net_b50),
    .c(net_cout49),
    .cout(net_cout50),
    .sum(net_sum50));
  AL_FADD comp_51 (
    .a(net_a51),
    .b(net_b51),
    .c(net_cout50),
    .cout(net_cout51),
    .sum(net_sum51));
  AL_FADD comp_52 (
    .a(net_a52),
    .b(net_b52),
    .c(net_cout51),
    .cout(net_cout52),
    .sum(net_sum52));
  AL_FADD comp_53 (
    .a(net_a53),
    .b(net_b53),
    .c(net_cout52),
    .cout(net_cout53),
    .sum(net_sum53));
  AL_FADD comp_54 (
    .a(net_a54),
    .b(net_b54),
    .c(net_cout53),
    .cout(net_cout54),
    .sum(net_sum54));
  AL_FADD comp_55 (
    .a(net_a55),
    .b(net_b55),
    .c(net_cout54),
    .cout(net_cout55),
    .sum(net_sum55));
  AL_FADD comp_56 (
    .a(net_a56),
    .b(net_b56),
    .c(net_cout55),
    .cout(net_cout56),
    .sum(net_sum56));
  AL_FADD comp_57 (
    .a(net_a57),
    .b(net_b57),
    .c(net_cout56),
    .cout(net_cout57),
    .sum(net_sum57));
  AL_FADD comp_58 (
    .a(net_a58),
    .b(net_b58),
    .c(net_cout57),
    .cout(net_cout58),
    .sum(net_sum58));
  AL_FADD comp_59 (
    .a(net_a59),
    .b(net_b59),
    .c(net_cout58),
    .cout(net_cout59),
    .sum(net_sum59));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_60 (
    .a(net_a60),
    .b(net_b60),
    .c(net_cout59),
    .cout(net_cout60),
    .sum(net_sum60));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output o;

  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;

  not none_diff (o, \or_or_xor_i0[0]_i1[0_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \xor_i0[4]_i1[4]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);

endmodule 

module eq_w9
  (
  i0,
  i1,
  o
  );

  input [8:0] i0;
  input [8:0] i1;
  output o;

  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[4]_i1[4_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;

  not none_diff (o, \or_or_or_xor_i0[0]_i_o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[4]_i1[4_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_or_xor_i0[4]_i1[4  (\or_or_xor_i0[4]_i1[4_o , \or_xor_i0[4]_i1[4]_o_o , \or_xor_i0[6]_i1[6]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \xor_i0[3]_i1[3]_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \or_xor_i0[7]_i1[7]_o_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);

endmodule 

module eq_w2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output o;

  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;

  not none_diff (o, \or_xor_i0[0]_i1[0]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);

endmodule 

module eq_w3
  (
  i0,
  i1,
  o
  );

  input [2:0] i0;
  input [2:0] i1;
  output o;

  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;

  not none_diff (o, \or_xor_i0[0]_i1[0]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);

endmodule 

module eq_w4
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output o;

  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;

  not none_diff (o, \or_or_xor_i0[0]_i1[0_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \xor_i0[3]_i1[3]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);

endmodule 

module eq_w32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire or_or_or_or_or_xor_i_o;
  wire \or_or_or_or_xor_i0[0_o ;
  wire \or_or_or_or_xor_i0[1_o ;
  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_or_xor_i0[16]__o ;
  wire \or_or_or_xor_i0[24]__o ;
  wire \or_or_or_xor_i0[8]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[12]_i1[_o ;
  wire \or_or_xor_i0[16]_i1[_o ;
  wire \or_or_xor_i0[20]_i1[_o ;
  wire \or_or_xor_i0[24]_i1[_o ;
  wire \or_or_xor_i0[28]_i1[_o ;
  wire \or_or_xor_i0[4]_i1[4_o ;
  wire \or_or_xor_i0[8]_i1[8_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[12]_i1[12]_o ;
  wire \or_xor_i0[14]_i1[14]_o ;
  wire \or_xor_i0[16]_i1[16]_o ;
  wire \or_xor_i0[18]_i1[18]_o ;
  wire \or_xor_i0[20]_i1[20]_o ;
  wire \or_xor_i0[22]_i1[22]_o ;
  wire \or_xor_i0[24]_i1[24]_o ;
  wire \or_xor_i0[26]_i1[26]_o ;
  wire \or_xor_i0[28]_i1[28]_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[30]_i1[30]_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[8]_i1[8]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[12]_i1[12]_o ;
  wire \xor_i0[13]_i1[13]_o ;
  wire \xor_i0[14]_i1[14]_o ;
  wire \xor_i0[15]_i1[15]_o ;
  wire \xor_i0[16]_i1[16]_o ;
  wire \xor_i0[17]_i1[17]_o ;
  wire \xor_i0[18]_i1[18]_o ;
  wire \xor_i0[19]_i1[19]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[20]_i1[20]_o ;
  wire \xor_i0[21]_i1[21]_o ;
  wire \xor_i0[22]_i1[22]_o ;
  wire \xor_i0[23]_i1[23]_o ;
  wire \xor_i0[24]_i1[24]_o ;
  wire \xor_i0[25]_i1[25]_o ;
  wire \xor_i0[26]_i1[26]_o ;
  wire \xor_i0[27]_i1[27]_o ;
  wire \xor_i0[28]_i1[28]_o ;
  wire \xor_i0[29]_i1[29]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[30]_i1[30]_o ;
  wire \xor_i0[31]_i1[31]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, or_or_or_or_or_xor_i_o);
  or or_or_or_or_or_xor_i (or_or_or_or_or_xor_i_o, \or_or_or_or_xor_i0[0_o , \or_or_or_or_xor_i0[1_o );
  or \or_or_or_or_xor_i0[0  (\or_or_or_or_xor_i0[0_o , \or_or_or_xor_i0[0]_i_o , \or_or_or_xor_i0[8]_i_o );
  or \or_or_or_or_xor_i0[1  (\or_or_or_or_xor_i0[1_o , \or_or_or_xor_i0[16]__o , \or_or_or_xor_i0[24]__o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[4]_i1[4_o );
  or \or_or_or_xor_i0[16]_  (\or_or_or_xor_i0[16]__o , \or_or_xor_i0[16]_i1[_o , \or_or_xor_i0[20]_i1[_o );
  or \or_or_or_xor_i0[24]_  (\or_or_or_xor_i0[24]__o , \or_or_xor_i0[24]_i1[_o , \or_or_xor_i0[28]_i1[_o );
  or \or_or_or_xor_i0[8]_i  (\or_or_or_xor_i0[8]_i_o , \or_or_xor_i0[8]_i1[8_o , \or_or_xor_i0[12]_i1[_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_or_xor_i0[12]_i1[  (\or_or_xor_i0[12]_i1[_o , \or_xor_i0[12]_i1[12]_o , \or_xor_i0[14]_i1[14]_o );
  or \or_or_xor_i0[16]_i1[  (\or_or_xor_i0[16]_i1[_o , \or_xor_i0[16]_i1[16]_o , \or_xor_i0[18]_i1[18]_o );
  or \or_or_xor_i0[20]_i1[  (\or_or_xor_i0[20]_i1[_o , \or_xor_i0[20]_i1[20]_o , \or_xor_i0[22]_i1[22]_o );
  or \or_or_xor_i0[24]_i1[  (\or_or_xor_i0[24]_i1[_o , \or_xor_i0[24]_i1[24]_o , \or_xor_i0[26]_i1[26]_o );
  or \or_or_xor_i0[28]_i1[  (\or_or_xor_i0[28]_i1[_o , \or_xor_i0[28]_i1[28]_o , \or_xor_i0[30]_i1[30]_o );
  or \or_or_xor_i0[4]_i1[4  (\or_or_xor_i0[4]_i1[4_o , \or_xor_i0[4]_i1[4]_o_o , \or_xor_i0[6]_i1[6]_o_o );
  or \or_or_xor_i0[8]_i1[8  (\or_or_xor_i0[8]_i1[8_o , \or_xor_i0[8]_i1[8]_o_o , \or_xor_i0[10]_i1[10]_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[12]_i1[12]  (\or_xor_i0[12]_i1[12]_o , \xor_i0[12]_i1[12]_o , \xor_i0[13]_i1[13]_o );
  or \or_xor_i0[14]_i1[14]  (\or_xor_i0[14]_i1[14]_o , \xor_i0[14]_i1[14]_o , \xor_i0[15]_i1[15]_o );
  or \or_xor_i0[16]_i1[16]  (\or_xor_i0[16]_i1[16]_o , \xor_i0[16]_i1[16]_o , \xor_i0[17]_i1[17]_o );
  or \or_xor_i0[18]_i1[18]  (\or_xor_i0[18]_i1[18]_o , \xor_i0[18]_i1[18]_o , \xor_i0[19]_i1[19]_o );
  or \or_xor_i0[20]_i1[20]  (\or_xor_i0[20]_i1[20]_o , \xor_i0[20]_i1[20]_o , \xor_i0[21]_i1[21]_o );
  or \or_xor_i0[22]_i1[22]  (\or_xor_i0[22]_i1[22]_o , \xor_i0[22]_i1[22]_o , \xor_i0[23]_i1[23]_o );
  or \or_xor_i0[24]_i1[24]  (\or_xor_i0[24]_i1[24]_o , \xor_i0[24]_i1[24]_o , \xor_i0[25]_i1[25]_o );
  or \or_xor_i0[26]_i1[26]  (\or_xor_i0[26]_i1[26]_o , \xor_i0[26]_i1[26]_o , \xor_i0[27]_i1[27]_o );
  or \or_xor_i0[28]_i1[28]  (\or_xor_i0[28]_i1[28]_o , \xor_i0[28]_i1[28]_o , \xor_i0[29]_i1[29]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \xor_i0[3]_i1[3]_o );
  or \or_xor_i0[30]_i1[30]  (\or_xor_i0[30]_i1[30]_o , \xor_i0[30]_i1[30]_o , \xor_i0[31]_i1[31]_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \xor_i0[7]_i1[7]_o );
  or \or_xor_i0[8]_i1[8]_o  (\or_xor_i0[8]_i1[8]_o_o , \xor_i0[8]_i1[8]_o , \xor_i0[9]_i1[9]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (\xor_i0[12]_i1[12]_o , i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (\xor_i0[13]_i1[13]_o , i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (\xor_i0[14]_i1[14]_o , i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (\xor_i0[15]_i1[15]_o , i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (\xor_i0[16]_i1[16]_o , i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (\xor_i0[17]_i1[17]_o , i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (\xor_i0[18]_i1[18]_o , i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (\xor_i0[19]_i1[19]_o , i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (\xor_i0[20]_i1[20]_o , i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (\xor_i0[21]_i1[21]_o , i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (\xor_i0[22]_i1[22]_o , i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (\xor_i0[23]_i1[23]_o , i0[23], i1[23]);
  xor \xor_i0[24]_i1[24]  (\xor_i0[24]_i1[24]_o , i0[24], i1[24]);
  xor \xor_i0[25]_i1[25]  (\xor_i0[25]_i1[25]_o , i0[25], i1[25]);
  xor \xor_i0[26]_i1[26]  (\xor_i0[26]_i1[26]_o , i0[26], i1[26]);
  xor \xor_i0[27]_i1[27]  (\xor_i0[27]_i1[27]_o , i0[27], i1[27]);
  xor \xor_i0[28]_i1[28]  (\xor_i0[28]_i1[28]_o , i0[28], i1[28]);
  xor \xor_i0[29]_i1[29]  (\xor_i0[29]_i1[29]_o , i0[29], i1[29]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[30]_i1[30]  (\xor_i0[30]_i1[30]_o , i0[30], i1[30]);
  xor \xor_i0[31]_i1[31]  (\xor_i0[31]_i1[31]_o , i0[31], i1[31]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module binary_mux_s1_w1
  (
  i0,
  i1,
  sel,
  o
  );

  input i0;
  input i1;
  input sel;
  output o;


  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel),
    .o(o));

endmodule 

module binary_mux_s2_w1
  (
  i0,
  i1,
  i2,
  i3,
  sel,
  o
  );

  input i0;
  input i1;
  input i2;
  input i3;
  input [1:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(o));

endmodule 

module ne_w4
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output o;

  wire [3:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module reg_ar_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(setout),
    .reset(reset),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module add_pu2_mu2_o2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output [1:0] o;

  wire net_a0;
  wire net_a1;
  wire net_b0;
  wire net_b1;
  wire net_cout0;
  wire net_cout1;
  wire net_nb0;
  wire net_nb1;
  wire net_sum0;
  wire net_sum1;

  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);

endmodule 

module reg_sr_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(setout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module add_pu9_mu9_o9
  (
  i0,
  i1,
  o
  );

  input [8:0] i0;
  input [8:0] i1;
  output [8:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_nb0;
  wire net_nb1;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;

  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);

endmodule 

module add_pu64_pu64_o64
  (
  i0,
  i1,
  o
  );

  input [63:0] i0;
  input [63:0] i1;
  output [63:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a32;
  wire net_a33;
  wire net_a34;
  wire net_a35;
  wire net_a36;
  wire net_a37;
  wire net_a38;
  wire net_a39;
  wire net_a4;
  wire net_a40;
  wire net_a41;
  wire net_a42;
  wire net_a43;
  wire net_a44;
  wire net_a45;
  wire net_a46;
  wire net_a47;
  wire net_a48;
  wire net_a49;
  wire net_a5;
  wire net_a50;
  wire net_a51;
  wire net_a52;
  wire net_a53;
  wire net_a54;
  wire net_a55;
  wire net_a56;
  wire net_a57;
  wire net_a58;
  wire net_a59;
  wire net_a6;
  wire net_a60;
  wire net_a61;
  wire net_a62;
  wire net_a63;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b32;
  wire net_b33;
  wire net_b34;
  wire net_b35;
  wire net_b36;
  wire net_b37;
  wire net_b38;
  wire net_b39;
  wire net_b4;
  wire net_b40;
  wire net_b41;
  wire net_b42;
  wire net_b43;
  wire net_b44;
  wire net_b45;
  wire net_b46;
  wire net_b47;
  wire net_b48;
  wire net_b49;
  wire net_b5;
  wire net_b50;
  wire net_b51;
  wire net_b52;
  wire net_b53;
  wire net_b54;
  wire net_b55;
  wire net_b56;
  wire net_b57;
  wire net_b58;
  wire net_b59;
  wire net_b6;
  wire net_b60;
  wire net_b61;
  wire net_b62;
  wire net_b63;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout32;
  wire net_cout33;
  wire net_cout34;
  wire net_cout35;
  wire net_cout36;
  wire net_cout37;
  wire net_cout38;
  wire net_cout39;
  wire net_cout4;
  wire net_cout40;
  wire net_cout41;
  wire net_cout42;
  wire net_cout43;
  wire net_cout44;
  wire net_cout45;
  wire net_cout46;
  wire net_cout47;
  wire net_cout48;
  wire net_cout49;
  wire net_cout5;
  wire net_cout50;
  wire net_cout51;
  wire net_cout52;
  wire net_cout53;
  wire net_cout54;
  wire net_cout55;
  wire net_cout56;
  wire net_cout57;
  wire net_cout58;
  wire net_cout59;
  wire net_cout6;
  wire net_cout60;
  wire net_cout61;
  wire net_cout62;
  wire net_cout63;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum32;
  wire net_sum33;
  wire net_sum34;
  wire net_sum35;
  wire net_sum36;
  wire net_sum37;
  wire net_sum38;
  wire net_sum39;
  wire net_sum4;
  wire net_sum40;
  wire net_sum41;
  wire net_sum42;
  wire net_sum43;
  wire net_sum44;
  wire net_sum45;
  wire net_sum46;
  wire net_sum47;
  wire net_sum48;
  wire net_sum49;
  wire net_sum5;
  wire net_sum50;
  wire net_sum51;
  wire net_sum52;
  wire net_sum53;
  wire net_sum54;
  wire net_sum55;
  wire net_sum56;
  wire net_sum57;
  wire net_sum58;
  wire net_sum59;
  wire net_sum6;
  wire net_sum60;
  wire net_sum61;
  wire net_sum62;
  wire net_sum63;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a63 = i0[63];
  assign net_a62 = i0[62];
  assign net_a61 = i0[61];
  assign net_a60 = i0[60];
  assign net_a59 = i0[59];
  assign net_a58 = i0[58];
  assign net_a57 = i0[57];
  assign net_a56 = i0[56];
  assign net_a55 = i0[55];
  assign net_a54 = i0[54];
  assign net_a53 = i0[53];
  assign net_a52 = i0[52];
  assign net_a51 = i0[51];
  assign net_a50 = i0[50];
  assign net_a49 = i0[49];
  assign net_a48 = i0[48];
  assign net_a47 = i0[47];
  assign net_a46 = i0[46];
  assign net_a45 = i0[45];
  assign net_a44 = i0[44];
  assign net_a43 = i0[43];
  assign net_a42 = i0[42];
  assign net_a41 = i0[41];
  assign net_a40 = i0[40];
  assign net_a39 = i0[39];
  assign net_a38 = i0[38];
  assign net_a37 = i0[37];
  assign net_a36 = i0[36];
  assign net_a35 = i0[35];
  assign net_a34 = i0[34];
  assign net_a33 = i0[33];
  assign net_a32 = i0[32];
  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b63 = i1[63];
  assign net_b62 = i1[62];
  assign net_b61 = i1[61];
  assign net_b60 = i1[60];
  assign net_b59 = i1[59];
  assign net_b58 = i1[58];
  assign net_b57 = i1[57];
  assign net_b56 = i1[56];
  assign net_b55 = i1[55];
  assign net_b54 = i1[54];
  assign net_b53 = i1[53];
  assign net_b52 = i1[52];
  assign net_b51 = i1[51];
  assign net_b50 = i1[50];
  assign net_b49 = i1[49];
  assign net_b48 = i1[48];
  assign net_b47 = i1[47];
  assign net_b46 = i1[46];
  assign net_b45 = i1[45];
  assign net_b44 = i1[44];
  assign net_b43 = i1[43];
  assign net_b42 = i1[42];
  assign net_b41 = i1[41];
  assign net_b40 = i1[40];
  assign net_b39 = i1[39];
  assign net_b38 = i1[38];
  assign net_b37 = i1[37];
  assign net_b36 = i1[36];
  assign net_b35 = i1[35];
  assign net_b34 = i1[34];
  assign net_b33 = i1[33];
  assign net_b32 = i1[32];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[63] = net_sum63;
  assign o[62] = net_sum62;
  assign o[61] = net_sum61;
  assign o[60] = net_sum60;
  assign o[59] = net_sum59;
  assign o[58] = net_sum58;
  assign o[57] = net_sum57;
  assign o[56] = net_sum56;
  assign o[55] = net_sum55;
  assign o[54] = net_sum54;
  assign o[53] = net_sum53;
  assign o[52] = net_sum52;
  assign o[51] = net_sum51;
  assign o[50] = net_sum50;
  assign o[49] = net_sum49;
  assign o[48] = net_sum48;
  assign o[47] = net_sum47;
  assign o[46] = net_sum46;
  assign o[45] = net_sum45;
  assign o[44] = net_sum44;
  assign o[43] = net_sum43;
  assign o[42] = net_sum42;
  assign o[41] = net_sum41;
  assign o[40] = net_sum40;
  assign o[39] = net_sum39;
  assign o[38] = net_sum38;
  assign o[37] = net_sum37;
  assign o[36] = net_sum36;
  assign o[35] = net_sum35;
  assign o[34] = net_sum34;
  assign o[33] = net_sum33;
  assign o[32] = net_sum32;
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_32 (
    .a(net_a32),
    .b(net_b32),
    .c(net_cout31),
    .cout(net_cout32),
    .sum(net_sum32));
  AL_FADD comp_33 (
    .a(net_a33),
    .b(net_b33),
    .c(net_cout32),
    .cout(net_cout33),
    .sum(net_sum33));
  AL_FADD comp_34 (
    .a(net_a34),
    .b(net_b34),
    .c(net_cout33),
    .cout(net_cout34),
    .sum(net_sum34));
  AL_FADD comp_35 (
    .a(net_a35),
    .b(net_b35),
    .c(net_cout34),
    .cout(net_cout35),
    .sum(net_sum35));
  AL_FADD comp_36 (
    .a(net_a36),
    .b(net_b36),
    .c(net_cout35),
    .cout(net_cout36),
    .sum(net_sum36));
  AL_FADD comp_37 (
    .a(net_a37),
    .b(net_b37),
    .c(net_cout36),
    .cout(net_cout37),
    .sum(net_sum37));
  AL_FADD comp_38 (
    .a(net_a38),
    .b(net_b38),
    .c(net_cout37),
    .cout(net_cout38),
    .sum(net_sum38));
  AL_FADD comp_39 (
    .a(net_a39),
    .b(net_b39),
    .c(net_cout38),
    .cout(net_cout39),
    .sum(net_sum39));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_40 (
    .a(net_a40),
    .b(net_b40),
    .c(net_cout39),
    .cout(net_cout40),
    .sum(net_sum40));
  AL_FADD comp_41 (
    .a(net_a41),
    .b(net_b41),
    .c(net_cout40),
    .cout(net_cout41),
    .sum(net_sum41));
  AL_FADD comp_42 (
    .a(net_a42),
    .b(net_b42),
    .c(net_cout41),
    .cout(net_cout42),
    .sum(net_sum42));
  AL_FADD comp_43 (
    .a(net_a43),
    .b(net_b43),
    .c(net_cout42),
    .cout(net_cout43),
    .sum(net_sum43));
  AL_FADD comp_44 (
    .a(net_a44),
    .b(net_b44),
    .c(net_cout43),
    .cout(net_cout44),
    .sum(net_sum44));
  AL_FADD comp_45 (
    .a(net_a45),
    .b(net_b45),
    .c(net_cout44),
    .cout(net_cout45),
    .sum(net_sum45));
  AL_FADD comp_46 (
    .a(net_a46),
    .b(net_b46),
    .c(net_cout45),
    .cout(net_cout46),
    .sum(net_sum46));
  AL_FADD comp_47 (
    .a(net_a47),
    .b(net_b47),
    .c(net_cout46),
    .cout(net_cout47),
    .sum(net_sum47));
  AL_FADD comp_48 (
    .a(net_a48),
    .b(net_b48),
    .c(net_cout47),
    .cout(net_cout48),
    .sum(net_sum48));
  AL_FADD comp_49 (
    .a(net_a49),
    .b(net_b49),
    .c(net_cout48),
    .cout(net_cout49),
    .sum(net_sum49));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_50 (
    .a(net_a50),
    .b(net_b50),
    .c(net_cout49),
    .cout(net_cout50),
    .sum(net_sum50));
  AL_FADD comp_51 (
    .a(net_a51),
    .b(net_b51),
    .c(net_cout50),
    .cout(net_cout51),
    .sum(net_sum51));
  AL_FADD comp_52 (
    .a(net_a52),
    .b(net_b52),
    .c(net_cout51),
    .cout(net_cout52),
    .sum(net_sum52));
  AL_FADD comp_53 (
    .a(net_a53),
    .b(net_b53),
    .c(net_cout52),
    .cout(net_cout53),
    .sum(net_sum53));
  AL_FADD comp_54 (
    .a(net_a54),
    .b(net_b54),
    .c(net_cout53),
    .cout(net_cout54),
    .sum(net_sum54));
  AL_FADD comp_55 (
    .a(net_a55),
    .b(net_b55),
    .c(net_cout54),
    .cout(net_cout55),
    .sum(net_sum55));
  AL_FADD comp_56 (
    .a(net_a56),
    .b(net_b56),
    .c(net_cout55),
    .cout(net_cout56),
    .sum(net_sum56));
  AL_FADD comp_57 (
    .a(net_a57),
    .b(net_b57),
    .c(net_cout56),
    .cout(net_cout57),
    .sum(net_sum57));
  AL_FADD comp_58 (
    .a(net_a58),
    .b(net_b58),
    .c(net_cout57),
    .cout(net_cout58),
    .sum(net_sum58));
  AL_FADD comp_59 (
    .a(net_a59),
    .b(net_b59),
    .c(net_cout58),
    .cout(net_cout59),
    .sum(net_sum59));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_60 (
    .a(net_a60),
    .b(net_b60),
    .c(net_cout59),
    .cout(net_cout60),
    .sum(net_sum60));
  AL_FADD comp_61 (
    .a(net_a61),
    .b(net_b61),
    .c(net_cout60),
    .cout(net_cout61),
    .sum(net_sum61));
  AL_FADD comp_62 (
    .a(net_a62),
    .b(net_b62),
    .c(net_cout61),
    .cout(net_cout62),
    .sum(net_sum62));
  AL_FADD comp_63 (
    .a(net_a63),
    .b(net_b63),
    .c(net_cout62),
    .cout(net_cout63),
    .sum(net_sum63));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w52
  (
  i0,
  i1,
  o
  );

  input [51:0] i0;
  input [51:0] i1;
  output o;

  wire or_or_or_or_or_xor_i_o;
  wire \or_or_or_or_xor_i0[0_o ;
  wire \or_or_or_or_xor_i0[2_o ;
  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_or_xor_i0[13]__o ;
  wire \or_or_or_xor_i0[26]__o ;
  wire \or_or_or_xor_i0[39]__o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[13]_i1[_o ;
  wire \or_or_xor_i0[19]_i1[_o ;
  wire \or_or_xor_i0[22]_i1[_o ;
  wire \or_or_xor_i0[26]_i1[_o ;
  wire \or_or_xor_i0[32]_i1[_o ;
  wire \or_or_xor_i0[35]_i1[_o ;
  wire \or_or_xor_i0[39]_i1[_o ;
  wire \or_or_xor_i0[45]_i1[_o ;
  wire \or_or_xor_i0[48]_i1[_o ;
  wire \or_or_xor_i0[6]_i1[6_o ;
  wire \or_or_xor_i0[9]_i1[9_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[11]_i1[11]_o ;
  wire \or_xor_i0[13]_i1[13]_o ;
  wire \or_xor_i0[14]_i1[14]_o ;
  wire \or_xor_i0[16]_i1[16]_o ;
  wire \or_xor_i0[17]_i1[17]_o ;
  wire \or_xor_i0[19]_i1[19]_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[20]_i1[20]_o ;
  wire \or_xor_i0[22]_i1[22]_o ;
  wire \or_xor_i0[24]_i1[24]_o ;
  wire \or_xor_i0[26]_i1[26]_o ;
  wire \or_xor_i0[27]_i1[27]_o ;
  wire \or_xor_i0[29]_i1[29]_o ;
  wire \or_xor_i0[30]_i1[30]_o ;
  wire \or_xor_i0[32]_i1[32]_o ;
  wire \or_xor_i0[33]_i1[33]_o ;
  wire \or_xor_i0[35]_i1[35]_o ;
  wire \or_xor_i0[37]_i1[37]_o ;
  wire \or_xor_i0[39]_i1[39]_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[40]_i1[40]_o ;
  wire \or_xor_i0[42]_i1[42]_o ;
  wire \or_xor_i0[43]_i1[43]_o ;
  wire \or_xor_i0[45]_i1[45]_o ;
  wire \or_xor_i0[46]_i1[46]_o ;
  wire \or_xor_i0[48]_i1[48]_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[50]_i1[50]_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[12]_i1[12]_o ;
  wire \xor_i0[13]_i1[13]_o ;
  wire \xor_i0[14]_i1[14]_o ;
  wire \xor_i0[15]_i1[15]_o ;
  wire \xor_i0[16]_i1[16]_o ;
  wire \xor_i0[17]_i1[17]_o ;
  wire \xor_i0[18]_i1[18]_o ;
  wire \xor_i0[19]_i1[19]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[20]_i1[20]_o ;
  wire \xor_i0[21]_i1[21]_o ;
  wire \xor_i0[22]_i1[22]_o ;
  wire \xor_i0[23]_i1[23]_o ;
  wire \xor_i0[24]_i1[24]_o ;
  wire \xor_i0[25]_i1[25]_o ;
  wire \xor_i0[26]_i1[26]_o ;
  wire \xor_i0[27]_i1[27]_o ;
  wire \xor_i0[28]_i1[28]_o ;
  wire \xor_i0[29]_i1[29]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[30]_i1[30]_o ;
  wire \xor_i0[31]_i1[31]_o ;
  wire \xor_i0[32]_i1[32]_o ;
  wire \xor_i0[33]_i1[33]_o ;
  wire \xor_i0[34]_i1[34]_o ;
  wire \xor_i0[35]_i1[35]_o ;
  wire \xor_i0[36]_i1[36]_o ;
  wire \xor_i0[37]_i1[37]_o ;
  wire \xor_i0[38]_i1[38]_o ;
  wire \xor_i0[39]_i1[39]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[40]_i1[40]_o ;
  wire \xor_i0[41]_i1[41]_o ;
  wire \xor_i0[42]_i1[42]_o ;
  wire \xor_i0[43]_i1[43]_o ;
  wire \xor_i0[44]_i1[44]_o ;
  wire \xor_i0[45]_i1[45]_o ;
  wire \xor_i0[46]_i1[46]_o ;
  wire \xor_i0[47]_i1[47]_o ;
  wire \xor_i0[48]_i1[48]_o ;
  wire \xor_i0[49]_i1[49]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[50]_i1[50]_o ;
  wire \xor_i0[51]_i1[51]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, or_or_or_or_or_xor_i_o);
  or or_or_or_or_or_xor_i (or_or_or_or_or_xor_i_o, \or_or_or_or_xor_i0[0_o , \or_or_or_or_xor_i0[2_o );
  or \or_or_or_or_xor_i0[0  (\or_or_or_or_xor_i0[0_o , \or_or_or_xor_i0[0]_i_o , \or_or_or_xor_i0[13]__o );
  or \or_or_or_or_xor_i0[2  (\or_or_or_or_xor_i0[2_o , \or_or_or_xor_i0[26]__o , \or_or_or_xor_i0[39]__o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[6]_i1[6_o );
  or \or_or_or_xor_i0[13]_  (\or_or_or_xor_i0[13]__o , \or_or_xor_i0[13]_i1[_o , \or_or_xor_i0[19]_i1[_o );
  or \or_or_or_xor_i0[26]_  (\or_or_or_xor_i0[26]__o , \or_or_xor_i0[26]_i1[_o , \or_or_xor_i0[32]_i1[_o );
  or \or_or_or_xor_i0[39]_  (\or_or_or_xor_i0[39]__o , \or_or_xor_i0[39]_i1[_o , \or_or_xor_i0[45]_i1[_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_or_xor_i0[13]_i1[  (\or_or_xor_i0[13]_i1[_o , \or_xor_i0[13]_i1[13]_o , \or_xor_i0[16]_i1[16]_o );
  or \or_or_xor_i0[19]_i1[  (\or_or_xor_i0[19]_i1[_o , \or_xor_i0[19]_i1[19]_o , \or_or_xor_i0[22]_i1[_o );
  or \or_or_xor_i0[22]_i1[  (\or_or_xor_i0[22]_i1[_o , \or_xor_i0[22]_i1[22]_o , \or_xor_i0[24]_i1[24]_o );
  or \or_or_xor_i0[26]_i1[  (\or_or_xor_i0[26]_i1[_o , \or_xor_i0[26]_i1[26]_o , \or_xor_i0[29]_i1[29]_o );
  or \or_or_xor_i0[32]_i1[  (\or_or_xor_i0[32]_i1[_o , \or_xor_i0[32]_i1[32]_o , \or_or_xor_i0[35]_i1[_o );
  or \or_or_xor_i0[35]_i1[  (\or_or_xor_i0[35]_i1[_o , \or_xor_i0[35]_i1[35]_o , \or_xor_i0[37]_i1[37]_o );
  or \or_or_xor_i0[39]_i1[  (\or_or_xor_i0[39]_i1[_o , \or_xor_i0[39]_i1[39]_o , \or_xor_i0[42]_i1[42]_o );
  or \or_or_xor_i0[45]_i1[  (\or_or_xor_i0[45]_i1[_o , \or_xor_i0[45]_i1[45]_o , \or_or_xor_i0[48]_i1[_o );
  or \or_or_xor_i0[48]_i1[  (\or_or_xor_i0[48]_i1[_o , \or_xor_i0[48]_i1[48]_o , \or_xor_i0[50]_i1[50]_o );
  or \or_or_xor_i0[6]_i1[6  (\or_or_xor_i0[6]_i1[6_o , \or_xor_i0[6]_i1[6]_o_o , \or_or_xor_i0[9]_i1[9_o );
  or \or_or_xor_i0[9]_i1[9  (\or_or_xor_i0[9]_i1[9_o , \or_xor_i0[9]_i1[9]_o_o , \or_xor_i0[11]_i1[11]_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[11]_i1[11]  (\or_xor_i0[11]_i1[11]_o , \xor_i0[11]_i1[11]_o , \xor_i0[12]_i1[12]_o );
  or \or_xor_i0[13]_i1[13]  (\or_xor_i0[13]_i1[13]_o , \xor_i0[13]_i1[13]_o , \or_xor_i0[14]_i1[14]_o );
  or \or_xor_i0[14]_i1[14]  (\or_xor_i0[14]_i1[14]_o , \xor_i0[14]_i1[14]_o , \xor_i0[15]_i1[15]_o );
  or \or_xor_i0[16]_i1[16]  (\or_xor_i0[16]_i1[16]_o , \xor_i0[16]_i1[16]_o , \or_xor_i0[17]_i1[17]_o );
  or \or_xor_i0[17]_i1[17]  (\or_xor_i0[17]_i1[17]_o , \xor_i0[17]_i1[17]_o , \xor_i0[18]_i1[18]_o );
  or \or_xor_i0[19]_i1[19]  (\or_xor_i0[19]_i1[19]_o , \xor_i0[19]_i1[19]_o , \or_xor_i0[20]_i1[20]_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[20]_i1[20]  (\or_xor_i0[20]_i1[20]_o , \xor_i0[20]_i1[20]_o , \xor_i0[21]_i1[21]_o );
  or \or_xor_i0[22]_i1[22]  (\or_xor_i0[22]_i1[22]_o , \xor_i0[22]_i1[22]_o , \xor_i0[23]_i1[23]_o );
  or \or_xor_i0[24]_i1[24]  (\or_xor_i0[24]_i1[24]_o , \xor_i0[24]_i1[24]_o , \xor_i0[25]_i1[25]_o );
  or \or_xor_i0[26]_i1[26]  (\or_xor_i0[26]_i1[26]_o , \xor_i0[26]_i1[26]_o , \or_xor_i0[27]_i1[27]_o );
  or \or_xor_i0[27]_i1[27]  (\or_xor_i0[27]_i1[27]_o , \xor_i0[27]_i1[27]_o , \xor_i0[28]_i1[28]_o );
  or \or_xor_i0[29]_i1[29]  (\or_xor_i0[29]_i1[29]_o , \xor_i0[29]_i1[29]_o , \or_xor_i0[30]_i1[30]_o );
  or \or_xor_i0[30]_i1[30]  (\or_xor_i0[30]_i1[30]_o , \xor_i0[30]_i1[30]_o , \xor_i0[31]_i1[31]_o );
  or \or_xor_i0[32]_i1[32]  (\or_xor_i0[32]_i1[32]_o , \xor_i0[32]_i1[32]_o , \or_xor_i0[33]_i1[33]_o );
  or \or_xor_i0[33]_i1[33]  (\or_xor_i0[33]_i1[33]_o , \xor_i0[33]_i1[33]_o , \xor_i0[34]_i1[34]_o );
  or \or_xor_i0[35]_i1[35]  (\or_xor_i0[35]_i1[35]_o , \xor_i0[35]_i1[35]_o , \xor_i0[36]_i1[36]_o );
  or \or_xor_i0[37]_i1[37]  (\or_xor_i0[37]_i1[37]_o , \xor_i0[37]_i1[37]_o , \xor_i0[38]_i1[38]_o );
  or \or_xor_i0[39]_i1[39]  (\or_xor_i0[39]_i1[39]_o , \xor_i0[39]_i1[39]_o , \or_xor_i0[40]_i1[40]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \or_xor_i0[4]_i1[4]_o_o );
  or \or_xor_i0[40]_i1[40]  (\or_xor_i0[40]_i1[40]_o , \xor_i0[40]_i1[40]_o , \xor_i0[41]_i1[41]_o );
  or \or_xor_i0[42]_i1[42]  (\or_xor_i0[42]_i1[42]_o , \xor_i0[42]_i1[42]_o , \or_xor_i0[43]_i1[43]_o );
  or \or_xor_i0[43]_i1[43]  (\or_xor_i0[43]_i1[43]_o , \xor_i0[43]_i1[43]_o , \xor_i0[44]_i1[44]_o );
  or \or_xor_i0[45]_i1[45]  (\or_xor_i0[45]_i1[45]_o , \xor_i0[45]_i1[45]_o , \or_xor_i0[46]_i1[46]_o );
  or \or_xor_i0[46]_i1[46]  (\or_xor_i0[46]_i1[46]_o , \xor_i0[46]_i1[46]_o , \xor_i0[47]_i1[47]_o );
  or \or_xor_i0[48]_i1[48]  (\or_xor_i0[48]_i1[48]_o , \xor_i0[48]_i1[48]_o , \xor_i0[49]_i1[49]_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[50]_i1[50]  (\or_xor_i0[50]_i1[50]_o , \xor_i0[50]_i1[50]_o , \xor_i0[51]_i1[51]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \or_xor_i0[7]_i1[7]_o_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (\xor_i0[12]_i1[12]_o , i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (\xor_i0[13]_i1[13]_o , i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (\xor_i0[14]_i1[14]_o , i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (\xor_i0[15]_i1[15]_o , i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (\xor_i0[16]_i1[16]_o , i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (\xor_i0[17]_i1[17]_o , i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (\xor_i0[18]_i1[18]_o , i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (\xor_i0[19]_i1[19]_o , i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (\xor_i0[20]_i1[20]_o , i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (\xor_i0[21]_i1[21]_o , i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (\xor_i0[22]_i1[22]_o , i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (\xor_i0[23]_i1[23]_o , i0[23], i1[23]);
  xor \xor_i0[24]_i1[24]  (\xor_i0[24]_i1[24]_o , i0[24], i1[24]);
  xor \xor_i0[25]_i1[25]  (\xor_i0[25]_i1[25]_o , i0[25], i1[25]);
  xor \xor_i0[26]_i1[26]  (\xor_i0[26]_i1[26]_o , i0[26], i1[26]);
  xor \xor_i0[27]_i1[27]  (\xor_i0[27]_i1[27]_o , i0[27], i1[27]);
  xor \xor_i0[28]_i1[28]  (\xor_i0[28]_i1[28]_o , i0[28], i1[28]);
  xor \xor_i0[29]_i1[29]  (\xor_i0[29]_i1[29]_o , i0[29], i1[29]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[30]_i1[30]  (\xor_i0[30]_i1[30]_o , i0[30], i1[30]);
  xor \xor_i0[31]_i1[31]  (\xor_i0[31]_i1[31]_o , i0[31], i1[31]);
  xor \xor_i0[32]_i1[32]  (\xor_i0[32]_i1[32]_o , i0[32], i1[32]);
  xor \xor_i0[33]_i1[33]  (\xor_i0[33]_i1[33]_o , i0[33], i1[33]);
  xor \xor_i0[34]_i1[34]  (\xor_i0[34]_i1[34]_o , i0[34], i1[34]);
  xor \xor_i0[35]_i1[35]  (\xor_i0[35]_i1[35]_o , i0[35], i1[35]);
  xor \xor_i0[36]_i1[36]  (\xor_i0[36]_i1[36]_o , i0[36], i1[36]);
  xor \xor_i0[37]_i1[37]  (\xor_i0[37]_i1[37]_o , i0[37], i1[37]);
  xor \xor_i0[38]_i1[38]  (\xor_i0[38]_i1[38]_o , i0[38], i1[38]);
  xor \xor_i0[39]_i1[39]  (\xor_i0[39]_i1[39]_o , i0[39], i1[39]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[40]_i1[40]  (\xor_i0[40]_i1[40]_o , i0[40], i1[40]);
  xor \xor_i0[41]_i1[41]  (\xor_i0[41]_i1[41]_o , i0[41], i1[41]);
  xor \xor_i0[42]_i1[42]  (\xor_i0[42]_i1[42]_o , i0[42], i1[42]);
  xor \xor_i0[43]_i1[43]  (\xor_i0[43]_i1[43]_o , i0[43], i1[43]);
  xor \xor_i0[44]_i1[44]  (\xor_i0[44]_i1[44]_o , i0[44], i1[44]);
  xor \xor_i0[45]_i1[45]  (\xor_i0[45]_i1[45]_o , i0[45], i1[45]);
  xor \xor_i0[46]_i1[46]  (\xor_i0[46]_i1[46]_o , i0[46], i1[46]);
  xor \xor_i0[47]_i1[47]  (\xor_i0[47]_i1[47]_o , i0[47], i1[47]);
  xor \xor_i0[48]_i1[48]  (\xor_i0[48]_i1[48]_o , i0[48], i1[48]);
  xor \xor_i0[49]_i1[49]  (\xor_i0[49]_i1[49]_o , i0[49], i1[49]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[50]_i1[50]  (\xor_i0[50]_i1[50]_o , i0[50], i1[50]);
  xor \xor_i0[51]_i1[51]  (\xor_i0[51]_i1[51]_o , i0[51], i1[51]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module add_pu60_pu60_o61
  (
  i0,
  i1,
  o
  );

  input [59:0] i0;
  input [59:0] i1;
  output [60:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a32;
  wire net_a33;
  wire net_a34;
  wire net_a35;
  wire net_a36;
  wire net_a37;
  wire net_a38;
  wire net_a39;
  wire net_a4;
  wire net_a40;
  wire net_a41;
  wire net_a42;
  wire net_a43;
  wire net_a44;
  wire net_a45;
  wire net_a46;
  wire net_a47;
  wire net_a48;
  wire net_a49;
  wire net_a5;
  wire net_a50;
  wire net_a51;
  wire net_a52;
  wire net_a53;
  wire net_a54;
  wire net_a55;
  wire net_a56;
  wire net_a57;
  wire net_a58;
  wire net_a59;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b32;
  wire net_b33;
  wire net_b34;
  wire net_b35;
  wire net_b36;
  wire net_b37;
  wire net_b38;
  wire net_b39;
  wire net_b4;
  wire net_b40;
  wire net_b41;
  wire net_b42;
  wire net_b43;
  wire net_b44;
  wire net_b45;
  wire net_b46;
  wire net_b47;
  wire net_b48;
  wire net_b49;
  wire net_b5;
  wire net_b50;
  wire net_b51;
  wire net_b52;
  wire net_b53;
  wire net_b54;
  wire net_b55;
  wire net_b56;
  wire net_b57;
  wire net_b58;
  wire net_b59;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout32;
  wire net_cout33;
  wire net_cout34;
  wire net_cout35;
  wire net_cout36;
  wire net_cout37;
  wire net_cout38;
  wire net_cout39;
  wire net_cout4;
  wire net_cout40;
  wire net_cout41;
  wire net_cout42;
  wire net_cout43;
  wire net_cout44;
  wire net_cout45;
  wire net_cout46;
  wire net_cout47;
  wire net_cout48;
  wire net_cout49;
  wire net_cout5;
  wire net_cout50;
  wire net_cout51;
  wire net_cout52;
  wire net_cout53;
  wire net_cout54;
  wire net_cout55;
  wire net_cout56;
  wire net_cout57;
  wire net_cout58;
  wire net_cout59;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum32;
  wire net_sum33;
  wire net_sum34;
  wire net_sum35;
  wire net_sum36;
  wire net_sum37;
  wire net_sum38;
  wire net_sum39;
  wire net_sum4;
  wire net_sum40;
  wire net_sum41;
  wire net_sum42;
  wire net_sum43;
  wire net_sum44;
  wire net_sum45;
  wire net_sum46;
  wire net_sum47;
  wire net_sum48;
  wire net_sum49;
  wire net_sum5;
  wire net_sum50;
  wire net_sum51;
  wire net_sum52;
  wire net_sum53;
  wire net_sum54;
  wire net_sum55;
  wire net_sum56;
  wire net_sum57;
  wire net_sum58;
  wire net_sum59;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a59 = i0[59];
  assign net_a58 = i0[58];
  assign net_a57 = i0[57];
  assign net_a56 = i0[56];
  assign net_a55 = i0[55];
  assign net_a54 = i0[54];
  assign net_a53 = i0[53];
  assign net_a52 = i0[52];
  assign net_a51 = i0[51];
  assign net_a50 = i0[50];
  assign net_a49 = i0[49];
  assign net_a48 = i0[48];
  assign net_a47 = i0[47];
  assign net_a46 = i0[46];
  assign net_a45 = i0[45];
  assign net_a44 = i0[44];
  assign net_a43 = i0[43];
  assign net_a42 = i0[42];
  assign net_a41 = i0[41];
  assign net_a40 = i0[40];
  assign net_a39 = i0[39];
  assign net_a38 = i0[38];
  assign net_a37 = i0[37];
  assign net_a36 = i0[36];
  assign net_a35 = i0[35];
  assign net_a34 = i0[34];
  assign net_a33 = i0[33];
  assign net_a32 = i0[32];
  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b59 = i1[59];
  assign net_b58 = i1[58];
  assign net_b57 = i1[57];
  assign net_b56 = i1[56];
  assign net_b55 = i1[55];
  assign net_b54 = i1[54];
  assign net_b53 = i1[53];
  assign net_b52 = i1[52];
  assign net_b51 = i1[51];
  assign net_b50 = i1[50];
  assign net_b49 = i1[49];
  assign net_b48 = i1[48];
  assign net_b47 = i1[47];
  assign net_b46 = i1[46];
  assign net_b45 = i1[45];
  assign net_b44 = i1[44];
  assign net_b43 = i1[43];
  assign net_b42 = i1[42];
  assign net_b41 = i1[41];
  assign net_b40 = i1[40];
  assign net_b39 = i1[39];
  assign net_b38 = i1[38];
  assign net_b37 = i1[37];
  assign net_b36 = i1[36];
  assign net_b35 = i1[35];
  assign net_b34 = i1[34];
  assign net_b33 = i1[33];
  assign net_b32 = i1[32];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[60] = net_cout59;
  assign o[59] = net_sum59;
  assign o[58] = net_sum58;
  assign o[57] = net_sum57;
  assign o[56] = net_sum56;
  assign o[55] = net_sum55;
  assign o[54] = net_sum54;
  assign o[53] = net_sum53;
  assign o[52] = net_sum52;
  assign o[51] = net_sum51;
  assign o[50] = net_sum50;
  assign o[49] = net_sum49;
  assign o[48] = net_sum48;
  assign o[47] = net_sum47;
  assign o[46] = net_sum46;
  assign o[45] = net_sum45;
  assign o[44] = net_sum44;
  assign o[43] = net_sum43;
  assign o[42] = net_sum42;
  assign o[41] = net_sum41;
  assign o[40] = net_sum40;
  assign o[39] = net_sum39;
  assign o[38] = net_sum38;
  assign o[37] = net_sum37;
  assign o[36] = net_sum36;
  assign o[35] = net_sum35;
  assign o[34] = net_sum34;
  assign o[33] = net_sum33;
  assign o[32] = net_sum32;
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_32 (
    .a(net_a32),
    .b(net_b32),
    .c(net_cout31),
    .cout(net_cout32),
    .sum(net_sum32));
  AL_FADD comp_33 (
    .a(net_a33),
    .b(net_b33),
    .c(net_cout32),
    .cout(net_cout33),
    .sum(net_sum33));
  AL_FADD comp_34 (
    .a(net_a34),
    .b(net_b34),
    .c(net_cout33),
    .cout(net_cout34),
    .sum(net_sum34));
  AL_FADD comp_35 (
    .a(net_a35),
    .b(net_b35),
    .c(net_cout34),
    .cout(net_cout35),
    .sum(net_sum35));
  AL_FADD comp_36 (
    .a(net_a36),
    .b(net_b36),
    .c(net_cout35),
    .cout(net_cout36),
    .sum(net_sum36));
  AL_FADD comp_37 (
    .a(net_a37),
    .b(net_b37),
    .c(net_cout36),
    .cout(net_cout37),
    .sum(net_sum37));
  AL_FADD comp_38 (
    .a(net_a38),
    .b(net_b38),
    .c(net_cout37),
    .cout(net_cout38),
    .sum(net_sum38));
  AL_FADD comp_39 (
    .a(net_a39),
    .b(net_b39),
    .c(net_cout38),
    .cout(net_cout39),
    .sum(net_sum39));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_40 (
    .a(net_a40),
    .b(net_b40),
    .c(net_cout39),
    .cout(net_cout40),
    .sum(net_sum40));
  AL_FADD comp_41 (
    .a(net_a41),
    .b(net_b41),
    .c(net_cout40),
    .cout(net_cout41),
    .sum(net_sum41));
  AL_FADD comp_42 (
    .a(net_a42),
    .b(net_b42),
    .c(net_cout41),
    .cout(net_cout42),
    .sum(net_sum42));
  AL_FADD comp_43 (
    .a(net_a43),
    .b(net_b43),
    .c(net_cout42),
    .cout(net_cout43),
    .sum(net_sum43));
  AL_FADD comp_44 (
    .a(net_a44),
    .b(net_b44),
    .c(net_cout43),
    .cout(net_cout44),
    .sum(net_sum44));
  AL_FADD comp_45 (
    .a(net_a45),
    .b(net_b45),
    .c(net_cout44),
    .cout(net_cout45),
    .sum(net_sum45));
  AL_FADD comp_46 (
    .a(net_a46),
    .b(net_b46),
    .c(net_cout45),
    .cout(net_cout46),
    .sum(net_sum46));
  AL_FADD comp_47 (
    .a(net_a47),
    .b(net_b47),
    .c(net_cout46),
    .cout(net_cout47),
    .sum(net_sum47));
  AL_FADD comp_48 (
    .a(net_a48),
    .b(net_b48),
    .c(net_cout47),
    .cout(net_cout48),
    .sum(net_sum48));
  AL_FADD comp_49 (
    .a(net_a49),
    .b(net_b49),
    .c(net_cout48),
    .cout(net_cout49),
    .sum(net_sum49));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_50 (
    .a(net_a50),
    .b(net_b50),
    .c(net_cout49),
    .cout(net_cout50),
    .sum(net_sum50));
  AL_FADD comp_51 (
    .a(net_a51),
    .b(net_b51),
    .c(net_cout50),
    .cout(net_cout51),
    .sum(net_sum51));
  AL_FADD comp_52 (
    .a(net_a52),
    .b(net_b52),
    .c(net_cout51),
    .cout(net_cout52),
    .sum(net_sum52));
  AL_FADD comp_53 (
    .a(net_a53),
    .b(net_b53),
    .c(net_cout52),
    .cout(net_cout53),
    .sum(net_sum53));
  AL_FADD comp_54 (
    .a(net_a54),
    .b(net_b54),
    .c(net_cout53),
    .cout(net_cout54),
    .sum(net_sum54));
  AL_FADD comp_55 (
    .a(net_a55),
    .b(net_b55),
    .c(net_cout54),
    .cout(net_cout55),
    .sum(net_sum55));
  AL_FADD comp_56 (
    .a(net_a56),
    .b(net_b56),
    .c(net_cout55),
    .cout(net_cout56),
    .sum(net_sum56));
  AL_FADD comp_57 (
    .a(net_a57),
    .b(net_b57),
    .c(net_cout56),
    .cout(net_cout57),
    .sum(net_sum57));
  AL_FADD comp_58 (
    .a(net_a58),
    .b(net_b58),
    .c(net_cout57),
    .cout(net_cout58),
    .sum(net_sum58));
  AL_FADD comp_59 (
    .a(net_a59),
    .b(net_b59),
    .c(net_cout58),
    .cout(net_cout59),
    .sum(net_sum59));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w12
  (
  i0,
  i1,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  output o;

  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[6]_i1[6_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_xor_i0[0]_i_o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[6]_i1[6_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_or_xor_i0[6]_i1[6  (\or_or_xor_i0[6]_i1[6_o , \or_xor_i0[6]_i1[6]_o_o , \or_xor_i0[9]_i1[9]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \or_xor_i0[4]_i1[4]_o_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \or_xor_i0[7]_i1[7]_o_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \or_xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module add_pu62_pu62_o62
  (
  i0,
  i1,
  o
  );

  input [61:0] i0;
  input [61:0] i1;
  output [61:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a32;
  wire net_a33;
  wire net_a34;
  wire net_a35;
  wire net_a36;
  wire net_a37;
  wire net_a38;
  wire net_a39;
  wire net_a4;
  wire net_a40;
  wire net_a41;
  wire net_a42;
  wire net_a43;
  wire net_a44;
  wire net_a45;
  wire net_a46;
  wire net_a47;
  wire net_a48;
  wire net_a49;
  wire net_a5;
  wire net_a50;
  wire net_a51;
  wire net_a52;
  wire net_a53;
  wire net_a54;
  wire net_a55;
  wire net_a56;
  wire net_a57;
  wire net_a58;
  wire net_a59;
  wire net_a6;
  wire net_a60;
  wire net_a61;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b32;
  wire net_b33;
  wire net_b34;
  wire net_b35;
  wire net_b36;
  wire net_b37;
  wire net_b38;
  wire net_b39;
  wire net_b4;
  wire net_b40;
  wire net_b41;
  wire net_b42;
  wire net_b43;
  wire net_b44;
  wire net_b45;
  wire net_b46;
  wire net_b47;
  wire net_b48;
  wire net_b49;
  wire net_b5;
  wire net_b50;
  wire net_b51;
  wire net_b52;
  wire net_b53;
  wire net_b54;
  wire net_b55;
  wire net_b56;
  wire net_b57;
  wire net_b58;
  wire net_b59;
  wire net_b6;
  wire net_b60;
  wire net_b61;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout32;
  wire net_cout33;
  wire net_cout34;
  wire net_cout35;
  wire net_cout36;
  wire net_cout37;
  wire net_cout38;
  wire net_cout39;
  wire net_cout4;
  wire net_cout40;
  wire net_cout41;
  wire net_cout42;
  wire net_cout43;
  wire net_cout44;
  wire net_cout45;
  wire net_cout46;
  wire net_cout47;
  wire net_cout48;
  wire net_cout49;
  wire net_cout5;
  wire net_cout50;
  wire net_cout51;
  wire net_cout52;
  wire net_cout53;
  wire net_cout54;
  wire net_cout55;
  wire net_cout56;
  wire net_cout57;
  wire net_cout58;
  wire net_cout59;
  wire net_cout6;
  wire net_cout60;
  wire net_cout61;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum32;
  wire net_sum33;
  wire net_sum34;
  wire net_sum35;
  wire net_sum36;
  wire net_sum37;
  wire net_sum38;
  wire net_sum39;
  wire net_sum4;
  wire net_sum40;
  wire net_sum41;
  wire net_sum42;
  wire net_sum43;
  wire net_sum44;
  wire net_sum45;
  wire net_sum46;
  wire net_sum47;
  wire net_sum48;
  wire net_sum49;
  wire net_sum5;
  wire net_sum50;
  wire net_sum51;
  wire net_sum52;
  wire net_sum53;
  wire net_sum54;
  wire net_sum55;
  wire net_sum56;
  wire net_sum57;
  wire net_sum58;
  wire net_sum59;
  wire net_sum6;
  wire net_sum60;
  wire net_sum61;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a61 = i0[61];
  assign net_a60 = i0[60];
  assign net_a59 = i0[59];
  assign net_a58 = i0[58];
  assign net_a57 = i0[57];
  assign net_a56 = i0[56];
  assign net_a55 = i0[55];
  assign net_a54 = i0[54];
  assign net_a53 = i0[53];
  assign net_a52 = i0[52];
  assign net_a51 = i0[51];
  assign net_a50 = i0[50];
  assign net_a49 = i0[49];
  assign net_a48 = i0[48];
  assign net_a47 = i0[47];
  assign net_a46 = i0[46];
  assign net_a45 = i0[45];
  assign net_a44 = i0[44];
  assign net_a43 = i0[43];
  assign net_a42 = i0[42];
  assign net_a41 = i0[41];
  assign net_a40 = i0[40];
  assign net_a39 = i0[39];
  assign net_a38 = i0[38];
  assign net_a37 = i0[37];
  assign net_a36 = i0[36];
  assign net_a35 = i0[35];
  assign net_a34 = i0[34];
  assign net_a33 = i0[33];
  assign net_a32 = i0[32];
  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b61 = i1[61];
  assign net_b60 = i1[60];
  assign net_b59 = i1[59];
  assign net_b58 = i1[58];
  assign net_b57 = i1[57];
  assign net_b56 = i1[56];
  assign net_b55 = i1[55];
  assign net_b54 = i1[54];
  assign net_b53 = i1[53];
  assign net_b52 = i1[52];
  assign net_b51 = i1[51];
  assign net_b50 = i1[50];
  assign net_b49 = i1[49];
  assign net_b48 = i1[48];
  assign net_b47 = i1[47];
  assign net_b46 = i1[46];
  assign net_b45 = i1[45];
  assign net_b44 = i1[44];
  assign net_b43 = i1[43];
  assign net_b42 = i1[42];
  assign net_b41 = i1[41];
  assign net_b40 = i1[40];
  assign net_b39 = i1[39];
  assign net_b38 = i1[38];
  assign net_b37 = i1[37];
  assign net_b36 = i1[36];
  assign net_b35 = i1[35];
  assign net_b34 = i1[34];
  assign net_b33 = i1[33];
  assign net_b32 = i1[32];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[61] = net_sum61;
  assign o[60] = net_sum60;
  assign o[59] = net_sum59;
  assign o[58] = net_sum58;
  assign o[57] = net_sum57;
  assign o[56] = net_sum56;
  assign o[55] = net_sum55;
  assign o[54] = net_sum54;
  assign o[53] = net_sum53;
  assign o[52] = net_sum52;
  assign o[51] = net_sum51;
  assign o[50] = net_sum50;
  assign o[49] = net_sum49;
  assign o[48] = net_sum48;
  assign o[47] = net_sum47;
  assign o[46] = net_sum46;
  assign o[45] = net_sum45;
  assign o[44] = net_sum44;
  assign o[43] = net_sum43;
  assign o[42] = net_sum42;
  assign o[41] = net_sum41;
  assign o[40] = net_sum40;
  assign o[39] = net_sum39;
  assign o[38] = net_sum38;
  assign o[37] = net_sum37;
  assign o[36] = net_sum36;
  assign o[35] = net_sum35;
  assign o[34] = net_sum34;
  assign o[33] = net_sum33;
  assign o[32] = net_sum32;
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_32 (
    .a(net_a32),
    .b(net_b32),
    .c(net_cout31),
    .cout(net_cout32),
    .sum(net_sum32));
  AL_FADD comp_33 (
    .a(net_a33),
    .b(net_b33),
    .c(net_cout32),
    .cout(net_cout33),
    .sum(net_sum33));
  AL_FADD comp_34 (
    .a(net_a34),
    .b(net_b34),
    .c(net_cout33),
    .cout(net_cout34),
    .sum(net_sum34));
  AL_FADD comp_35 (
    .a(net_a35),
    .b(net_b35),
    .c(net_cout34),
    .cout(net_cout35),
    .sum(net_sum35));
  AL_FADD comp_36 (
    .a(net_a36),
    .b(net_b36),
    .c(net_cout35),
    .cout(net_cout36),
    .sum(net_sum36));
  AL_FADD comp_37 (
    .a(net_a37),
    .b(net_b37),
    .c(net_cout36),
    .cout(net_cout37),
    .sum(net_sum37));
  AL_FADD comp_38 (
    .a(net_a38),
    .b(net_b38),
    .c(net_cout37),
    .cout(net_cout38),
    .sum(net_sum38));
  AL_FADD comp_39 (
    .a(net_a39),
    .b(net_b39),
    .c(net_cout38),
    .cout(net_cout39),
    .sum(net_sum39));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_40 (
    .a(net_a40),
    .b(net_b40),
    .c(net_cout39),
    .cout(net_cout40),
    .sum(net_sum40));
  AL_FADD comp_41 (
    .a(net_a41),
    .b(net_b41),
    .c(net_cout40),
    .cout(net_cout41),
    .sum(net_sum41));
  AL_FADD comp_42 (
    .a(net_a42),
    .b(net_b42),
    .c(net_cout41),
    .cout(net_cout42),
    .sum(net_sum42));
  AL_FADD comp_43 (
    .a(net_a43),
    .b(net_b43),
    .c(net_cout42),
    .cout(net_cout43),
    .sum(net_sum43));
  AL_FADD comp_44 (
    .a(net_a44),
    .b(net_b44),
    .c(net_cout43),
    .cout(net_cout44),
    .sum(net_sum44));
  AL_FADD comp_45 (
    .a(net_a45),
    .b(net_b45),
    .c(net_cout44),
    .cout(net_cout45),
    .sum(net_sum45));
  AL_FADD comp_46 (
    .a(net_a46),
    .b(net_b46),
    .c(net_cout45),
    .cout(net_cout46),
    .sum(net_sum46));
  AL_FADD comp_47 (
    .a(net_a47),
    .b(net_b47),
    .c(net_cout46),
    .cout(net_cout47),
    .sum(net_sum47));
  AL_FADD comp_48 (
    .a(net_a48),
    .b(net_b48),
    .c(net_cout47),
    .cout(net_cout48),
    .sum(net_sum48));
  AL_FADD comp_49 (
    .a(net_a49),
    .b(net_b49),
    .c(net_cout48),
    .cout(net_cout49),
    .sum(net_sum49));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_50 (
    .a(net_a50),
    .b(net_b50),
    .c(net_cout49),
    .cout(net_cout50),
    .sum(net_sum50));
  AL_FADD comp_51 (
    .a(net_a51),
    .b(net_b51),
    .c(net_cout50),
    .cout(net_cout51),
    .sum(net_sum51));
  AL_FADD comp_52 (
    .a(net_a52),
    .b(net_b52),
    .c(net_cout51),
    .cout(net_cout52),
    .sum(net_sum52));
  AL_FADD comp_53 (
    .a(net_a53),
    .b(net_b53),
    .c(net_cout52),
    .cout(net_cout53),
    .sum(net_sum53));
  AL_FADD comp_54 (
    .a(net_a54),
    .b(net_b54),
    .c(net_cout53),
    .cout(net_cout54),
    .sum(net_sum54));
  AL_FADD comp_55 (
    .a(net_a55),
    .b(net_b55),
    .c(net_cout54),
    .cout(net_cout55),
    .sum(net_sum55));
  AL_FADD comp_56 (
    .a(net_a56),
    .b(net_b56),
    .c(net_cout55),
    .cout(net_cout56),
    .sum(net_sum56));
  AL_FADD comp_57 (
    .a(net_a57),
    .b(net_b57),
    .c(net_cout56),
    .cout(net_cout57),
    .sum(net_sum57));
  AL_FADD comp_58 (
    .a(net_a58),
    .b(net_b58),
    .c(net_cout57),
    .cout(net_cout58),
    .sum(net_sum58));
  AL_FADD comp_59 (
    .a(net_a59),
    .b(net_b59),
    .c(net_cout58),
    .cout(net_cout59),
    .sum(net_sum59));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_60 (
    .a(net_a60),
    .b(net_b60),
    .c(net_cout59),
    .cout(net_cout60),
    .sum(net_sum60));
  AL_FADD comp_61 (
    .a(net_a61),
    .b(net_b61),
    .c(net_cout60),
    .cout(net_cout61),
    .sum(net_sum61));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module ne_w5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output o;

  wire [4:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3], diff[4]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);

endmodule 

module add_pu5_mu5_o5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output [4:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_nb0;
  wire net_nb1;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;

  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);

endmodule 

module add_pu32_pu32_o32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [31:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module lt_u64_u64
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [63:0] i0;
  input [63:0] i1;
  output o;

  wire [63:0] diff;
  wire diff_12_18;
  wire diff_19_26;
  wire diff_27_35;
  wire diff_36_45;
  wire diff_46_56;
  wire diff_57_63;
  wire diff_6_11;
  wire less_12_18;
  wire \less_12_18_inst/diff_0 ;
  wire \less_12_18_inst/diff_1 ;
  wire \less_12_18_inst/diff_2 ;
  wire \less_12_18_inst/diff_3 ;
  wire \less_12_18_inst/diff_4 ;
  wire \less_12_18_inst/diff_5 ;
  wire \less_12_18_inst/diff_6 ;
  wire \less_12_18_inst/o_0 ;
  wire \less_12_18_inst/o_1 ;
  wire \less_12_18_inst/o_2 ;
  wire \less_12_18_inst/o_3 ;
  wire \less_12_18_inst/o_4 ;
  wire \less_12_18_inst/o_5 ;
  wire less_19_26;
  wire \less_19_26_inst/diff_0 ;
  wire \less_19_26_inst/diff_1 ;
  wire \less_19_26_inst/diff_2 ;
  wire \less_19_26_inst/diff_3 ;
  wire \less_19_26_inst/diff_4 ;
  wire \less_19_26_inst/diff_5 ;
  wire \less_19_26_inst/diff_6 ;
  wire \less_19_26_inst/diff_7 ;
  wire \less_19_26_inst/o_0 ;
  wire \less_19_26_inst/o_1 ;
  wire \less_19_26_inst/o_2 ;
  wire \less_19_26_inst/o_3 ;
  wire \less_19_26_inst/o_4 ;
  wire \less_19_26_inst/o_5 ;
  wire \less_19_26_inst/o_6 ;
  wire less_27_35;
  wire \less_27_35_inst/diff_0 ;
  wire \less_27_35_inst/diff_1 ;
  wire \less_27_35_inst/diff_2 ;
  wire \less_27_35_inst/diff_3 ;
  wire \less_27_35_inst/diff_4 ;
  wire \less_27_35_inst/diff_5 ;
  wire \less_27_35_inst/diff_6 ;
  wire \less_27_35_inst/diff_7 ;
  wire \less_27_35_inst/diff_8 ;
  wire \less_27_35_inst/o_0 ;
  wire \less_27_35_inst/o_1 ;
  wire \less_27_35_inst/o_2 ;
  wire \less_27_35_inst/o_3 ;
  wire \less_27_35_inst/o_4 ;
  wire \less_27_35_inst/o_5 ;
  wire \less_27_35_inst/o_6 ;
  wire \less_27_35_inst/o_7 ;
  wire less_36_45;
  wire \less_36_45_inst/diff_0 ;
  wire \less_36_45_inst/diff_1 ;
  wire \less_36_45_inst/diff_2 ;
  wire \less_36_45_inst/diff_3 ;
  wire \less_36_45_inst/diff_4 ;
  wire \less_36_45_inst/diff_5 ;
  wire \less_36_45_inst/diff_6 ;
  wire \less_36_45_inst/diff_7 ;
  wire \less_36_45_inst/diff_8 ;
  wire \less_36_45_inst/diff_9 ;
  wire \less_36_45_inst/o_0 ;
  wire \less_36_45_inst/o_1 ;
  wire \less_36_45_inst/o_2 ;
  wire \less_36_45_inst/o_3 ;
  wire \less_36_45_inst/o_4 ;
  wire \less_36_45_inst/o_5 ;
  wire \less_36_45_inst/o_6 ;
  wire \less_36_45_inst/o_7 ;
  wire \less_36_45_inst/o_8 ;
  wire less_46_56;
  wire \less_46_56_inst/diff_0 ;
  wire \less_46_56_inst/diff_1 ;
  wire \less_46_56_inst/diff_10 ;
  wire \less_46_56_inst/diff_2 ;
  wire \less_46_56_inst/diff_3 ;
  wire \less_46_56_inst/diff_4 ;
  wire \less_46_56_inst/diff_5 ;
  wire \less_46_56_inst/diff_6 ;
  wire \less_46_56_inst/diff_7 ;
  wire \less_46_56_inst/diff_8 ;
  wire \less_46_56_inst/diff_9 ;
  wire \less_46_56_inst/o_0 ;
  wire \less_46_56_inst/o_1 ;
  wire \less_46_56_inst/o_2 ;
  wire \less_46_56_inst/o_3 ;
  wire \less_46_56_inst/o_4 ;
  wire \less_46_56_inst/o_5 ;
  wire \less_46_56_inst/o_6 ;
  wire \less_46_56_inst/o_7 ;
  wire \less_46_56_inst/o_8 ;
  wire \less_46_56_inst/o_9 ;
  wire less_57_63;
  wire \less_57_63_inst/diff_0 ;
  wire \less_57_63_inst/diff_1 ;
  wire \less_57_63_inst/diff_2 ;
  wire \less_57_63_inst/diff_3 ;
  wire \less_57_63_inst/diff_4 ;
  wire \less_57_63_inst/diff_5 ;
  wire \less_57_63_inst/diff_6 ;
  wire \less_57_63_inst/o_0 ;
  wire \less_57_63_inst/o_1 ;
  wire \less_57_63_inst/o_2 ;
  wire \less_57_63_inst/o_3 ;
  wire \less_57_63_inst/o_4 ;
  wire \less_57_63_inst/o_5 ;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_10;
  wire o_11;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;
  wire o_6;
  wire o_7;
  wire o_8;
  wire o_9;

  or any_diff_12_18 (diff_12_18, diff[12], diff[13], diff[14], diff[15], diff[16], diff[17], diff[18]);
  or any_diff_19_26 (diff_19_26, diff[19], diff[20], diff[21], diff[22], diff[23], diff[24], diff[25], diff[26]);
  or any_diff_27_35 (diff_27_35, diff[27], diff[28], diff[29], diff[30], diff[31], diff[32], diff[33], diff[34], diff[35]);
  or any_diff_36_45 (diff_36_45, diff[36], diff[37], diff[38], diff[39], diff[40], diff[41], diff[42], diff[43], diff[44], diff[45]);
  or any_diff_46_56 (diff_46_56, diff[46], diff[47], diff[48], diff[49], diff[50], diff[51], diff[52], diff[53], diff[54], diff[55], diff[56]);
  or any_diff_57_63 (diff_57_63, diff[57], diff[58], diff[59], diff[60], diff[61], diff[62], diff[63]);
  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_13 (diff[13], i0[13], i1[13]);
  xor diff_14 (diff[14], i0[14], i1[14]);
  xor diff_15 (diff[15], i0[15], i1[15]);
  xor diff_16 (diff[16], i0[16], i1[16]);
  xor diff_17 (diff[17], i0[17], i1[17]);
  xor diff_18 (diff[18], i0[18], i1[18]);
  xor diff_19 (diff[19], i0[19], i1[19]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_20 (diff[20], i0[20], i1[20]);
  xor diff_21 (diff[21], i0[21], i1[21]);
  xor diff_22 (diff[22], i0[22], i1[22]);
  xor diff_23 (diff[23], i0[23], i1[23]);
  xor diff_24 (diff[24], i0[24], i1[24]);
  xor diff_25 (diff[25], i0[25], i1[25]);
  xor diff_26 (diff[26], i0[26], i1[26]);
  xor diff_27 (diff[27], i0[27], i1[27]);
  xor diff_28 (diff[28], i0[28], i1[28]);
  xor diff_29 (diff[29], i0[29], i1[29]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_30 (diff[30], i0[30], i1[30]);
  xor diff_31 (diff[31], i0[31], i1[31]);
  xor diff_32 (diff[32], i0[32], i1[32]);
  xor diff_33 (diff[33], i0[33], i1[33]);
  xor diff_34 (diff[34], i0[34], i1[34]);
  xor diff_35 (diff[35], i0[35], i1[35]);
  xor diff_36 (diff[36], i0[36], i1[36]);
  xor diff_37 (diff[37], i0[37], i1[37]);
  xor diff_38 (diff[38], i0[38], i1[38]);
  xor diff_39 (diff[39], i0[39], i1[39]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_40 (diff[40], i0[40], i1[40]);
  xor diff_41 (diff[41], i0[41], i1[41]);
  xor diff_42 (diff[42], i0[42], i1[42]);
  xor diff_43 (diff[43], i0[43], i1[43]);
  xor diff_44 (diff[44], i0[44], i1[44]);
  xor diff_45 (diff[45], i0[45], i1[45]);
  xor diff_46 (diff[46], i0[46], i1[46]);
  xor diff_47 (diff[47], i0[47], i1[47]);
  xor diff_48 (diff[48], i0[48], i1[48]);
  xor diff_49 (diff[49], i0[49], i1[49]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_50 (diff[50], i0[50], i1[50]);
  xor diff_51 (diff[51], i0[51], i1[51]);
  xor diff_52 (diff[52], i0[52], i1[52]);
  xor diff_53 (diff[53], i0[53], i1[53]);
  xor diff_54 (diff[54], i0[54], i1[54]);
  xor diff_55 (diff[55], i0[55], i1[55]);
  xor diff_56 (diff[56], i0[56], i1[56]);
  xor diff_57 (diff[57], i0[57], i1[57]);
  xor diff_58 (diff[58], i0[58], i1[58]);
  xor diff_59 (diff[59], i0[59], i1[59]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_60 (diff[60], i0[60], i1[60]);
  xor diff_61 (diff[61], i0[61], i1[61]);
  xor diff_62 (diff[62], i0[62], i1[62]);
  xor diff_63 (diff[63], i0[63], i1[63]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_12_18_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[12]),
    .sel(\less_12_18_inst/diff_0 ),
    .o(\less_12_18_inst/o_0 ));
  AL_MUX \less_12_18_inst/mux_1  (
    .i0(\less_12_18_inst/o_0 ),
    .i1(i1[13]),
    .sel(\less_12_18_inst/diff_1 ),
    .o(\less_12_18_inst/o_1 ));
  AL_MUX \less_12_18_inst/mux_2  (
    .i0(\less_12_18_inst/o_1 ),
    .i1(i1[14]),
    .sel(\less_12_18_inst/diff_2 ),
    .o(\less_12_18_inst/o_2 ));
  AL_MUX \less_12_18_inst/mux_3  (
    .i0(\less_12_18_inst/o_2 ),
    .i1(i1[15]),
    .sel(\less_12_18_inst/diff_3 ),
    .o(\less_12_18_inst/o_3 ));
  AL_MUX \less_12_18_inst/mux_4  (
    .i0(\less_12_18_inst/o_3 ),
    .i1(i1[16]),
    .sel(\less_12_18_inst/diff_4 ),
    .o(\less_12_18_inst/o_4 ));
  AL_MUX \less_12_18_inst/mux_5  (
    .i0(\less_12_18_inst/o_4 ),
    .i1(i1[17]),
    .sel(\less_12_18_inst/diff_5 ),
    .o(\less_12_18_inst/o_5 ));
  AL_MUX \less_12_18_inst/mux_6  (
    .i0(\less_12_18_inst/o_5 ),
    .i1(i1[18]),
    .sel(\less_12_18_inst/diff_6 ),
    .o(less_12_18));
  xor \less_12_18_inst/xor_0  (\less_12_18_inst/diff_0 , i0[12], i1[12]);
  xor \less_12_18_inst/xor_1  (\less_12_18_inst/diff_1 , i0[13], i1[13]);
  xor \less_12_18_inst/xor_2  (\less_12_18_inst/diff_2 , i0[14], i1[14]);
  xor \less_12_18_inst/xor_3  (\less_12_18_inst/diff_3 , i0[15], i1[15]);
  xor \less_12_18_inst/xor_4  (\less_12_18_inst/diff_4 , i0[16], i1[16]);
  xor \less_12_18_inst/xor_5  (\less_12_18_inst/diff_5 , i0[17], i1[17]);
  xor \less_12_18_inst/xor_6  (\less_12_18_inst/diff_6 , i0[18], i1[18]);
  AL_MUX \less_19_26_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[19]),
    .sel(\less_19_26_inst/diff_0 ),
    .o(\less_19_26_inst/o_0 ));
  AL_MUX \less_19_26_inst/mux_1  (
    .i0(\less_19_26_inst/o_0 ),
    .i1(i1[20]),
    .sel(\less_19_26_inst/diff_1 ),
    .o(\less_19_26_inst/o_1 ));
  AL_MUX \less_19_26_inst/mux_2  (
    .i0(\less_19_26_inst/o_1 ),
    .i1(i1[21]),
    .sel(\less_19_26_inst/diff_2 ),
    .o(\less_19_26_inst/o_2 ));
  AL_MUX \less_19_26_inst/mux_3  (
    .i0(\less_19_26_inst/o_2 ),
    .i1(i1[22]),
    .sel(\less_19_26_inst/diff_3 ),
    .o(\less_19_26_inst/o_3 ));
  AL_MUX \less_19_26_inst/mux_4  (
    .i0(\less_19_26_inst/o_3 ),
    .i1(i1[23]),
    .sel(\less_19_26_inst/diff_4 ),
    .o(\less_19_26_inst/o_4 ));
  AL_MUX \less_19_26_inst/mux_5  (
    .i0(\less_19_26_inst/o_4 ),
    .i1(i1[24]),
    .sel(\less_19_26_inst/diff_5 ),
    .o(\less_19_26_inst/o_5 ));
  AL_MUX \less_19_26_inst/mux_6  (
    .i0(\less_19_26_inst/o_5 ),
    .i1(i1[25]),
    .sel(\less_19_26_inst/diff_6 ),
    .o(\less_19_26_inst/o_6 ));
  AL_MUX \less_19_26_inst/mux_7  (
    .i0(\less_19_26_inst/o_6 ),
    .i1(i1[26]),
    .sel(\less_19_26_inst/diff_7 ),
    .o(less_19_26));
  xor \less_19_26_inst/xor_0  (\less_19_26_inst/diff_0 , i0[19], i1[19]);
  xor \less_19_26_inst/xor_1  (\less_19_26_inst/diff_1 , i0[20], i1[20]);
  xor \less_19_26_inst/xor_2  (\less_19_26_inst/diff_2 , i0[21], i1[21]);
  xor \less_19_26_inst/xor_3  (\less_19_26_inst/diff_3 , i0[22], i1[22]);
  xor \less_19_26_inst/xor_4  (\less_19_26_inst/diff_4 , i0[23], i1[23]);
  xor \less_19_26_inst/xor_5  (\less_19_26_inst/diff_5 , i0[24], i1[24]);
  xor \less_19_26_inst/xor_6  (\less_19_26_inst/diff_6 , i0[25], i1[25]);
  xor \less_19_26_inst/xor_7  (\less_19_26_inst/diff_7 , i0[26], i1[26]);
  AL_MUX \less_27_35_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[27]),
    .sel(\less_27_35_inst/diff_0 ),
    .o(\less_27_35_inst/o_0 ));
  AL_MUX \less_27_35_inst/mux_1  (
    .i0(\less_27_35_inst/o_0 ),
    .i1(i1[28]),
    .sel(\less_27_35_inst/diff_1 ),
    .o(\less_27_35_inst/o_1 ));
  AL_MUX \less_27_35_inst/mux_2  (
    .i0(\less_27_35_inst/o_1 ),
    .i1(i1[29]),
    .sel(\less_27_35_inst/diff_2 ),
    .o(\less_27_35_inst/o_2 ));
  AL_MUX \less_27_35_inst/mux_3  (
    .i0(\less_27_35_inst/o_2 ),
    .i1(i1[30]),
    .sel(\less_27_35_inst/diff_3 ),
    .o(\less_27_35_inst/o_3 ));
  AL_MUX \less_27_35_inst/mux_4  (
    .i0(\less_27_35_inst/o_3 ),
    .i1(i1[31]),
    .sel(\less_27_35_inst/diff_4 ),
    .o(\less_27_35_inst/o_4 ));
  AL_MUX \less_27_35_inst/mux_5  (
    .i0(\less_27_35_inst/o_4 ),
    .i1(i1[32]),
    .sel(\less_27_35_inst/diff_5 ),
    .o(\less_27_35_inst/o_5 ));
  AL_MUX \less_27_35_inst/mux_6  (
    .i0(\less_27_35_inst/o_5 ),
    .i1(i1[33]),
    .sel(\less_27_35_inst/diff_6 ),
    .o(\less_27_35_inst/o_6 ));
  AL_MUX \less_27_35_inst/mux_7  (
    .i0(\less_27_35_inst/o_6 ),
    .i1(i1[34]),
    .sel(\less_27_35_inst/diff_7 ),
    .o(\less_27_35_inst/o_7 ));
  AL_MUX \less_27_35_inst/mux_8  (
    .i0(\less_27_35_inst/o_7 ),
    .i1(i1[35]),
    .sel(\less_27_35_inst/diff_8 ),
    .o(less_27_35));
  xor \less_27_35_inst/xor_0  (\less_27_35_inst/diff_0 , i0[27], i1[27]);
  xor \less_27_35_inst/xor_1  (\less_27_35_inst/diff_1 , i0[28], i1[28]);
  xor \less_27_35_inst/xor_2  (\less_27_35_inst/diff_2 , i0[29], i1[29]);
  xor \less_27_35_inst/xor_3  (\less_27_35_inst/diff_3 , i0[30], i1[30]);
  xor \less_27_35_inst/xor_4  (\less_27_35_inst/diff_4 , i0[31], i1[31]);
  xor \less_27_35_inst/xor_5  (\less_27_35_inst/diff_5 , i0[32], i1[32]);
  xor \less_27_35_inst/xor_6  (\less_27_35_inst/diff_6 , i0[33], i1[33]);
  xor \less_27_35_inst/xor_7  (\less_27_35_inst/diff_7 , i0[34], i1[34]);
  xor \less_27_35_inst/xor_8  (\less_27_35_inst/diff_8 , i0[35], i1[35]);
  AL_MUX \less_36_45_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[36]),
    .sel(\less_36_45_inst/diff_0 ),
    .o(\less_36_45_inst/o_0 ));
  AL_MUX \less_36_45_inst/mux_1  (
    .i0(\less_36_45_inst/o_0 ),
    .i1(i1[37]),
    .sel(\less_36_45_inst/diff_1 ),
    .o(\less_36_45_inst/o_1 ));
  AL_MUX \less_36_45_inst/mux_2  (
    .i0(\less_36_45_inst/o_1 ),
    .i1(i1[38]),
    .sel(\less_36_45_inst/diff_2 ),
    .o(\less_36_45_inst/o_2 ));
  AL_MUX \less_36_45_inst/mux_3  (
    .i0(\less_36_45_inst/o_2 ),
    .i1(i1[39]),
    .sel(\less_36_45_inst/diff_3 ),
    .o(\less_36_45_inst/o_3 ));
  AL_MUX \less_36_45_inst/mux_4  (
    .i0(\less_36_45_inst/o_3 ),
    .i1(i1[40]),
    .sel(\less_36_45_inst/diff_4 ),
    .o(\less_36_45_inst/o_4 ));
  AL_MUX \less_36_45_inst/mux_5  (
    .i0(\less_36_45_inst/o_4 ),
    .i1(i1[41]),
    .sel(\less_36_45_inst/diff_5 ),
    .o(\less_36_45_inst/o_5 ));
  AL_MUX \less_36_45_inst/mux_6  (
    .i0(\less_36_45_inst/o_5 ),
    .i1(i1[42]),
    .sel(\less_36_45_inst/diff_6 ),
    .o(\less_36_45_inst/o_6 ));
  AL_MUX \less_36_45_inst/mux_7  (
    .i0(\less_36_45_inst/o_6 ),
    .i1(i1[43]),
    .sel(\less_36_45_inst/diff_7 ),
    .o(\less_36_45_inst/o_7 ));
  AL_MUX \less_36_45_inst/mux_8  (
    .i0(\less_36_45_inst/o_7 ),
    .i1(i1[44]),
    .sel(\less_36_45_inst/diff_8 ),
    .o(\less_36_45_inst/o_8 ));
  AL_MUX \less_36_45_inst/mux_9  (
    .i0(\less_36_45_inst/o_8 ),
    .i1(i1[45]),
    .sel(\less_36_45_inst/diff_9 ),
    .o(less_36_45));
  xor \less_36_45_inst/xor_0  (\less_36_45_inst/diff_0 , i0[36], i1[36]);
  xor \less_36_45_inst/xor_1  (\less_36_45_inst/diff_1 , i0[37], i1[37]);
  xor \less_36_45_inst/xor_2  (\less_36_45_inst/diff_2 , i0[38], i1[38]);
  xor \less_36_45_inst/xor_3  (\less_36_45_inst/diff_3 , i0[39], i1[39]);
  xor \less_36_45_inst/xor_4  (\less_36_45_inst/diff_4 , i0[40], i1[40]);
  xor \less_36_45_inst/xor_5  (\less_36_45_inst/diff_5 , i0[41], i1[41]);
  xor \less_36_45_inst/xor_6  (\less_36_45_inst/diff_6 , i0[42], i1[42]);
  xor \less_36_45_inst/xor_7  (\less_36_45_inst/diff_7 , i0[43], i1[43]);
  xor \less_36_45_inst/xor_8  (\less_36_45_inst/diff_8 , i0[44], i1[44]);
  xor \less_36_45_inst/xor_9  (\less_36_45_inst/diff_9 , i0[45], i1[45]);
  AL_MUX \less_46_56_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[46]),
    .sel(\less_46_56_inst/diff_0 ),
    .o(\less_46_56_inst/o_0 ));
  AL_MUX \less_46_56_inst/mux_1  (
    .i0(\less_46_56_inst/o_0 ),
    .i1(i1[47]),
    .sel(\less_46_56_inst/diff_1 ),
    .o(\less_46_56_inst/o_1 ));
  AL_MUX \less_46_56_inst/mux_10  (
    .i0(\less_46_56_inst/o_9 ),
    .i1(i1[56]),
    .sel(\less_46_56_inst/diff_10 ),
    .o(less_46_56));
  AL_MUX \less_46_56_inst/mux_2  (
    .i0(\less_46_56_inst/o_1 ),
    .i1(i1[48]),
    .sel(\less_46_56_inst/diff_2 ),
    .o(\less_46_56_inst/o_2 ));
  AL_MUX \less_46_56_inst/mux_3  (
    .i0(\less_46_56_inst/o_2 ),
    .i1(i1[49]),
    .sel(\less_46_56_inst/diff_3 ),
    .o(\less_46_56_inst/o_3 ));
  AL_MUX \less_46_56_inst/mux_4  (
    .i0(\less_46_56_inst/o_3 ),
    .i1(i1[50]),
    .sel(\less_46_56_inst/diff_4 ),
    .o(\less_46_56_inst/o_4 ));
  AL_MUX \less_46_56_inst/mux_5  (
    .i0(\less_46_56_inst/o_4 ),
    .i1(i1[51]),
    .sel(\less_46_56_inst/diff_5 ),
    .o(\less_46_56_inst/o_5 ));
  AL_MUX \less_46_56_inst/mux_6  (
    .i0(\less_46_56_inst/o_5 ),
    .i1(i1[52]),
    .sel(\less_46_56_inst/diff_6 ),
    .o(\less_46_56_inst/o_6 ));
  AL_MUX \less_46_56_inst/mux_7  (
    .i0(\less_46_56_inst/o_6 ),
    .i1(i1[53]),
    .sel(\less_46_56_inst/diff_7 ),
    .o(\less_46_56_inst/o_7 ));
  AL_MUX \less_46_56_inst/mux_8  (
    .i0(\less_46_56_inst/o_7 ),
    .i1(i1[54]),
    .sel(\less_46_56_inst/diff_8 ),
    .o(\less_46_56_inst/o_8 ));
  AL_MUX \less_46_56_inst/mux_9  (
    .i0(\less_46_56_inst/o_8 ),
    .i1(i1[55]),
    .sel(\less_46_56_inst/diff_9 ),
    .o(\less_46_56_inst/o_9 ));
  xor \less_46_56_inst/xor_0  (\less_46_56_inst/diff_0 , i0[46], i1[46]);
  xor \less_46_56_inst/xor_1  (\less_46_56_inst/diff_1 , i0[47], i1[47]);
  xor \less_46_56_inst/xor_10  (\less_46_56_inst/diff_10 , i0[56], i1[56]);
  xor \less_46_56_inst/xor_2  (\less_46_56_inst/diff_2 , i0[48], i1[48]);
  xor \less_46_56_inst/xor_3  (\less_46_56_inst/diff_3 , i0[49], i1[49]);
  xor \less_46_56_inst/xor_4  (\less_46_56_inst/diff_4 , i0[50], i1[50]);
  xor \less_46_56_inst/xor_5  (\less_46_56_inst/diff_5 , i0[51], i1[51]);
  xor \less_46_56_inst/xor_6  (\less_46_56_inst/diff_6 , i0[52], i1[52]);
  xor \less_46_56_inst/xor_7  (\less_46_56_inst/diff_7 , i0[53], i1[53]);
  xor \less_46_56_inst/xor_8  (\less_46_56_inst/diff_8 , i0[54], i1[54]);
  xor \less_46_56_inst/xor_9  (\less_46_56_inst/diff_9 , i0[55], i1[55]);
  AL_MUX \less_57_63_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[57]),
    .sel(\less_57_63_inst/diff_0 ),
    .o(\less_57_63_inst/o_0 ));
  AL_MUX \less_57_63_inst/mux_1  (
    .i0(\less_57_63_inst/o_0 ),
    .i1(i1[58]),
    .sel(\less_57_63_inst/diff_1 ),
    .o(\less_57_63_inst/o_1 ));
  AL_MUX \less_57_63_inst/mux_2  (
    .i0(\less_57_63_inst/o_1 ),
    .i1(i1[59]),
    .sel(\less_57_63_inst/diff_2 ),
    .o(\less_57_63_inst/o_2 ));
  AL_MUX \less_57_63_inst/mux_3  (
    .i0(\less_57_63_inst/o_2 ),
    .i1(i1[60]),
    .sel(\less_57_63_inst/diff_3 ),
    .o(\less_57_63_inst/o_3 ));
  AL_MUX \less_57_63_inst/mux_4  (
    .i0(\less_57_63_inst/o_3 ),
    .i1(i1[61]),
    .sel(\less_57_63_inst/diff_4 ),
    .o(\less_57_63_inst/o_4 ));
  AL_MUX \less_57_63_inst/mux_5  (
    .i0(\less_57_63_inst/o_4 ),
    .i1(i1[62]),
    .sel(\less_57_63_inst/diff_5 ),
    .o(\less_57_63_inst/o_5 ));
  AL_MUX \less_57_63_inst/mux_6  (
    .i0(\less_57_63_inst/o_5 ),
    .i1(i1[63]),
    .sel(\less_57_63_inst/diff_6 ),
    .o(less_57_63));
  xor \less_57_63_inst/xor_0  (\less_57_63_inst/diff_0 , i0[57], i1[57]);
  xor \less_57_63_inst/xor_1  (\less_57_63_inst/diff_1 , i0[58], i1[58]);
  xor \less_57_63_inst/xor_2  (\less_57_63_inst/diff_2 , i0[59], i1[59]);
  xor \less_57_63_inst/xor_3  (\less_57_63_inst/diff_3 , i0[60], i1[60]);
  xor \less_57_63_inst/xor_4  (\less_57_63_inst/diff_4 , i0[61], i1[61]);
  xor \less_57_63_inst/xor_5  (\less_57_63_inst/diff_5 , i0[62], i1[62]);
  xor \less_57_63_inst/xor_6  (\less_57_63_inst/diff_6 , i0[63], i1[63]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_10 (
    .i0(o_9),
    .i1(less_36_45),
    .sel(diff_36_45),
    .o(o_10));
  AL_MUX mux_11 (
    .i0(o_10),
    .i1(less_46_56),
    .sel(diff_46_56),
    .o(o_11));
  AL_MUX mux_12 (
    .i0(o_11),
    .i1(less_57_63),
    .sel(diff_57_63),
    .o(o));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o_6));
  AL_MUX mux_7 (
    .i0(o_6),
    .i1(less_12_18),
    .sel(diff_12_18),
    .o(o_7));
  AL_MUX mux_8 (
    .i0(o_7),
    .i1(less_19_26),
    .sel(diff_19_26),
    .o(o_8));
  AL_MUX mux_9 (
    .i0(o_8),
    .i1(less_27_35),
    .sel(diff_27_35),
    .o(o_9));

endmodule 

module eq_w8
  (
  i0,
  i1,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  output o;

  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[4]_i1[4_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;

  not none_diff (o, \or_or_or_xor_i0[0]_i_o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[4]_i1[4_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_or_xor_i0[4]_i1[4  (\or_or_xor_i0[4]_i1[4_o , \or_xor_i0[4]_i1[4]_o_o , \or_xor_i0[6]_i1[6]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \xor_i0[3]_i1[3]_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \xor_i0[7]_i1[7]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);

endmodule 

module ne_w2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output o;

  wire [1:0] diff;

  or any_diff (o, diff[0], diff[1]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);

endmodule 

module ne_w3
  (
  i0,
  i1,
  o
  );

  input [2:0] i0;
  input [2:0] i1;
  output o;

  wire [2:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_2 (diff[2], i0[2], i1[2]);

endmodule 

module add_pu8_mu8_o8
  (
  i0,
  i1,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  output [7:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_nb0;
  wire net_nb1;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;

  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);

endmodule 

module eq_w7
  (
  i0,
  i1,
  o
  );

  input [6:0] i0;
  input [6:0] i1;
  output o;

  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[3]_i1[3_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[5]_i1[5]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;

  not none_diff (o, \or_or_xor_i0[0]_i1[0_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_or_xor_i0[3]_i1[3_o );
  or \or_or_xor_i0[3]_i1[3  (\or_or_xor_i0[3]_i1[3_o , \or_xor_i0[3]_i1[3]_o_o , \or_xor_i0[5]_i1[5]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \xor_i0[4]_i1[4]_o );
  or \or_xor_i0[5]_i1[5]_o  (\or_xor_i0[5]_i1[5]_o_o , \xor_i0[5]_i1[5]_o , \xor_i0[6]_i1[6]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);

endmodule 

module eq_w6
  (
  i0,
  i1,
  o
  );

  input [5:0] i0;
  input [5:0] i1;
  output o;

  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;

  not none_diff (o, \or_or_xor_i0[0]_i1[0_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \or_xor_i0[4]_i1[4]_o_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_FADD
  (
  input a,
  input b,
  input c,
  output sum,
  output cout
  );

  wire prop;
  wire not_prop;
  wire sel_i0;
  wire sel_i1;

  xor u0 (prop, a, b);
  xor u1 (sum, prop, c);
  not u2 (not_prop, prop);
  and u3 (sel_i1, prop, c);
  and u4 (sel_i0, not_prop, a);
  or  u5 (cout, sel_i0, sel_i1);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

