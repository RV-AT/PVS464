module ISA68Bridge
(

);




endmodule

